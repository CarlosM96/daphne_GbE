

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MndbkmQgTx8/SiPqHkiZOQc2Og7HsnPGv6R762YhZQlkd4u7VGdD8IGkiw0uWRUu6oQdsfM1OaG9
WPWL29c2eQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uYgUbAMBWB393Bxd1Uwwk/JZMU+8OgH5Ff0hIkY7hTLYcp2m2I3qH7c3ic4QoxZ6Al+voEtVdAk5
Bix21hRZ2Y0am1rrEihQmx4ePyGPrmsSNCEQjGFVhcuS2jdqxYRbcztvxPnMnmA7z2sGgxlBvDca
2LUCcUabhGetrgqLRPw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oqgsGo1FvkqYDJXZwYKAlm2GwQouVHyr3oWltCkQfy4eDiq8e6dZtMYTvS2OptsCXxwhnt6dpFkV
aQPwWgI4M/EeWoFl0sJqSpzuKxw3clkzso1m+60ALM2kbDdmCRiPzqUp/agesGa5v97tktn3T6EU
BgYvmTcBujJumX/2YXO0JCzvDgj15zfmbIwFlBOPlf+5lHj1TDCyJHsleQSR9Aw+OaqgMxpV4mhY
KIV04+MC8ksfeSYXqZM6GbEdoTuQXQAZJzv3f93bNIadB93Qjw1ApTq3glmk6F504OeL4H4uFhb4
yrLA/+YVagpERJJyxq8aF8jV2cf8ecUQVWApJA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ot1qpsZGNYyIou1IaCBBPbZ84syWy7TKG1f/JPbtBkfaCKsScSnESpPe9sIEyscYmg2MtRaPN7AW
pPElR4ydaedMQf+P1JcgNOAfE7pZRVY8nidFZsYHLk1yqIYc7kZjeBd60Wo5rAwgqRN5Z5tVa1pI
Gjf6BjkRcJxSd3Tu227hWTzk73NbqcSK0eUT2OmuNYVI9IdHb/PF5TW46MpIdHW1dZegcarbIwLR
bwe2vnrYpJNkH1MPBuSnZN/mmW0kK15ZEUBpz6MZhQu6b5tP6+p4qUumkx43xvPki86TqWxHvjKy
yulQ+bFIKH7nyGHyWzM2izLOJ93wG0vdK4K7/A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PbJi+boZI6/u9MDnTENt2Rcb6pD7iRjIlP6ME83AndD2K/54TLrMalMeI7LTsr97UwTKUFhzjLF5
XKAzaDRI1Z/F0TOStSdDbTq2p7N+l9ugTgoLpWX5Yq3/aGpk6L00r2Fm5gSOceZIoCI6E6rvaEZq
2fE4A2nqlGPY7nD6Tgo=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
U41YN1XD2lvq5ZBC1dknnD/8+1FHs+DzbJIA/qcqrsNBOVhBgQ6QTIJSI1PPcUQpjrGr3zoN/eN6
Otg8vQ/qNLepw2AqzWc7J3PGDNuxYxVfXvNgBR5Y7czpYRo+g0OQqGUkdOAQbsfL3tC1KFD2mwtB
IwQwjBoP8jx29oDmAEUQ9T7Iv6Doit8ulo310hnw1KbbW18kAqDiczZLAdBvdWm9gmXduuf/XGv3
ekAT/xoctRBzyMw6/KLSAjnx7HBmWiwx3WDkoPfl2jfgWMmneVre3c+6nnHhmu+fZbx1P8zovjz+
gTiE+625Rd6WtxpBJM5iJaRSzwPBrlPDT72Lyw==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nvjVjtChOYYPiT3W2qQsbIogwQPRl90aNdsik9o6NVpzDFwS6AEfklc1U9kUuyE5ZqdYMi2XL264
4VfeTmZOGLAnNXvF+1qv2dH7JpycefgUtOdavuUUL9ES5QLHVP+imBnabbIyNbOtVt6lIBXhicmr
kwmT+J+dRdC2FTZ7hZhDfQRX/66b033JcoXE+EZj5yf7r6DC1f/IWvDOHfISdsXcUdlU3PbalCDy
94/1SFMc9/N/dnqYuxDczKydEBuchZeIouIdQu2vtSsoO9qNv8bH9eR3vXW8VzdH+Yf3W2d/FyMr
rwEaWhDQ+Ftm+RGc8A4ZXAj8zW/r/RMuWf8/cw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_11", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
brCdM6vu8hnAr06KwbGI6icCY+Q4rv/VITZPcy7/Z6aDlmsxgz96AuAPZVs7C2cafXg5UegZek1Y
EFhkIirLmjoPsTYAkmrMf2l/v/HwIusgZAU1KpriPLypXgjyuEXntQTnYIx9hNjVe9252xXf36vH
/XDflv9Z1YumzU4GMmYcHJiz5UHFxwk/87AWqlH6Hfn7fhCGrHoz984ffImxmPHL+cbGdzbcyh+v
kmF/lckbOBTnBfu/92OknPpBQFhAw8ZFwNyM2v9TJyZTwHgdfLLgG1H3nipJGCSh52D5OjoGsBQz
bXFA1ydpE9R+BTksgUhjJig5Oiv3yWHuu0PIyg==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BS6u5oDcP7egGpSYOQ+FbufBNbtK7LQ0P9+kszA+El74e/Sv6S0VyssuMGoaSJ8MnvgdnMFwhjxU
mZKo0GLtlzpNaE0RBile+d2hI8zREBXIwJcwXHDJKOQadE1wYhW+zsKRkjDgzGjLDicBbCi/grvC
r2LKMhUtHrtscGeT/udYOYiKOanwk+8PtmKh8shfZY9uvWocb8mfvEN4lwpxkl0c3c9X73MofBU4
9uPLacxSDOEsH201WRf+r5psiNmY0WmDZRFtUVIJwa12M73Ug2NEF3Lctmn09U/EtiPZHXEhFxQ4
ilXx2ACgw52aYJnXoGowv67zfz1dMVKcT9W63g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74240)
`protect data_block
HM4juvqhP/gHt02garvOODs2FCvZVj8LSdflV46ocRKSsVTgUMjlkxZuMY85pUZoEgW2ZLmXHwCJ
5qgqStd+TRU5JwlX8Dfc9uKHl4SyahNt3PZ27Axa4EGg3o4Kj5Nn+DkrdEJkDvQE77pqYGS1eTPC
5HJ+IlOj9gucJkUqpO4Y3f9vUz/XQKIrvWaMZH/VwIHJucREBX+b1b/5e6Bz6jX5CauYGDInwUVJ
K6H0z176gaU2kP84U7ltOaSRk/MFwh31cSZ8PSLt0dEi5UgJ2BeAAKO5O5FZ9GGMFHzaOIbAO3p7
ZUdDVbIh+COJJoK3PuqarcmWuyfwhth5Detok5+RDjBa5oDgQ8IUPuKfDwZTaPWyIPirFSSP0YLS
p48+VrbivNy41j8KFbVHcBX8/1Fs2lEEAMqAj3RRV+odFLbcGI6yRcdEYhe6g804sz+CUm5+TRlZ
55RwCnfAtnr2gIo+JZr2AaZpmO/4NUiOCcWMuyRWpuP/ZuxIgrZun5iKD1TRqXRsR/PhqR31UmVt
dxEalyBrExMS4jhj9ahDRGM5O9Fy9aVNN2erTvIGTxs9/VADqBok9zOkl88YByDGkK7u6GqJMWLE
BueHUjM5L0oUSd4RHgk3kvMunjF0mGdvOyBc92QYjSyRtVGeniqZ+raGK+p2NaXQkXmP+2imhDvs
3Gbf++KuSHFuXR55Ufk5fQShaxCcRSQC6yIzyzEIx99p2y2SzLS9DCZ/cdPPulODL4mWpmRRBaqA
Fv8jEbJjUDD94950uC2jB7zL2ODBT+nwUWQyR192mCwCNLAeClzM31Myw8unGM1fzg6JZtCwf/lS
45RWVKH0hbvXYvoUgaKirUW8onsPrYGsDbUm/a3OznTvAlMcS4QVheGcyUAkfvDsPR3fQJf6D1Ef
mbZSkMXQwUUSzNca5e84FaHQ7dIG/eSfFNx1plAMjkcCp8b9LcYRg2G5YE9ObQtH6yUR3UVwP3SS
3z8Jkd34BKtv4fT3Rj+wYDN1wpUkbth7y/aCCDXgWGFVUGvpMf7JBYT/fI1edfeyUw8F0ppNG6Lv
4+6yWuGHFgJsPL7JHcGJm1AtDn9HXPMcZ8NbElcSyXXkJ8ABtQ6unLigmZ5/43iIwgzhm07JWTxw
deUlVbxM9Jr7QAJzChx8XbCDY8ukyZvQueJhNWcDS1ttRkUxNSgF1gnjKoQqO4ShFwA7RSdYDEL6
gt97wXGhVH9WQ0vVPmxAAvYQ6pR3UY4UHR9+jOa28Y15OIgynrQQnXHZIQV68ghFK0+sY30sy04W
3cqMNrzP7AvRdyC0koSReKFnL3YL2kmati2XSwVXGZqkgvFUAKI1I3PpDoFYuuuJyIBus8+CY9Sy
uP5PlrJ6SydCRZ0c830Sr7SC6xwuMJm6Y+qvvBTZkpHsP41gxKwTbDiD/qSbIHf34j6nwWCColkf
60zTQMLjifcWMcV8tLtUneP7tJ10voAD4ILrM3Pxc/vZa21sTNYbXarBRTBxNtqDeT0gdNy1mpEY
IoBUbWzxcL1q6S1lKnyAu7DBmSTBnXY/hXa4NA/bKvLI8fH9CHA1GAKd3S+wsw/6SzeSS9aRTZ63
VNBmYXdZB4rJTudbC+2gNve81Y9tZaydH/TbZHwotCjyDFc0kM/A+Irf5F1mdMO2h4mjF86PasZ9
3zW6DoS/n6qMScAhPE/H/cVTzig4GN9D6YH+tVB1FdOPvBs8LNrQMJmPSl/wdOa5s88vW25K0vSh
ASjvLAoFO73yO/SZg/ecg/7QE0O512oeQ1xFy0wYauSgjYEDiV7v/aD/pyzIPILXmS2Pv1MRlbpj
x2BUf9FlgkY0mJ+G7jVbcdGTrDwwvzjzfO/EB2yor3N4AjsPC/Hfli2YRt64Nv++zTWhZYHjsg49
3ku3S6aOkvJgAritu1P1dv8oxBRvEA8rfQoNxZhtSOIBAdM++5c627HuoqORIeEBQRSUDmGxRqog
vAnPR0I4c6B3FAJ9PY9Jkw1M5U9KmwgOJBGUGtN7x3iXPVXgqo7oKbwO+G5P9Ogk5VeqGxRlLE6v
LhabK3JEVfViaWFnAkUZ7MR47MPikc3AkdjUt1d0WwaltUdObta+8HoAnOdZTvub3lJMQGnt3b4B
N0FHyX2JTjieV85tZpl8l+nEW/Wex0Rt3AoWVbzfUUxTsJiNJpXbpFtdEcSgSGB551if2q1DMQ9L
JKiWZH6iYckBULHqzHTgxTx8zzytZyMFAKCBxfXCTiwXBT2UZxJJ+qZxdnoa27OqNxj3AMqgUFcE
lp7nzh3Dh/2EGmdZnImE+cStjbm/TEZXjKbbsGaKu12Sd5jsWPP295ILaSkXImbGclvswIhmP7fk
NThUU2IrGD7GyY7hRefzqgLJwF6A4+0AKiX2t3sVwGR4tOlAqkOZAEaHCaWNZJWv+JGYgYLOWMP+
ckcX394xl98LZiQLka3yXzzJZLFmP3mIGquOnaOzWhfE1ZJg1fJGLWuxQTywQcPA6cbUY/wwh5/E
nDX3exmXVM9+tXivKxIYOZs19xRssAOFn427zFTgbU3ERe2lLVDVhJFsth1+4C3KkrP9dwK71c/P
x5YqjPyuzdkPE9WMy27BdBfrt8huhT93YtR2sCxFeGVthn7zAbe+df6zl7GAarMuT/VuUaXzN0kB
ASefahV6lif2i1Y6ezFK/mzNUrLiwnHrARf72qT7gYmbyLROq8S/UxWoPV7lxbm6nftEgsuWUnR9
+12WrN3oS/v3EPF0akkilu9ItZS1+PDPLOyKXgInghuZQxv8OgTBCkR4JaRZad2A3NW/02WtiaIT
j19BiPbXleacky0qzzSiFHmCbmZqzXDvyW+sc3z5XWGUdbcODgO5z2sgsbBcOWQ9f76S7wJNUEXV
gJ+v9utk8ViDasa1Ng9djI18gsuzM5cpqd2NYMJBCBlOkV0K4sTy8it+LnceKJ2L3HRSoryEd8rA
WcMAt1ndv0UpflvIz1alKByws4r7Do27ZrDhzJymZhRSS6A9qYM2nSBndeVeq1FsY+mVvvyXqzh9
AWbG+KGzQN4M/NjNAT4W4vW36RGpwka49kknCfOukx1JscE9/qRCv20UFyoA9WPqbPuJMbYpok3y
JHlAPohglJEpgFrF3xZxMOsQbftBoYsTkgmySLInvTTURBDmSN3wyfFITnMg/mNGcHXnou6riBjx
WMq8/dcWk3gkdPDAPN4E5L5ReVGF1iVzQP+exMkBdLOIso68Sed/hYZpDAuAvKkYbSmw3/0OKGii
C3S7AqRt4wkkLcZUH0RYHz1uD+4VF3+ACMdCebLujM7V7QBGc6weqm608IdCZCR3OgHI1QzA+aXX
dCSfjPj2ZQkx13F5EcWEqRUzxpzwZpIR9hszWjODYGKFeNQ/jHMzkNRuYQvHsnCA8JkuymLbJHO2
kmO3zxutyb+LXUJYKr3UCSyor6Rm3OQC93iDt6ih99dw7Lcg03vUiDPhGDNU1G530GzXjNaqAZEA
dNTcOCH1Kq5kybfJ9rdj05vdz/HyjP55iZIZYnQOm1U9sgF02rOBTGf14QS6gs/VOAFIlDVIiwd4
8n/D4kk3jN/uqOXuldonmAxHf9u7pYkfcpm3tBnRIDWib85BHUKLIsg1JVUtSBQFVoQULbZZINSE
CqXlUO1u94tv8Ugb6LI7dMiTacwh4TN1lqo5dk/nO+LFa3Adayw8iMLvkxnsL342UFnDVc1uD5j3
lWMSolewXMdPBkUO8u/iOQL+XD+2gbHsfU4Clal4CbQTRnmDCYkANndg5TKbdtaligySKFGG5dW3
uniw5UeHRu7mVql+XjKwRZw/VuH4/yB69TIGtNVfsM4VXT0mKNcUv6dbYLP6FXe8Zs0FgfuBVcBM
mehBM1Jhyhpxs1PWBeOLPXfQ8HFE4ZdX3C5aPtd5ao5YMtG1GszwzZPhuxqP/H/c3BVUYxbscqJy
Nk+KctfSAwKNQZ/YDZBSVk4n5yhcdKxsSGibaC3mzr/0lCdjFqDVR6ujYWBSqEyhTuVyVSUZQa7g
XkZb/vgAqvgw70nqnndKsoM2Uuy0+YcsGdpcZNXukEo6eN5vgfZq4UY7hSkDZFLGiMmzJmcyFd6c
HsT4kZV7RWRuBiXpqdXTskBFFDaiRcIilqpOS2pX6Of+tYbNy7pdz2Jesl92RbaBGtrRWKZPpMHl
xsPPFGgPE1N+j1pWmSAlEzmVnfr0v0PGrvxVdjPynwoVUwy6hhNjQysw7p1kW9t5tytK8dxrNgLl
XpNHHYtesndgTWg+p15vwjjwn5H8fFu0HsqEnYskaYDC2pgszqxcbUEFUPtKkHT/Ge6/xxYIprj+
NPcRbBp8QbDjKQoBa7G6/NrMbi+Csa2W7NUq8lnrhIezIP5p0P/+bSoZ4BH0op/PYbHQX49EE81x
mMEIzhcb6pE/E5txDS3sznKVBZplWun5Ui56b+6hMi92F0dudsbwdUfGdLPRtUI4oVNxOmWmsU9q
g7Bx4B6NBTS1J1zQXs+i4T5mwhdUxH8vro3IorUhirljghpPs6glhzeqLizMyOJXI4HZ/aAgetr1
z0bk/SrQZ4HZtmadtRjOOIC2LWswVC0opqxHhALnzzvqFoe/qRINoVSwMt9AkJNSI4ApqeljMGQQ
NYO9lbOa3IkJY5sNpwJKHFXQOqtv/1tIbmnR9emhBjuW8oV1choO61XWfEAJ8+c2GsCY7FT7aZEB
UUyVMx4CgYo7h4/TAxpmZn9AUruKaGXnBSby+fg69bo0pv7yhURjAmiCQSLa5xxFvSz/RDZ/C70r
0M+m3d2vJUFAvjFWl6GLdRvgOTdZ2jJ1WXFZfzE4S+DtwbQhPp81cydDh6ZiHbRU0fE3oomM1cVi
0nfo8LKAkJZ9cg7ozeBcLMelUi5NDSkcLG2dnmmAxBRhra1HFfHO5n1ofVv0Kq8GR7w/A5OzTTlU
H3ybu2v7CD1lVA10ZdVwQIxYhOB0+yF3PSStBT3bHDCxdFiZ27KkS1Tj+QZYQ43mGJV1YpardQ0y
7YXttvD4iLmCVVhZmSaCEQfPIk40/jHGmOzzKHNsUSdw1uJqYxhQyPOYOVhra3GBzE7muDuFLqOe
8a68ClT/12cc3zCR28FQrwIc3HI0Qg0EabYBZc9qeNG39IZxzN+P2Le16meHRo/CFO7PqXnyAukH
PwaDWQkyLIHVA2c/ypOxqJ+kEXgzthKpZe11sqI3ARWE3Lx/TOcu/uzDCB3phVNszKIuELae2ri6
4g1PTQhT9gPHVPjWAKr042uu7jFquybyVcSrifiDSTIN0oK+lBoJFqdOqvt0ugvIrCibxQ2WI7J9
MUeugJpEGKKKST/kHntmUnlPfrF4vSPjKCgZrlQnT3m3KD2aeRR62nS88y7aKSEHx6acD2brghFj
OyGkQrBMrGwGNKQ74cv3lohdsVYfJPThDjIVYGZO9y0gcQLeiyVH6ELN+umbb6tBaE6P2qxs9Avt
T1RB5QBx8Ehz8x2jW7leAdblGbP93byt7dbIqB2Tg7y53ZPAvBwq+0Fl9OqNMNYITTn8qXmuszWG
auFwRQUbXo+VWFgffRQ6bIRUVlBWzN0snnoRjkHOmeW2s6VaGUwfnPUyPQwmLJ5sNU4WwjDogUVz
oB4INvSL7DHzioR9RfADOq8+vS9l5eKDNrRenEL/WkXa2FBeB7DwRNZ7gAeScQio+wS5oZE/kCrQ
iofR9LrZjlFf8AD9UN8KrV3rvU9U/sptAE96mscvgGKcrNqXRh5J56JT388VcO2ZJZO89Zlfdzui
UjP30LmyZ46bpe6YzcMJDPRHso7ZPcvu7rR0jh+b0K+huXtENNNd/PqIJEZ/edrYTFZE1cpcwbsW
DNpctlmSKL2fev/ffqz5ur952uZnkNlyuT4Q7LJ8Z22YDfzU8+zynN2YaONkC/VI2URTNJT/htNb
VpLSBDYvdWixC2V8lPRM5jVfcVpUcZ4q4LTORlbov8V22B275TDxfBcgy5UB3eF0G60tRRGQznbd
L4QSUvZz70jFGFLpR58SfT7ZtCQC5Um2Row9roHUOH9ZOUvpJHaOJKDX1n1hTqMGhQ9MIC0zadIK
tjuFD1t4OsReFsNk7Qi0WBiI1qMNTt7ClxzFQjtBD6JWXjuqwkhfcAfDuc8bwxpAMnxdhR6S4EYz
AAF2AUWR9BvgebE5ZAsAB2oI+UygdMTIzUhiti89K/TpMRjRqR+CSVuSS1n1c6dkoPnWk5vHBwLf
F7C98gvwpJAxv0s0KH8KzcLjwOWsaRbKBNYKCKrhwuil59WrIsUIiU8NJq9aO1TJe3Dm7SpfgeMe
Ce0Rg64Jex0S3XwYavHgX1+phj3fchK1ERudTwmXurNNMV/X8mFGp1XB5OpoOaoLOrBHsQY80lF9
nSTNofN2/HVfi+5WcecpB5qsfm/qw+tG7kg7PePeE2TBPPlWsP1GzqCvErdOtP9t2JkWtOa0HYwX
stRs4VE1g7NoIdiyn3Ejxed8OM9K3hSM/Ln+qFFtbYLttvVVUUy4WfsA4v25xWV80rBAuIraFzvV
MgoY1zDznU7QatDS2CzUwIL/sHB+76awymNL6n2McTIjnrmEVTRdxsN6jUC6TNODGCuq98CWq2D1
vqgGfl4B//kI3xlxrKmdQ++pEFkfBmCwwsJSNTUZhegstJkXJM65VXcvqWkRLvTPkAtGkGv0lIzd
VMfCinEalKKNMULDUxAFRLeb0HjF7D9hu00EtvxHpgMMzlEuQy3dDpMuU/jQo/wojMwGCdNZNYvu
vKry4EmrYgspaO3jv2fChfIUCHUw/5JwMVCFafZMyMSR2tqvb25KRKXP0qysXdO44av8GQK4DTsh
UwBh7jWJCZ+TR5XepcOWEeiPk8H5ZH6UB+bbe4gWuyjsk0R8UuIbCaeFvO3hJXkF3kwtWSmzQxyz
tyM1BJ9wnBPVfWyQ7ViY1TCqMp9tOln4WrpXJbrjN4HM09psl6pdNA97LwALPLV8sM8FwVxrh+yl
wCqC4bi2vHaLHfcpn0GfkPdN/7KCsY+NcFT+8d6T6EBm28w5OsR5Z8H6lZM8nYeZLrcfPcV3D3hb
ARl0ezgZWffHTpMwFxrWWY6tCVbribpIBtrIgigIoPpWR5MXyreq1DTt7ujRcU3AvHXmU1hD6D48
sxQqlzK8Y5dXqDIOPztvHmtMT42MxROmkeiS+IM+IZHlWfJ3nLb4WBMF4vaizXJgSP58uHQUgY1Z
gZLCb+RZKDiTdK9yhtarTUwvyZ5Gx4EpoVOfXufpn0F9958v5avGhFXff1ZtGtAAzioG8+62rwQZ
Z0oE+36zBJsAUw/8zWMANAMCixp7CTPqH1ja0lK0GvY3rOthEAkvHMjVGLWarS/ujWTg4w30fJWi
NJvDE7LG35nN6xfvJM2nm/+RY1n0dOJh7js36iN7vU97Ngd7uKK9Zhq8/PTsmuVJc3rYEY/tEal4
lk9fp3oYo3dyetmeDMLCJMjhAknkM/ycJQHmPbq4TZiPH/mAemRlnZfXHS9O3Jhi3LlhlyJ+BsRF
XRMcAtaMSgY9LUekjvFuU9Y3OAtzHgAgYsv1A119Cb3qYEgFMDvgRw+9Bx3BO8MtPDvwtu/h/2cM
UnEPNiju0gS/V24j3q4OdpsS294McVqGDlnmay7n9b2j0MeIwWPRXlKO22RpOWHA52Ukruyou5tO
WDllTSxgOrpuuqZRrnrUBwjw81t+LbKsJuyEdA7b3R/mgGHdBdG9MvkF0Rf5ENuziEbXRFEFK9C5
K1WmP8NKEbg2c/2dc11YfwFMhjiwMj5ianlznmyEVuDmXzfkULndmyfbFWA1dnVzKxqyex4Ppp6n
Sr95nu0MiKzLoHhPZlpRjERhW1q0nNCSkckAb3uEu4MgYRsJDNge/Ho+pAY6CQC1rindZdy6dP2z
oAVV2scj9y7iRj5KmWFR9Rp8wPn4v8YhVYOxC9aCCGrSzwuC4jlXs6z8dvcF7K2VaZGQXdTrgxFR
zhfOKIeM1ZzxTNJfcFQnb7zLspZNZ4EbMH2GtJOqgcQJn1jKwcVdKmDs9nDv4BxpP7e/ahxx6GWp
gyVEXUpy7Tjhjg83gzaBN8C+Nqml9o0UsGOMgxdANBjH+lLRC7hFMSLnrQ5fQf36eRl7+UYk4llv
N5i9O8QG0Lv7QEBuDnmFW6dCWRJqzjDrk7NDX1VvGAgBLVBu9LmrDwXn6S72ndgRxuVqBDwxARfu
2iABf+txnte/ycsW8nRGfJgVa2jkXzDAxT4eHhhcE0rPPbjBmW0jFz6lSQFcjXPG1TP/o+Zx3SJN
7CZ8sUDBZNnI7tnN1rLD3wxoT+cptMG1OVsNHtki+bOBYdi1tbDZrEXOfuyta0IqHw9zjXmf6N31
xKfcftWt4EK0mNViNaPKCs3llCTDNZxI3KthIALm5D4YEAnfNdeCEUs1NxWGs8Sw8FuBhdB5QV01
YzXpaMGZtVQBd4BvtwxTtuiBbXHeh9aaSogQN2Ot+HMlW+F1jrPW6BOAf9nbgIB93a9fZaGLvx6C
9O6sUiI9h1KyBlaLN5wZyVw87npZo4vyWNuCHsBcsqnN7CvWPyjLahvta6syBXSlIQRA2HqgoJAR
0jiAeZmrgHbx5xmijD0rZu/AJ2OxDJNbWwYV6TDntaZTafx0hjibRZ8StZQUrfnVmiIplSnabi7w
JNcpPLX2UQKuJRHa8hJrn0wIEYrpQpaafj0drAg9C5q/BGnM/V4ZnHInZXRxJhb1j73K3oWBUd3W
nAUdmK3PjcA4tDbwIT7faP2hpPOw6XmKyeMBuh3PdZ9XN0J4bDJNkUeYC0Mt0ZG72lh2oMSQkwhr
tgXqnbMMPcOhv5HPJX8p1BcSI3X3Vd6rfADgXf3NWS2/rZZAuJvhmFvhJCDUlcs+g7MZkc5OXrkB
GDE+gcbl+Yos/fvSYFT1XyQRay+3mzzzssvMAnZB/1aHKrjvErrkGrU5nyST/EElkWqTjSNt0UHY
4GQUzRiE5zMPXbfEOocs3R4woAzyf+eh3XCiGbFYRXW3J5Xv2nkrNCqBHEF9OygKiD2kzU+W1JJV
QVgcS5aQADfmzd9cf/JyH+6TEQQArh6GjBz0VFSoB7+L9LOCqZKcHVh4ZFwnIiYNdj4TGpTlvi6a
zo2gCKr/wm7QX64g7tUzJqYWM61MiAik0FJ7h+Xa0Kx7IhTpoguUCXFR8ZOAQ6Or9CpzEdHhI8g9
yOoW3sviqFKqfHPrxuVOryP8gaVh/8nLmlIb6jKmwL11qV2+gHGDsSOer55K/uVxllzZxjwZeXV7
aXxf8PU4cbkGFtKWRqkv3lQRyTFLkrdQJ6LnTyniY3qNZEDSZYZ7gd0IylPszx4BeaGaixvITavx
hXTA5CZiwK/cRa79m7W945iouQltZWHLwlya8DjpEgsBzSxHhQfJyli6tIF4UEGZ30VeJQG8Rh5T
IUrX77beLh+T2VkcK5gr0DBNf87gI714tatM1520mIKabXapIaZ6LdqTNFPklOqEfGzhpxPGxDBq
r1ayOVUP0te28Yj9Ync8qNMSK4yaGMSNS+zfqjaUbjEWMHBCmTSWRI3rQIz5md1uPRx0LaAr6qsu
eYdCq1r9K46UkY+Qfg6oBqkLlo3HN0z7m3dFaT5KGu5Iw1tw3rMQ42U/SVMpUKA0iGMEdNZjiiui
d7u0BMEVl5lhrm0JUno36Q4ee7ZYpWbgPK9Ai0fH4fnU5QgjTNCoygERxTZz3wI6DaWjulqsfFl6
L9Fb6WxMPoAX421IytWSrEbfK1EPqpyMAmV/EpdfsFPM7YgIRk/7r9MCfFRDDt6f8+qUCTE7jsq0
WZwnSVN+9Ou/JErAeTVi+C5MHluNGxDTPZGB+T6sCv5pR9dGaz00ztAhdSlGGbxYswkxhDLTi24i
CH+5VlIy8JcfLKJ3pWWxSWTZypu4FFn3y0kIzM8ksgw5wihKk8VcNfpo/MJvlIFU+hyRHxgwEEBJ
2qcLRtKtrSmehdpV+fN/kY+IIqapGqD+IJ1a8Ogq5Xa2vaGWh1DjR0QZvHQmfwApagmGtRDJDYa8
pjQuHfG47ZJfCwPUMuHJVKS8D5LZLrW9w5UKdO0b1+Pht7fUV2b5jEkvKljfjT1Q6hrB8mHJo4iK
MOMFT01eh5sMRObfhvU/kd517+Oz4UufKgWoqDYBPL+IELwtyY0jVPIvDRHoxhyPvfzEmlLCeu55
ZB+wPDwTmHXshGGKPTlaOWWNG8uIs+BDX/Igm0v6s9TJuUMHt+syaZyG1XPQyRfXPeeeWWBsmAJS
pdH9i4yiEld43qc1DJrA4SY8qm4gLUZ4d1HSJ/b0nTaNckQwSc31CRSeBJ0OD61UYPCfwQRv70cD
bB57vBYeOHP2vj2ilTjUl7aOrwyFnE1i1a+3nu9o4oHRD63l6egdsXIiOYx6BuHESxSv66negN6C
kSu49fK/tNvWyKYydiyf8/m92lYjk1iS4AoaMWWtQPoVX0E8+tQT+gDC4vi2rCOkpolvh4DXQhbb
ue3JrdekhxThmRJ2T91D91UZdie0J9WBlNlNuPjxhtTu4mTz85sdWiYnwWbfxdO9bemWWnc/fdoA
WOg2eUn+UXoeF/ICAGlrJdYr2mqZfa791H44G1RkYURlX3EhEOrPlTGx3z0hEzEUnpMK5YPyV8QH
ujsQfDcXJVXvr7Wm7y6/plsnjBuaWG/kDwrSxhsGflodRGcg2iAnugIvHxn4Ikg9LGvdrW5Ev76w
Kg1rYIKWys87dyIoyEOcYSPk+WCtDjSlW4aRPVulo0BELmESV+TFvz+3H4AFb9sqUE2LYdFpY1Ml
6kkt0BgL9ekntQVaOJCuQC4EvCqGwvXWh0TWj2jKY8PoFkgS0VDq9KGTGTATuhT6f2mzefCn4z3s
yJ1BKkOCed14V4YPWzEYO46l7A6JFnB9zbX5h+3hQbx4pkUmLhdlJNQHsTnYtT8xxk/L/WgDRjXk
Q1Sx6fEVWKVfG1ezjsR6nWSNeOX6h/EwzKOIpq7Q2LQ39rJdiDbUsLxvWATW4kZTjPhg62NNUAss
D6EHb5f/ubOhnPBO8MxKphipG8+vVEw9b4pqiXDlmpp0QjRw3lZNs8fUmuZU0pK/97RUVpfKovwQ
GAKrMJc1IS3EVLK7lk4MLOj7kWT0/43xhclw0fqWbehiNu46DxPXfFqEjXLJa5QnakRHpX44XjXh
omP28QUb6tHjr4qtYevufuV5UCLeMaww48JKzXGzMmTMYWFIqXoIypGWJsnMe/Q13gAcwILoV1XZ
n5PWl/uQMdZDwm2TuLayPls8M9QPn5nH3/79SKlyU5PXzsBkMakSE8Hf2OaUJWFohw0kk1HLwhSj
9r238yz4HmwNT4YMWqBri5xqPKO8bqQlpFNVXlTk3c3KwdfdLpHYmSPLvQvwxlGkZpjXdwtI859e
OrUoPotVL0GCTUSe+2KUXECtA1wrv43Vcc00W6hIf7clJ3BYTWJd8B33zig+SNkXWSULeXGoc+yG
TJRmadkM/JSQfhexqPMty4aRT87x6MgZgnQN1yP+Wwsd7tXrdzR3CiXzAflb5Shy+SQm9UfGaHhp
iVsTbUDZU2uTg7AluqCxOGC6vnzTiNWCqsFxnW3fRvAvHvUOKCLVYrgPUB9NrnjeEE60bjXFwR2e
z1VKOvgplPlaVlHXSbNierbjwyh5HKoe6CVB2MxXUqNk4vPKWOCX5Ji7B9o/iiBVckGUPdEApsa5
x3y8/RndsjjYXVMJWX819GvRYNJX5AJHStlljgZNxUoUzNIOiYtAiQg46UwR4CdIAFZ/VD8v0BiW
Vl5yEiDR090DSxIUb/lOGx2rhvqH4FPEhPwdRa6VIztS9OvDUcHEWqm7UOJXqFXWZtAPqU/XEdWS
cqLKtazW77SsvcVkdjtZz+FAopboZSJANvIyK+zrUj6kN6Yga6NzRlWDos5pOUd2DY5JznrXGitI
ewj5hXQI/uMEfHenkzZkfBGW4iou998011algbH6mcsPLAoEXh5uQB9XW3C17pzn7NSmDembg3UZ
5ChXcN3O8gyAyYbpeAi3MuFGNSp1kyob7S85g5Pnbb7ftyZoRD7cB3QR/okjYDuMcCTNAF+iix2k
MBZq66FjKXgK3ESDAwD6l1Lh0G5PBVvL7tsuVg8AldaeKsZ13D8+As5ZjO7kQ9F1Rb8M5YPMFaaL
6U1VPd173IUyrBN6Zkc4jSt/vU6YD1itBhBCogt6uRVuSTYZc/E346UhM0pr3/LaJubfRvx0XYM0
cBzAS0bodyvAlloqTaO585dGBXkWoYL5PXpxg6f1Ss0ViArbuavkEgQvsMiOiCu5aocI3Clq8lwT
/CCXc6bgvIBJlmvSxq1zOcWq51QZ4Ruyzm/igPXYN1m/ov3EJZWsFUqvTw2qSLpWn+U+WBd1g6M2
S3jW052ravR+92yCyxQqZEg71EQg0K0AWk4CvbI6dAMpdXvApA+Da5DQWm213Zt0QDaHrVkCWA23
4i7AZeXewRI3QDW+QZ5+uzafW9ImoVlWP4yWKDcfivPnW1ch/GMunNUc3xloGY/6HcPakZ7+RajF
DJrzh6H6TM7YFFdpIEAm9QkaHfH0Xq4MWtgFLQx+9rgSIWrs0zuI3d43UASgaQgVNi09EgmO2dif
yVbyfRmqP8pXNSj/BAxJvBDnvyzfVsAgj02ftWNkWxgpUgeR1TPfquK4ovhL6QWuTc3SzUk1z2fo
MrxRNz3obaguJDSrPKw6vrhmhhPKplk74RXJd9Yw8IX0eQXjRWHkxKddZ0e22SCw+a+f8MuAzkkn
51+j0ZznE1Ae+QlWNZ67Vjyo4RNAZ3VqZhla/YEl2k8/s8Xy9YBNCL0JtF/uR6GCwn+6gjmNpCNK
ool2/Ui2mgZv3onzwxGyjnKy1gHnls6NlwGebOKjSezKbf8AXlfzvQLItc4IWLgCxLcsdmCzvJYH
fpKYRTxfMISksnwsu9EqfL1+9ysY6p4Wh9t//+wLJfKW5Jhmwwxr4TTY4Q2A0jBEwliGW61DrYh1
dz05VgIv2VaVGyO+7Nqvl2zHOiCqVlK0sD2/7chW0hUca0GwTmAHabmQscDizylbD5cHh304sKzb
Q0aI+NsnuNmw7YrhT9lYQKPooCIper7+2S02JSFqjdLWurkSDbjiBelIdvpiiG8+DQ36dUzS3W2z
RfuwEfJiHAKfwan+OR9tU52Hql/OMHHkkzL29FnV+3eTXX6qAu++hbThGRbZOfTgDyRz7cYrj2Fh
wJLiVNRpM1SPB02SlBT0ef9pUt5l6d3wWzbMMk7hNzlDlX36PQ4CSdGE3BIaZrpKPmhR6ifMY2kl
4Lrlwd0JI2yLXJYG9T5rYwNBiha+222Cv5NdevMhIcfVqGN5hmlfMPap0e4VvA2Y78sgWt+VcmkG
LmpT/PYdxbkjgtHXUaqRZFBSyUoTVxpl5SSlx2iemE2nwcEgs05lqLhltiqxcW7yZXZBEw1nYzUu
AEPytKIk3IKbbbahSTait7wOb3VCh2E7gC2AAY+0oJh3Qz0/6gSLLo1JVbJ9HJf00OHlnyT5LvTC
n2yvBDjAW/LZw5ZFQl04ou7gha07A/naq2fnr2hzR/jvYh2kYTqAMlDMTLIG724b+M5Do4G85+R5
1uZmrUNi1ecqq91b3wKCvVRitdsgRWNgACGrCF+0ijz/Xk7RPGDJDtJSCp6yfRJoH/BHiKIH23ay
lvG/TvJI/PF3bBdSXQF57cihKjN9is6VsgdAzHx5J/x+ZdZmAk7K/cyur9Joa975VEodCA0BDAhO
wsbd0WzXhkCOiNHpeMxdrthmxuHcZ4HpHLfY/YoqFBzY3pNJnaqI6QmJ3l1GZqbFXf/6JxV+2klo
iLzr9s6DdxSg2Vc7xyUqrIqXSJuLx1lVsvW6YmAeKFWF40IqxYuya8AjFc33CFXbbBV1I/6yTR8y
46FaK/DszFo//Iprt2csa0wbfOfGX7mBAmIC/6Q5bYBOHx/nv1v+7MP+mcfq3jBs8Xk2EjJOiL0e
prG216oiVFogQZUxHTdfw2Zlmn9itOIq7YuRXdAAMBDs6iEH9D+TCe8kZ5I8x1AfoESiI0OnnbS9
c0C0NkBUPhEne1ohRAoaKowHLduRuHi3YR1joXUxDurht2TUErIVp0R7oA7C8KDfYPneN3pAUrW8
lYB/dvDGuzcthVdYn7Loaol7zMVaoQW5NFSeAk4geJmiCKgyht8/QBll88vcpZzeTdsDMoshmb0d
kyqU/LWSGVGkA87rDetVvvZhahw6W4aN2rU5HnrNBd3rPDH9NkrJkTlvBp4sXNVHS4MBcwD0brOO
t38lwumVtzVhS5Ha+b3HXLqoMbiOeuuHvbzjDdjGpXwg+CAKG+GDbIDx3X2V714vEWcK6qEbFN4Z
Mh0pjRtKz93HrooVbAw7wGZ0iDmkIypszsmMEdg6yQ0q4BvYI3VlpokIFyZNMtN6LsaZq97AZZ6a
AHGIvc/dVtwuwY7jOM9+B0uOWxTg/76dgGC41bK9p7305H5B4PP364ZLOsCuyYyVBVZAoJAO3uMo
GLtezvcKPuMWxSuEScSIGufm6ZxQ4emcncRf3K1bHkogi+Atm/G5VI8T7r1i1+50z9HnpR9nf4pG
hq4kDOWjq6XnASBMANc9ro6/1w9ZxwqbG/3yur4zfwvceSVonT5WO6Ae5errW7SdYX6im7Wp4xEh
0aRLLDRDBGkjhUklu+xiqlHmwtv5hHRahuRjNl3TRY4F4q/tGlBF07VkEvTei1+Z3FtlstanATQB
UgqYAOddfgt03byI9uZf3sTWNR2/3wW15q6dca+JpxzxsRePMbCuVXbvV61wuhC3QYz7IDVHgOk8
FwFotrNIe6ZA3tNzSfWhjZ0Gl11qnMk2faLxDVBF2somTkJASxVNRPUBLuOpJE8pgtGtIwZ0+g1R
H7XcxP3igFZZHrvp9bV4IvZJt57wGjalFMVjlOI2qWpeaPmDX0JDfG8qppmKRodK7PVLPEHFrY4d
DXM0YJYubEHVPNLW8zLm9TKBTNF3KgiEUZRS4omec0aF8Ct1qqX+6xUE+aVj/p+fdm5tCCL1CHkf
j6mE5MlQ2IBSWb6OuI7ZSDgbYIkoAKfFCqY1O/CJ2h3olrUjofcN8yJM8337nZ36svS7r+eldG+w
cvQHbxvn+NLjm1N7lRiKV7en2uAmzQHqG0QXBwrIEiQ78s9ltX6q1cERdwmba1vZ6CgR7yTtw5MW
+Uu6/TF/+eZLt3zF8cB2UOw28bs/F6kce60QtAWMsyxTuaoFA1JNNnxzU39RdEAvBBAcFUfEVYnm
aVNDs4mR5tEJ2whUN9vjPzIgVzYbBpXvFnkxZy7gkw09xfVI96HpIFYoqnJD2I7o5lGY9ukplqOv
SRuEtAOyQtZVQWkDjTgosvhwAvZpis4K6Wn5aQ63CNhohXufBpmgNwF/vqY6VCX4am80Kt6A65sc
tOPed8+C3yEAgBzjaSujfAoZPtvknwmiG/UJdo99Glz6tfUU40LfG2dGi42caSOdGTGFXvDlC4Am
c9cYxp5ZqrLs8TD4ZMz0DfqbYB2YEX4W7TglasoJ+Bi6AtLQlB9HkGmtKu+djDm0hXPxuCWfrCRY
+GqNbGcb8kc9/qC/0X8UkBH7Pz6MFYONbIBx81woC46/7YJQCS7a3fNr82VhOtZfsfKBovx0ICsX
dTG4NleX27rq5UQNl2v9v7Sv18La41h69cTEpfFR/XT/pMs4lnh5wTv4qlabRdnU52EHg418DJS9
HQW79lAMWf7KpCjuYjK/V3PDyyzVbS8Jqe1ENeLvxMTxb5b8kLGTqIYyKGNpVEPg3PUvz03FrgnY
IHyJM8b3IV+fxBffj8KLBTocijiZ8wfSxD1FR8i9m25j4mJm4hWnGx/NW1NRnEMsewp8TcpsPZZR
JbbrVi8GY+yijOdAT7qDFTKKivZCXf3nCRo7vQ2NSr2JVT5urkB2LknhrRQsDui4X9nKoxGQgLjj
ZELNBCQVcktJVGSGADI51kULXNhyRmxY9rDhegTwkRtsY1qAYeg/VXiJTg3ru2QSaYjB6OcUI39O
BlhpJRrqVPSBbrrQZMgGblFXZNfpt4r/CynZnOlGMpO+sc9/vGPyf3snhuYM1qi925QhigHraHWO
pw3oAsTmZfRwFG9dyJ5LwMgTcD8Wm20OPwERbTNPZVxAa+ITGt5k0S/LXuTrtfLl+QLB5ScQtvzM
7QlhtASmZtH2XHtrTJl16Yx7Z6Eu5Vaxe4WJqg0lkmSOJ6aL7xZIkjeCd5mehl28zij8lzyciZwW
EUmpCdh8O47gQ4ytd8kmoLxrtclZhi2R4HZ6oLHb/VOX2NCgH7WHVN6/A943oEQTSVFVL3DAfE1H
rz5KLAlnCWhnef42sTf9mee3gYasu/0b0GrKRU8RcbCzonuUR/UG7h2Tz6UwxKeLu4tEqzYzE4d6
Ru997EnQ22QKXIiMMfvJJ3TXx8EHip/DW/j9HCct8CErWs1GpJrhf5ozUqPrA5EcC0LDQuCn0lr8
g5eX8nTtMJLedkdcxCJGUO23WNEN7yDD17HXSnpuXd0ugFQi2Ez67d5MC1/yBPZGgXWx850QlQI5
btAvmBjYZtgFo4PHNx5OP9PP0sgddvoo496vYqv1EtSSv6UkFXnmVrNl9jLJ7x9G1pCOaBnullX0
oIe12oaXJy728hmgYvIJ+ciBEBfQ5sd5Xle2TAoP+hNpQdMD2u7O63gezzE1WmOwQanyJ/Vos6qX
86POXOqLinDlB2HR3OzritgdFgGpQJipnqHQJDRFXee5ziCAEEtRfertO4CJlUYjVFQg4HqAXFra
ij0pW8gGyPb4NJ98JKIkQau+YvuzYEoCQ/TX/nBbQWIQ2+jmyTasqxIxZ3Zr/4PJbbhnv6g83DzJ
4HRezHtWoU1nVl1DoDv4EJTedoyxa8Gn4/HCx9nnmO9n8q/GO3gNLdWK/GbzaZWAGLK5MRM6GTVb
F/Cw3Z5OH7f7Sm7AYKjUK9W9e8PI32rfAjGNbUyo3sgJia+hN/ziLqaXDl7WEefKRmqysVUjxs/N
v6/ucYV4+OLwTCDE6g8RLsgWh31cK+3xHt6YjgxXq3EG1DIH/DLlEl52a3odmm08wXy0EsTh2CLC
vyY5GlcBeNAaY0twEq2vdBStw8H0RX9Do6Se/RVHabyJ/EDwlSLq9Dj/xlHcRZGt9bt0MzNzJ2uC
kyGbTSiZ1bswJYRedJ6i4CPXLry3iQjOnNIY581hPn7uEveekJNuO0gin8N3R8yb2Vt2j4mdLsB1
4jnXOCPBtnDAAiS1fCOAJBRp1GCkws0pA3RKMdkhd+WGjvmuelseuXeFe2mASXsA7o4JGwuYjlnc
i3JW8bJdU5QnwXUcvB2EQ190KU/bbu1h9q7Juh1os3mSWv71WOvVevy4vaX8AcDKYoIC2TMtQpNx
DS5F4tXJHVK1k7kwhmWaeuBjsYgoUuTemYYG3T4F84Tlb+hLudnTKDudE70JDAyguiFk7JPp3KR7
zAnf0NfVlkVWpELijTeQ1KdIYNMrgSdyjf9ELviBWt+1culmA+1ftJjPbNLKRs5n0wRSTxtPG8FB
vP1qnB63AfmiQaNiIiH7tEcK50qncq52A/3JloL2iRZ2wHJnLfPXxX+J+c+0NU/OC7UUbvypEBC2
UvnRrNtQBw82Vnd6avF/4OjnKQUVTNSBQaO8UPKm5ZUF4hI5c2JNwuFvurViC9IT9NsRtlD33dn1
NO2Zh0RAEod3w7+S5o17w53YGaOdZ9EbatDninepdKHKwMkEXz8HnNy43kzk9ud1rNcx7sfd8zi8
WGBvp12ai1e33508m7IBxBqLePLhBAOAFQ+BZCXmhW1ZGJngc0xU3/POZF3UC3365s8WyBWhL2Wv
prjGPz6yDY+6PvIfdLSQHa/qVZlKm+GOCVDQMtqVybGkiemHaQWUR/60618jcCio0r+QybqCkLXb
Qe/UWTMSgoMBlJdb1FNmDqj4PlKzYwPwn4ckcqeaYRB7tB33+xNRuAFx4OgW22fbctkTy8fXeCbS
zwUKnfNOF2Q9KsnRDXImIUH/P1R9GpBAudgWNMwTAGafpWzNX3qDUgqC0wNuPD1d5aey2DYk+b65
ZFwRlMdXN81kDc999p+6iPHdtLcDqOkbxNraCjIEE+R2RzCStyzT/fihQN+YKtVDq5ot+T7pVaX3
ojpv92Imed7fADw0aiJCNJe/Q6rQiEIzfKfYzFEaDbr7zxPNJG9Q3ISStVqWremAzpJDvi+05iJ5
+nqalQ8ID7ANkcBmGD22xDINXkgAHe6qCI16YxYQZdcMHAHYOssOrgzFqgW/74XcaG0jLXe4Jlku
+eWnJbOTmWL+ZsuNmrAX02d5c2KpGPcHXFFx2mhjWp7eTKwmN+edE5ku98UEAISOU4Nk8jE5MWxI
Q4Z7OtCgmpJo7E7BUHZrbzFElP1JhlGp/92y45bRXe0xdqGa9v31wCXjfffwUFdXGGID2aF+dSFx
sbPnlQRSn95sMfAEwfXwrHUJOKh7PJsD3c/l22/InHCB+tSas9q6euxX9qn3JjSEPiZ146PvbPiz
QLD64FNJHuuZbgKMrOvagGQaMkTjF90Fh9XXWM8RcfLYQBsTRmGws6U3/8EZRZpFvPSTy1CLrOVy
oX18c8wS62ClkSP1JSE8xUHOedJHMFo2ZJt6G4UeUSex13VOnoG2Y3wDIONlTplyIGSiQIXHuCVu
YBO63pHReiPhwf65hCJK4HJL/lf4aAO5tzbsaabK2EfM/vOqce6d+/s1ryX65KykgexPX4lRnghW
H1umimlmav3g4CkqnW8qSsjua5mvzMaPfQfIBWgBxpRS8o9VsjL/gk1bTW4dkEuidnU9Xm95T74T
iOGL0S5b0ZuWWB+XcXprfxPV2sylC7mG3+M7m/YVsCXofg783jp0JjI8rY1liCewGobKvXuLY2Kd
duQtkHYYWjaqqtMBJtdmEZykcjM+bNnP6PlpLRCJOHxUUfsuM1v/ifAccNE6s6GOFqOMy/r0ENSd
pFCjvWSVOc0hVNU8rj4ltncanDkHdOUV2irtm55nMLMpBziNQlS1DI0hIZbxeXIDCSwtTYtvaOKk
6/HeTYRGC+cBK7psqOWYYFxMSxIMdfC83DpNbbs7JuVxL+i57vvEBzwCj2a57DAHsCVrt+V1arzI
3YIZUiWIv9V8fqo8lCqhzDWSlJL0cK0dG4WOPdgsgsr9aE/aOoLvFCes3I+1LHtd3gIsuLKQNPfz
lFQt+x+YlAW9yB2fEum9JWO3cyMawGHcxxkvJUEQXOU1DvvDHrGgOiDr1E8NMJ79HAfJyi/Cvkiy
fJwY7OHmrcMO7iwZnD68FrHPUB+NoLFH2K0yvHDy3MPZ7m6RWHPkZruQ5lTTMz4Jx83vyDTm1MPG
G5fTJaDR7FMHJ2tFH3hix6FLBlJt1/bTWHErAul+DjeXkI4l5ij2E58al4uVJgOarB7F459qznP4
2WE936I2cYDxMymbcfNTJq5Eq0RZ8AlehveZFWYlCI+WOlmauj+ouMD6zfY6zeHcDo9PXXpdoutF
7qKLr3plIzAUr9lJMP3WTkxLV8IYgnDhVU2HzKed2xarsJkxppdrAeHdhE9I1uOjcN4Cz9Mh7eA4
e86elGW8PDD3X54EOcQHT3jmSz25XGP/58wMfYwee5pI6Q5asC0cy019Ea5eZ0iuDPKHD0VTyfFd
XxipC8iQQKSeY13cgMeMj8ZnEF3iQ444v0KaYD42KWUAML2leL77GyupD32KXeqwkZYSiMip+98o
xHFnZLwAn+xJEZRmwqAZu30DItyPBWKQMh2TTMcT/btPGyYQ7EXmHqN0dgNqrsCEghtmfjdwf3xC
Y6vWPjLBEuvCVKBzMDa1BPy5VwKkEQt1lacA+meu9Z7KuhSmJUFvZmBIA/4YRFuTLu18lcrkk7pr
Zi6dtHfAaOch7RbHEmJJ9T/2XusL7jen6iCQy8PgwIQtrsUGNLoGQY7z+5JGise6UsQFquAxDVaI
VZE30vxNRdfryu5jd77+BK7KKZKLXGknL+eosfrW2UwH7P5x/qPgZDAyL4bTQydIactHMrjH2VKF
/84pyxhY+figuFv4MieWnc7HnZmJ7Up03AMUf1cF+nlcg/EHXlz+SEh/smVNKCWsnIhGAWtk++Q5
JiilarxDir/X9t3fJfXYZHi3t9Y7/TVoiznwj1IY/iGonYLH4xUw9/1m8gHhfK8+AHMQil4sPFWi
AM046d9kcEt6lvMixd3SU6mRyFImeuWHjltRdXJYZYfKGLeRL108Nrgd9aC1G3GjapE2yJUK2j8f
UBWcQAlEAYpcO3ZB++IVGGexT+GlP1Yh4WWxgFRVJdhZbYhEd7cku7X+c3p9oi1R5qTUIoBiZnlE
GN8UQWMQxWoxaH3C/SMfzxaCVQDk6jT+wuPPVU9TG86Fu+rog2FEZsLo/duQ7S27Nf+KPBs1BwWQ
PaNdhHudZhpUZv1Q93+1d3mRxELEHT/OCc2HemtND9NryEDMbCKf/WtQb7EUsInPyGdpgTxKP235
dvaJyij5Gpp+NtCkr2CZmMnVxCEskLldYWGITFD/LDKIaNS6Rpfid8+ajtbbSSYIhVYt+d2Qq7Wt
RejRPhAf9d65ze1G5YE/PhcDAIpvUSybMtC2AtSWWO2DBtP8kXiVmSXArYsy2zqcFHqTLV8IhJjp
wg7eGs/J9uMt0D8R4v1cpZHqTfuwpncc7/Gdj58VJNH4AMu86O3mjVQiSTfMjN9FXHQS2jcNK0t2
7JMq7Qim48M7TcvYIM6jbPCHg67QMxlkEPrcf6qVVsj+WbEPI8Qcwdz4kOQADvKyITeSDDKIMIXC
k0ZH5LfOHCtBgxjRgdjJGKczTNxbrZw6adIlW8ss2sPKCWDQ/0sCr8eFgKfi5MyRE5JtB+LEJ+vf
CNvGgrOUSQzxQQSfBmSRUtb7AzvlzWVH7EPHocoVMbXYiBnGN+7iI/+xEBv9HBAU1HKFGYUACn8x
6HMsSjZ8jX0eugk4I0kSapU3Y2/cfygKLOkl1kaeHrQzyONtfOGMTXW1lkJErhKjo6dgtUBYqrmj
DZz7agkyASqg3MyWIJ2A5fl35dOiM3O0xatBvchqrWkyFZ+d1M3fynGcFHqp7C1i5jlHEimC6I1+
kbdDjLZ7nQgoeQCSpF+iKslDpLmqyXlMfB5cbY5VFlzK1v0eKO0BtO2ICkmMOGJ9H8ZZIgNWSvCU
bjLqPb3eWniUKSf9UX1Jxx8gSN0XcteLWyRR/lLHoyFvlqHhhq5qAuqZOu94v1k6Wd1BHJekdc9+
sWBE/KfKojAwRYX89jXNE1VHpGMdvv+otmdf6yXlBoMwQdd68fhBLJ+ZZkyXeyi4TymhpS+Eodau
cQ3eyFG4jDEUx02NYI/QTgn1HmTK0up/o6K/KI0vFMkkKeeU5AWS1EumMyQyvQLyDpnYOiMPRdvW
8Q7kE3WA4Pid/4dYccfKUk7CsQOXHFB0SGkLmrvuAJFDRKVc3HGfmsYWN6lVej/RzfkRXcO56wp2
90ufHcoyeGdps23yMHIaxt6mtTN/nPfIu2wQMEQquslMdLuEUiEWgJG0RQjroC2UQ+NSoR5THXRQ
ebsvSTy3CmZm55Wkk6op5Hm2FU4bnV6sTAxGXV1pqizxcHTobr2//FDsIiUhNHQewoFm2f1DzhTH
O/BcuP8q4vuobl9ywP0XqJGM6YgiHWzWv8AAS8cd7DzYstvFVdLlJg/zzb1rlf1ltmSi+fiF0GrM
yZyx6NKp32HaRUiB99Sz3O4Gxv87FNf1dbk/hFWspRcTU/pOe6yOFC6/2iq2LEoyg41VW/ehB7tG
HeqlgwiUupPxm7RUipYz7u2J46ANwOUTuczeBACGglQ39T6GgyqeM3ldHxi5LJds5xxQzAh9suMh
WHtsjM4Ilm/LbJTw3QmeGDQIhboyCXxqR29N/JiSU6HcJy0T9PvY5itmwa22MKtSqSLYvU8HK1KL
lDiVrQBIGLOIAC3KaH+/CUJzG50p2jh6BuJHqbt2dWNqT1JupPNU2nrR9BZ+8MnrYwmlnMN5hBGH
kI5QC8lsCX5tMubCNnVtY53XQg2o7SbTcCwtUtZWz1G1lyWzOHb5M9brLrrqjERR+LI3SJOXQAqZ
TSxizGemQNIksFZJlvsDJoDamg3hAtpeHLckWiiMAUja8yAB3vly3PAnDbSE/dRQ2KuUiwTrifHu
sMyP0T8hcxqBFSmr+dzRGetRq/mjdN5+nm6U+LJZThm3onZLAzu2UhdoiFZ+tSMetg9IgJk0n4o6
69xmEihMPs3A/5PHIkO39nyUBJ6O2qdhNJjXABvkBoua7SQpI3dE1VgyKYz8kL3XaR7CY4hAh9a7
s91DL5U8K+7jS/HxVarfulh9gUVC1zhR9NLKwpp13tW5W4nUX+IzU89/+egc1H54iKsKgSsXLSYD
943lTORuwTbTDu3TXcwino2eMymq0dHaGnIth1jSNF8zoy9kgS1pvG5FiVZsIu4wHjLDJnveuS8h
+L7rKQje0Ypx2qg5RVSeTjF4blEyVQ50DTlG5z4ME6gWABKQ4bNq2UiWftnEwB+WbpEZXqQGBCvR
mhcm5ZsBghxpn+y0U9E4XwXDhxpFVSV8dWODg38QGhVZKMF78/O5lc6OifIuMA4HDagQtO9ui7k/
Q2tHmCGMyOlNvladHXS40FGi6LGLH6mVUAUE+j7dl44H4ssr8ZIzPx4kvFyfIRR2u2sTQg6envVm
mYvvCHpaEsnlQtx44Z7WHz4GwDb7qTkLuLOLvZk0s8wwYByAdLeezs2NhrNAY4XStoTshmP1yUWb
zI1JXd+1ZswJFY+KF/f4LwK+jEKp3MiF8TKpkQoNiVmodmQgnJR+oJnQNDGyj1X2JTY55HBLnfum
+gtmNKBPzalBKkcAdhWqj0MDhtC80n3ejuoNo9WIUW/GWG3Dw/wnFudw+kTe18D/YkqzZeVZD3UL
LNgHdNadudbopVH7F0T6SFCEf+RfiuO5DjEbxQO2EzhIQZAyL6ab42MqGzySnKrHvBe/d74cGVSg
uD4Twhwq3bGb2bL7D3oC1ICM3AXDgF5BXjgrrnC8TSU0+OrLMjqFzRfHTvTkXNQpPpfNHxKjcNTu
Dhm6/zaEPd6NgwaCcDIqlhutFaEe0AphOXVPerGQVPrgGBHbeb8ryJGMXBdNARCKV7clWi/nywKI
VO9pCqaOpi7jtoKI0YkGa1RUWEdj6xawQPrxNjB4ALgH7iFxilxC7BpYWrEo0JScLM6jOLVWJbba
kAGP4esTzLYZIh8HFrbZrXeKL9U0ccrzxJecqfUeXosUoq1KX+Kk32xec0cKlZHA3nhmwfE4cjci
X0JaAhpUaWAxnb7AZsWvDAE2vNq09d2YWNrlDMEqAM11V8MnJChxRpSSFTBTIW7Rc06O2pEqU94t
t3DicisWHrheDdLiLmWH1QH9H2zdaqL0bDIOyNIrjB3Pb097JKfZfice39uheOIBky1CFvoOYMpR
b42qeB6tY0Z8S4PlqP6mCUm53z6z9qdVgtZy2fmojrOnABD0fbyZTV5g4hFg6bnkEe0icA9/EcS3
nQytAmGflPubL3GSAe+uhq6wOZQgVmsXJx0CM52M3WF0W0jsaPNiiCm+OFdXSGfQ9X+XfAjJFwrN
2K1xSdF4Fe2aNrHdalEtjvKUCp76QttnlFUnseEfuERlUissZ417q4WjkzBI7C6cACLioiILrUvC
bltlKyQNwkggHmpnfHyRru8KGC87rkIVQD8po3Osch1SMzoJjC8K/0aNZ5ZjcBJjO/QNL+QrDpT/
G2XE73pSASfvyhfPEfdwgxbRFKagc/mKK1XTYuUz5/O/+AeB549Xf5qamiouNu1OnG+WvXWwZJqx
xUIizmgv4R7O80fLitKw9+Ixj69CBndccgWAo8UOeAp+5CNA7O3R/ADEGdY8GeQO4P33sZH6zP4k
U5nT03kAvp+1PNzebYKpvMstm1AYoo2jWBPnakUtt7L+b9E4ho8JQKsLZK7g8kiyX8W0eiull2qf
0rTb7D35xePOaOkh7BAX40uVz2IWApMI0TO/l8SmxrHngndgND2stu77JJhXrtn0cSmbLDxFBxt3
WqrlSdz8dAA8/M1KxX471Vg6bqaBum8TaTzA9Al20cFL4TJFpY+V6ontkGrBkqEE5qpTMF6zZ1rw
3rZdHmsWqBNyBUS9/V7vxDvEqE9XUvvNm6FQ1dyw/GA8ve5eBQTl3Lxa3R2xaTQzaw5KYlk+0kma
xNteAZ3yWWTOtrRlDXbSV9pH5381tgVnUKRPpRLErjkC/0xmYaixyQXmnQi3YdbJuYgo6/HfK19K
C2cVFXdry64InCUUeYOaWFCCVvNz42uX8Snvl4Z/SIKIKNSJDI4SMHUWadt0w2VGSybySCYplj6P
jHZVVV7dBumUvV9QJCC7Mvpn7Xp176S0E9vkZLz0/FF/xZ3GSQYdhMLRy2uet9iMy48JMb7e6bfc
ZAKmAmeVixt2Fahrvo7NGfZYUKDkaMNUkd1jHnB9QbdAn0Ifxv7pNmQVpKGIwTOXUYyL4j/TRhVB
qk6XJlqGZsvwhHlaetl7pr146Fry8ZCAJjXG3RMkV9uyznWPmefLvhtNmauqOHeIQM+7pdInp74K
2nENUHErLOJ66dFMnMCdgbHPIjnoYgyeQMoX0cH5oFIbe0BxHrjCFFT0t83YHTaGJV8G8M83R1fO
Iy5CSdWkT+9c2J12U7yQh+QArM90tvtc3NesvSgDVF6OvOpL8VTX1M1rdzNbIi4dl6a2Nuzr9p6H
OyM2Q1sNHY+Z7QBnKRY+L9XbYcnRjIcYJntIPNWZVpVKj3PWQmovyP3v9Savh5FrKGH8CwmiH32w
OiXKhHyYlgds1+tw2UlzQxRe28O07hOKjUWSFIomuLnyO0RJFCPbBplA0l6YWnOB3MkUUu2w8L/t
zPGkp9hLgLwC6ueSxGxOfbaZvJTl+kwt+7jMbP97fw7ytYRJ0TAZVuHry7x4CePmJ+tFNgKHpyFJ
yYVlfmMqbVd7tkFkWV5IdXLv7IH5sFQz95oosvHfTzixc+GxNEx9UT6fpert3X24TrqdXdcPSkXA
gSGJILVZugZmRwZMMMvsZyKLysBE4MnrFoVgSn+zDxVYYkqvSfjnvPW4TlZA+nqi7H7dFxFZuGWX
SSdyDbx6rGB7mTu4RwkrHZ0OlGAJUViyfrrWmZ7LffGdN9nEn5v7kC9KocRb/YrXS7uFB/VBE0Kg
O8GSLYWn9BVzwFKmLoLrj8SWSE8o0K85qKr409+Da2Z/p0ogXwk1z7P3E9ud4EFcaskrgcbnPuP7
nhIUpDexmfK8Q3WlF3G6oFNKMWvD6AXd3TQQXPrD481Oi/ErP6I6QWc+K3l8J6a3AcuPg8eCIdP+
NFOJVBsPGXr42jMd26oN8ZzrEkgM3y4lHcARJtWOLK8eQK0M+xtWIz6N9YZFpuiLrHJqlglUSFQ0
rLfefP8xgXfhPxAMs51jdvywiadyDIODvRfhIbuX7BIWgK7QRrfZg91BMrQhIeglxokjdcYLS3SF
El5rwcswqixwE7Bmjrjl2S/YPkXp/qvdEPnTbz1tC4Td82CPg1rPFx12V9lB3gy5fNVu54NynDDd
WBtfSlali7TMxDYt95csS0dx7LjeWZg5D9K5G8oo02ACtkyuh67KgdtTx9SX2zHWzLN+KMjOob5W
+7J0W0SBNBwPGQkNWzjjEhz44np1trrzHE/QmmNj6FvT9sdeN08LC6EoBA3DcCdGwDS6lG2FZkum
vE1T0w5oh+sd+ID4M3uDHvqXssFnc2Y7z9fVxDY1ymgS2jTTRBm9cqIDV6TuVU3SW+c44HyBfBu/
/5ib/g9zAqbFq/+AERmJboM1T4Tid3gOTHisLnUA8ZxSIazehG+P1JU3bQotqsBduVV0w3O+o6TX
mZgbiprewEpTauU/UyZxeaIX79WQSw2fxwntYf+c6ITV12d9/LG/DgSHtRV1AJtt82D0bOcB0jvh
Qso2M89Ei0QpnzmtaMC6CdJ6GlZg3AKj0NhBFf56Ip8e760024aUEiNpISmTsEpMnp5AZHGxHyke
rb8gEVp5i8VbubGH/wMZHm5o8blkWLvZktQDuYUn+agxAgZClGWM8o0+zk9K+F4HXMCRZwX8VyJ7
WT/LHP6W33tGsxb2Jns324QbtJ4pFBYwtTb3VHy5CKPxLFPLMG50a4j1H3m2MY2T5L0KFkUq9pVO
/qokCP0+oLrMXD72g1wG/78qsN74EUQ5Wi47tELxVTbWmnw4akTkMPdcMM3CMkIKdBpgaM+/45ob
+JLQxwUac64393mc+kpxPi3RYLxGkolsuB3QDOfI3B8a7tAhSN+h3Foq99sLYKB6O6ZhT2VkZvJq
uF0+AXpKV9f0gGceLEmYHKIkY6bVSfTrmeeUo6c/3/Jve11jDNUwCnBINva8JsYER6ARVlJ5EmUk
3rSXsqnmUFkgABZBmCjWUTqUGJMbzmLfMbtT5QYPHsrFsIscLOb3pFlPmVZbxXK/crOUfG0TEmyV
zEJtziudVnUAV/vWzKRSoCnE8ErIKpkhpj68Q1AsVplCo182Ferb8O2vNj2txLMKUs7YsCoWk1WZ
BxORZRfnaXqF2ywRiHGp1Pp82fsIQo0inTYjGjF6FT+3mwaEF6OFDaUH3dNtpiqeUKcq/sI6bfZ8
t5+v1nNVaGSJSU287DUFaweZ8+nQia2IpX/FgDt6ggImnSWdnVmtomlPb4GbR7B2FqtxOJ/WZWyr
ordnGoYFLRHa9DxAfdm57r44QOpaYP/jxC7wtg32T0rdpfYz1iVmmoovc6szLuE6dA2e/1it9onK
pUw4l7hkVnQ6UwmEMPhF6WBAAsW9nJZS56g5AAb6c0yynVgAUqKec+rMp4iX1hW33hxGn8DrSXLV
6rwXUVZNdX83cCd1aglgMPogiYXawRCVEhpRC7NFw2Hur/ZKVHqJeQG6AXQwN/kuwsdujptgG8sD
nliT05F4AlNmpk2wXAKSFqW/v/xmUvp7rCScIaEPhn5vphTlnm3zSz7QQ/AdBOHMfn9SE5TSQ8k/
13qUx9A606XnYkH7DZSkAp56FC8HzKtwTJHUEYk/GDR31MgT/It0bPLgLmamaDa/d/6T6hlyh/uN
IOOlCpoQhaIKRJP/98r7kgqEdDURHlrqrq+Rk+e5yzFuosflw3KFeAnSLZdIMbKypAKyPLza6jFp
tSnRWwD+/8/8xHzyu16uHnken4Vk5JLigldTmnmlxPUeqZNg0jCs5touUgxne67+W18UpYjPuroH
p+BoJDiO1NAcy1+9lIbIPPJc/EwmPQrQhgQOw7hMuUco24GeSF3ng6F1RVRRqqd5vw1J4Qtt/e3g
cMHWvnPHLpSSFfAamcsHGOk69azlS3VdiTNBUr8q6Zn0SpoEnJZK1M19gibBUCB7VmuW9bWuvhvh
Zg+At5QhksUukzG3Uvr4z/LbetsrLbqnco/vgtbtJrqv5HHITPOiEL4NcutW4v5AZZZ+GRydPVQ/
NvTAHjIP3QyZ1nxtAS5DusIn9SFDnzD9KDSbcYm/xv5aussI8HJ3baWkGcsn3L5hzvl988nf+Ti+
rKh9IZ8F6RaVDIaCrSAQV/MfE8PU/kqkp+1XfWPt8qV2s4ai93rwHzeOpsx1YqYcDTbnM1QZhzWc
d97j+s4frGygk/hUwdikfhFYE75AWkpn0uh7GNRLOz8aKoMYqhaHc5ofkerWBsvCFmb7uNCkLT81
dTmrhPffHm3Vr1uT5l79SpGEjq3bgm/XAyhGkrnR/XsiI3ltJpTuKD51O0KSZzIzcKVoFlnod3yy
6qOZ8Y8TiFHbrtceEhriEFcmWb+8aWG88pezZ33bU0SpRgxb5uoAE+lFbwN8hpauBmgdXFz1ZvMJ
mnMO0OfKlbtlkW4g+K+Cqygz1rJaaQGJ0BW2mV417BQfilz6VhiXVnDfuRA7LyIcA1CtrTWIZJRB
k95Yojwr6IuFZYOG4AsWeMxOwZXJc+qMs/LuYI7NNd+meFYgdh6VmSJQrRK3A6NXnNEQTxiW0HvJ
u8+YHbjDnZ5qrXFCjmvs/oTJ6zCdwZgZKLkXtm9DsFzlcJpkN7tMHeTl1FhZ+eNWGngF0EbGTAtJ
rA6hSCZziPt1aqE9szKmRfFpWX4K6gI9ZWE+COXqQprGVevoTSUY+jiTa+T2bs6UsRlJ5bcFLnGZ
S14Jcwfi3zm61bj/VejcXFDakVH1XFXbn/mVn7t90aYPPrsu9mPrbMxdE35UbYmQ08XSX5J1FHH3
jalk4rqIVBuyo6zqx/RYz7S8gLuDbuPQycz/3Aa45TnXzoAxTg5sxRNVaObWoE0GGDS0mKcEkar5
8T98BIhp3zF8PCbKwMhfjP64rIvgiy8wCkl+3/MxG3iwJEXRUzlWrAjYylXPWA0jvqeLsQfyycdJ
KHkBtwo3NxB0DiRhfJw9LuQ/DnMgAP6XLuxla2yEAJKRyDKIJdf9BT7hSo0ZnywF4DcZX0yLe3m9
1rWx4Nq4P7OcSlfaqKTFRxU+5oIQ+U8SiaVaRagiJMvvl/wX/pASBa5QL8v7wALoHYPLBt8Zbpuf
k2McszskfPysy4ZLltuzzuXTsoLgqMeSQp+WmydPxYnFkmzsGXZ2sxjUaKMRQ4vSRabuThhSZIOF
VMHrmXVqaZJT3BCOU7X3WnAlao3bcbUfUPZF5xtieUm//TzOP4TC6dyC3Zyo1OPj3BQnd+smwTwI
uhGisM5nMJU+dAJbBIZ2Y3ehUN/nyJJ/KqK+NycYwHol8+zWMicTObUTJJTo3BpmbdbgC79fv+NQ
qmO8H05rtcZjR+oA1dNeciA7MvZFKNb6NSLLoEghyVCTW6VRDqIEHbhbrkPutijYQUBqEH17+jJ+
0TcxBiySEbdM5KZagCZHjhpeHFEdeJHyu30HYuLwPKTI8w4Nl2eXfReklXTFrKBr63AiiGsutJCG
eqFtA9OWt2UkBad/b2Cb/f+jUrfKyxLedptlxjwUiCpycWoILHfQeNWw9VpMkpw/gJ54qKaw1u2Q
nZm5bbdiq29XgWoeWEFrz+npMfHE+J1s/84qfb22sh151dV3QuebnGG3b2rz4KtfLhd80tmgdHgZ
WDZ2jd9VnKA+5bMMFysGxW2q9lysWsUAoZAsYdx6iEWO/31nuJ7p0gVnMtvSAhYAnD/mtQT4U89T
GtsLkPy8bwCBq+nhC9VuYiErYLsuzr4fn4rLubqa1S8eCJFCEKPbLpD+6iu9i9F+y25CfK52VZua
CZOKcP1JxYV6hWV08SP0w0nokQ+nZrgiT8bq6gV+qNI1oNlSzKPLc9Ycmbl4EVzu4OiS/DbQFKBc
hB5AE2GReXmkbJ4151LBJTwQZ1ZHeJ5+cqEoMkStaG9Ay0yK0qpE4B5k6S6bjXqaRTlFiYTbCIjM
yIyQQA+igO93NdViYgfS2D1XSRWNHycYKuxeh49OBMzLLWkw6+/wbrvpJpQczN7KGmFfrwvufKVg
/cMrjJeH9+6Biu6WsXasacQ8CdC5QPb+f/4REyWDNC1rGmnFwIiWrSd1eEEi6HtqgylipLaAFwKY
S+hrVLKLThwdfyUNv6kK0FYFiMlcNBWUtsW1UwnfQJbxOXsv4W8NmKd9hVaPpJbSuC9P/r4mRpRw
5i9f7MMPw2unBb1EGd64Tp1YUDEQrg3pCzv1u6INOGHt+oeEqMPmE8KztsSNqieLiubGP5gjEKZM
V9b2yQUVE5/WQvGsTBIgoOWqhhZhhiJV3ZMaEvWL+ZxYxuWadbfhOvAzdpjXXTFwiARTlZ1oBqCr
3yqhNIAYjYylTGq3tfQHQ16tt5WM1O9ShFMVwczwOFYoIxy6481pfrHYWy9YEAOENpRTh+HCfG9q
yA8fHitIDBVYPybg1AKg7Qp4tSSMbp1dqYSlz7uPl+bJQupDXUPJT+vTSYBJfx/DfaJPMDUcavyv
31s0BhIXXzJG+X83E/tj8GKvSHms1xim7YSf/UuOjI6YmgaMeOTCeDJdBE4pzPPDIYL86m1y4zuV
anJRrJu/Iu64nm0NFY195ujdbvk5FS5AjmxhfEhWjEbav4aAFN8KT5lP2j9+7JM0qawsJsiOvi4Y
NdJ95IR2vtV3I6DVvB9RgfRTsLPmmcmMIqWqHqfjRPyBUPMYnGBIOzDKHETdpdif1o+VBGXAhlPR
jhGV4zT8/RMLtG6H7TuEEg9Lm/kO/JnE/3kduQwSZQqXG5W5lfk7r3eAcYFWuEj1JqHxjOH4Rmtg
US5YmsCv6tqhv7RQZEt4qd8ISsi61yT/1e9mGQ5Un8dZGV1AT6/rhIhiWmxfsfeDHcPOge7Dixyl
HiwV3I/UENm3Ev+YsWGQ04pqIbo25I9k6SB7sKHP+q6k4IcuJEIg/z5eGgRqyirMgtyCb5WCwSGt
O++CjfDsbFP9+DSJRIdJoPQbg/zG2jPGi6ICafUSs162W1k9qFfHmwp8DZQMQVpEnGYGKNJZna8H
WgG3z+gz+xJ4dIrp8j8kJy5eYfNfdOy/vKoQIF8RqpdWSHs6SfY5TNXGv8I7X0nAJbjojajqciEl
KGIBypK1YKcGrv3b4YUgNK+sS0CEP8NmxjywWYjaCjWR6lP44pIIcJgPaNGz4l6KB7FlcW/10sGK
T5ccpdWwPrlosSMa4UpL6eywpIfRRNM/tK2awMgphHs63RKD2x/Nz6qni8vwWIOLYCYYI6ndJnmL
DYnHsMrsC9jmSIBlGjd6345uLrjQTw6YyIT7e4GllQb2qsH41QGTJOzAjS0Tf048uq7FqI7LX7Xi
Vw+xsdvOdI4qXOBJ8LYttL7BG3NdJcq83MxcOAMMWTQC1wEdO/jg0DdEnn2TXqi1kH8fdl1gsqDH
Jc8kN+fTYAa5Xt8VA2FtLLLIsX82OxpdpJ9FEMTWokQwhPpv1MuJ5oDKFwt2T8uiTkiGIjmQUt5j
g4FKiroS2GWqjvSkeeWgNsvHjR3xifrCCFNug3IzKItui4529KGTLq7iBeZ0T3WN0WP9tVm8rFgh
SknH3p95oiHSatk5GyVbRACyylFRoSlZSG9GXTXS28N1+J+plQasiJUH4OfB+M2u5e1HrjwmDTz0
8/mjkmY/9QCHaqQEMY3wFtzdZSN5+b+jLdbwtgzffL1nf9hsovQX+eV2Dn+SvIamaC/X67j/SUYS
rgqwdTPf8BhCfhfHK7Rh1uJ9JwxlCYI16IxcfOxgqIl/t5BsCW6KuVvzsJfAb7xvzKa5XysN23+S
d/KiouHbCNGk9ITSpDh8PyDScgnGGXACm9YAc1KFkKPd/ZzVZXnsE445b7biolSat472hAzHffpe
+9iLrLZ33JixsS+zEA57fbeB6T6qohWJKBS6iuNIY93wDoaU9C/82a5H+qbdOZM+z83fxnyG2A8B
lDfHBNnYCmgIgJmCA/kJu78YUcGTb69U2XNLf8ha2Hy5YbrUar5k52vVlXKjECa8wNko98d9Tz52
RQW/xTLf78juplAA30ru+FRZBSBccQLnYAC1nuYAUhTg5I9k0R9EK+wh9FVJSVCMWhp1wAzLexKx
FsYiThoGYBNDdVFkVbGvEX8P6SVXmXcq8lLw2xBw5RByrOELkRwH0LmtokgfPCCz8Ja/1iucmCpa
Rm7IOBuSxEhmeRhIRenuJG2zNaP//QEvMxxt6MCuCLHsVkU0BaO7RqPi7BnH/dVFwexhNAL9QZuC
EpN1OCHzTIrvTT2HZE+ayQh9bUdtY3OVSzOUFPVqMhHuJa5jYw3FULNFiQhKZTuztP4W4J2WYaAP
Pj8CZmHncok3ouMUuTq9C/R4peYYJK+i2y/Xsvb0cATh/T29Y5DPqyLImR7OF4FhkadcCAkAUUfk
geT559RDCAi1oTedL3ryTX+t130AKG724J56Wod/TSuuMtoPK6syjE0tnhJKl6NUfgh8YIiMDOjW
15iZIV8xJ/O+fDYobxsac1PffUCHaxfm617BTuGfJybGSHwghpOS0it7pvDySD1gFMFWzkn+EWBG
3WlNIAzwM9jjjGkx5b8/Kq708us5ZPiyOdgJn018WXg9LzAq4IS7E6o1G747R5084jiXmAO6dHI8
uYrv1q5aAbJs4vaJMW4zddhifmBX9UAYjcd4fO/GOA+GxsbA/Na6ZwkFAQQm3YI3UyIYV8kguMbO
aRMN+ie/7nNq4RLsFnI309KlqAnCoTQUQq1OsE1iVMliUbSPh/cY1eH2ctv/HtkLRGi/GdcxR+z5
uMWzeam3gCv45BbxUGcwrpL+0WEWsC8NI+WnMOSyAvwOQO+XJXRMk6Mrrk+VtErfEKKFPiRZQnY6
dm/foXiIb8HqQxFK2qICWraVxdxAY4b7xILw7JgbKtmQtPjIUUwAtetYND9qJ1gqXFIxMp1pduSN
2QG6dzbqY2ko24Okg8OZEtA0LKqeGqMZgwgHS9s9RFNUEFWrPrgZFvzomNmbvZPJWfp4fKdCkV74
/xzftWmJYEIfSLDpv+yo5iVtFvcXGVVSTqSTNd5GLms73++b1K9eMOqS5WrRjQZMWh7nZy8VCCVp
nxSrz50UPDBQcaEEHQgcR8cLmAlSkopUAUp/Xi1Qdx2m2s80M5qEnRZGJpT7wSJ4ldO+Rx5jR4pj
yIUkOjwlZJ8WdhxI/vl27EM2yCmdeLm8toS+dt93v6ZA0EOTCAMl59d1xZUsf/GWbRlzQ2w29dVy
SeCHD6qGrc8WEpdfxrRGdtgCsmh8G35mYm2R7yKHM1NigGeeG5VKSo6kQsM5noye04uA37bQkCgW
9M8G0FMYI1UPOPy5QR9h/qiLz1680QpcH3Ln8ozWqDwK2LNoSvNcfrNPrqcI6g4PRWXsB3r8RCSR
ZCna967F0yy/CBpi5dan0bE2hVsLOBIfE+JnaSmddA/gI0vXjST3S5EZy5aRTDJlWYo2LyChNT7o
pYGKyJh04HbKFZAv9bUpJhCvcagu+PbGNUleOJ20EraIPIAruZ0lrKNZqaqvC1IAkmB88CxZ0Q4z
27JjnXAcD4KTvOes1Rid5GUrTngpTvqV35VHKqn60yvvkJvgDu57545Tkm2GJ4KsWqsAW7Tg16QO
PaP6EqJzQEymAjUeP3Jrn5aWfSeJtDeL6bjOsi4iwZ8GFt5EW2f8WflKj5cclij9mFkqaex5Z4ym
CvfsJ/BE8WSXOvypSzNUaIfpDzeUkGMcpnXHVWXBFRgYPtPkf5KP6mdps/U8gFnDJMvpQnU0tOvi
UorLWGal6FR7f4EN9cAjwiTZCY5B0qKhqknabLhChDb3oBXMHfprYgZuWQNdHlLBon5Tu1lTPIlD
ECeN6RaU1O/TZTiD7+bPILSeZ5xAQNefbJS9xy91/cNEcMbSg3t7v9WoUf1B551WRouN4FwSk4ot
xFLS1M2r58LrILfMRwq9Syzkdflr8YYB7huBkEJKt22lxZhz+8k4PPQCiLRCpKKVhTeO0Bdx79Ps
fGK84ZX3DMlk/zbYS9bKY9WOc1diVx7OMJInuLhe4x4oI3Yy7GzE+1/ODxKMvFS+wCLZ65eFu1+l
cmP4tAr9q1rBtBYdfpsmKT3hylcdZWFnYWb6RmzmGVBPYvE89osusBw7W9J5rxRWLJRZZhwZDdls
l/mwiA071Ahe7EDd6SkqvEBbuFbQzrRUqj48aDdBR6H1cMVdr4u0kXmZGv0v3Cl/Hc92UObBEu+G
E1Fk+zbEWECQ9717yKzkhG79MIeAEZh3YAJYX/K2iuF7fk7VuyYqnMAetkNKRmnxL+oMoBwb2ul5
GxOjmlpFN96Eup+xwZFLLpAV6Gn3dmDan5RVMkT+589q8zWqIdsxh32PqmCUgnqSs6RNAkJAIvBX
mi522W8+UjQpgQ9qcICwOpB0oKs8R6yTH5E2T80yp8jQerjzEZ14ZwySl4FMMAPYOjD7hIKLsY5c
ckL0whyZccAzgYBxR4d9VUkmHXWnoT8KgrIF3xw+Y4ivii4njvKwn3sr/Zs0Vq39G9P0Q/stRXDF
FlkDAQugTsrqZcKZ693zW6wt+BHysJSHzmzRnr48nWQD9q/qgmdFv0aALAYVTgcAI6CLVlKD0h2w
NgXWjX0abuq68MN3e1xS7hqt/Z1BNsDQk482Sr/s+nnwCd3xcw97c0Jth1BSRFcVjuVAefoRE9n9
MeubjmkGwSkWpADRjZLby6qDREHW8zuUwOfVCxbNynrDKHPY/BLaYjHsPkzIRIDAsqFRdmlyKW/U
+UCyJD0ce/01NLNO7HDlUXZDRGdt70IqAqg38GfYUIBtssdRn1W7wgDiRp1Krrr4GIRS63MZOjlv
ETWmqsMGS4lSmPz6gowA6nbXlADuXV/PUy7NSWdk55W27jF4VKOuLyghvuK1VuztPE1IDIow7cFi
SI0JXCOknSGt+hdDr1O7rTY7D8pNVBrjD5mjg84Bu8MAeREMormGBQX8iyqM7iXfgB9IsDyVm+VG
kDID9KcjXO59fjVNFpbsip9nnRbTKCPeYSZhRUI3OIzZypryEhpYoi9nQnYBruGX/zE8GMRS62kL
l9UdzxaPVN7al+yKabXfK/1QoqMauOZNSFxwYdgfs1tNSL2YtVGwEgZA/xoYDUgrhG/A3VxvaNMg
Js9H1P96Coo02KL2cWEI0Cb0x6z6FPoxQoopE7StWebOI62kr+w53ClIMRxWsw+OQB3L4zPXsIaj
wEZ8rIogdEmRO6FKPWsI/I+G8tq65wUCXM3flah7/H/9c9XT7KyBBgGaLNwU9Qo7/dkvQmbKnXMG
ZDhVO09mWIK6JI1xq7hdU4YD8kjJrDA8bvcpG4cAMSEivLywKzAgYoisCk6ExHQqRiANTWpmTgak
nkC8QfMR+IC3LEx9+kDPY6hOZ4Z4HPN949CZ8SfJ5SefE5CQmxxsTIpFNA4esOlC+4/s0VBeyIMb
Na8K+P8g1iy7rKonT7jJhuYF+PpfgjhP2R8RG24DLX2dI6FF54cumdfyWCD8jqGZR4hREHtwJ/2M
4bp5vG4wiEoVhibjyFBL6Esb5cyOp4n2O3oYMusrCM2iSFrwgwVdylgXZmkznh2MEWURaMV5BcVi
a2J0rpfGvzdCTFUf5W/jpIqkMOgWUSSzSa96MS7fHQN9SZMufU8bGacwQTjM/KKFx5wATaSnUQTx
oFNhY1QXuZXLcOrSdeWUf0U3+KBLpw+cxmvcCe5KXMmVXgUcKnWOI7FCUZWstCSEfDCRBIC+upYk
p2ASaG9Gh+vAYPy8wOSGsptokjh5EBq72GzkQuUp846ooLcj66em3qM+RaxLpqKeEokM9iFBiLmF
H+SjrTFqym3mxMvyZCZM1icI30YVwcpPkaX62bjEV1bocUrkUZfprjeNRlwtPASReZBxiNWhuL2a
71K/pjqLW9Izote8wCUjT/gPMv8vyx1jh2rxt1ciO+9AEmU26kq07SU0i914Wgm1gScPFk4TTQta
GHo4WYnAFqWUdYOwOvHBSG9FqqJvjZJRXGoHjBIixir+Hv9x70kDMIg+yKm/0uL7m7qeo4xZP/CD
LdxT7xN2dWH342SK7XlHZPfozGTrF69cKN9PhskPqGVidZiSaRfsqziWZ0ZmayREy9WHjj0Bzp9H
rWbYv1Ea4BbuBn9ei6aVtaTWaAgW6Q2cTd1WX4M7+JxwVsYfA/mabwinmsWekzdZX1L5bVobP8ap
q+4Ix6Q9bxnF27WywWTJePWlXjRTDp4oyL/DxprgcRzgEVpjUzj9hwayn+6hJ6kCmn7fLJip/wDc
fJg+UBUa5wS9qNK2q93iJ0oqmnFvC7PuzTRi4D/V7b1GoXJWQyt7fidJaM58KhEmAMR5OBWVx/Yc
GvCXudW42/NbvSV+gi2RIU/9aji7tT1JWkE9Fa/MH6uwbOmnuEmMAwxO8Ad2d3Xlo3qe1TiGrREZ
DL23NL8hAcjdGLYUyES56nd3l2aeZ+kyOOa/XZ45ZgB2VcXFuXkqPGhlBw2mFDR/Ti8G1wz7FyT1
v5VneubyWae8RqJee6ThsOwQiDbOw/0RLOfLdI3zsOmVvP5mJJC34JLPfMQhnEb1tcG55gj7xBMP
RsjbbNCb9V4njBE5RU1+qseAwKHYMw7caZnsXUmQdTCVcIiGDuejG0CRucTMUjzYXbV+zXr9rzgA
vx1omMjZ9M+RDb5r6TPhuw+AvNbHwLQcdbAawn5xEZAuKfwa97sFOU1KLMdqPbmAMA8msPb3ez+i
xQrexhMbyBVHRSliBrC8XUiB/ms+AK3Onr0vbAxMj59mf17YfwxiJg41DkPavnfMveDFWC71OCFa
ajtrUd4H32bq7wdR28EVTaifKABOFJaw4t/D+JlfA5lbo8cAZhUHmDja7Pui4QWyQYs1cuveUPPC
NzwdbJQ8EPrHk4cyYaGzSk8SVoygFMEE7Qr8D86mUwNVpq8H9Zds5oRFjqXts/hVcDtvq/SmUqS/
w/4MS+YJm739mr+2T0Xi7sw78AfnwzQzXkbtuSTlqgH7RjEKdWrniVjrGaelUAwO1iCQcb6VM9eS
2fEnmTW6f/eUmbjNTrAx/ZFB9ktH3NFzO2bJjqjWF9f1bGbilK1vbAG+DDLCXabvdv1LjuK8J/wx
yMcKwKoTYt1Xok3Y3+UM6xm8LdvmFhK7v+hyqZBNLYfaFlVW0TJK1PdJTXuWUDN0wmuqR+MgXUEx
8G8N60PPsB00U9vg4WANmPrOqnReUaAJx17Lo9X/Knd2jdjt2X4VHy8NZGpjOHLbO9kMCcfVOrZe
jizBK6FTPDVZLZ2V9ThZziHEzVtIjPUfw06hJx9oKEaqMexuKdwZmRyYIhChGmTCZK4MC61PfUbM
CrOj+/pdBtZWarsDC9q33MPmvTqwfinxaU5QM5wDlfFCCYw273Yy+6gUi2N3aW8uTmutZvDEyCgt
KIMyHs0PtuBNxIY8JLkPJBFl1LkeHkJHZSNdGXG8IaPSX1I79ydNfuhQ5vvG8pZChTcUfMpqLhjS
BwbqYg/U0+wascsUYnhNfr7h4/bpAmwQa/PFJjBh+iMhRJ3QdFUGwXA5zU89Vg/OOUL8UzxJCO4v
PjmvBYaKnq7zwnuA/8onHQd7ZGJiEKS036fCinEP6ZpMmB2ywBOkAdYLImh7HT+cHWPj2N54Vxth
26vYkRE9udtEYpjfUzDcM+JK9yziRdpwjHq8+E3OiltvZcGKtyOkwgqwFzdwT1Yy+UELZ9KYrkST
fVaOd8KCcaemHOW89ntTTW9cVT3JYfMV3F9HNolbqsOH6SnQ3zVy0zBTDs66i/jKH/CIDID/9QXF
mqGujZTin75OjAJg3F9ZE3J+qcO8mAMohYJnCKcRLCsajL1kgzOscPtm3HAkRvEoTG+cmJxmjQZP
ntl0cNSRKQchxglkEzEU33TknVdyWADx4aBpcYqDGrEf6FaiR1xILh9VVTioM0DgfQwHhwXiyF7c
LptKIv2CYIIOCTzI4chKqVTmax+WZ37esmz70a96Gmjav8m3DZrPiMcVuajbK/KAkm0lA9RuOQ1D
MVaf54FhLNQqZeaNNMYaCpnUYIE1QvH4EZVVCTvHvOdNzK1DsHjVbAK3URs1HAwYHpxj755B64xU
/Aw0vAwxPh1pyUwTnaeXTwTv+Rh/u4MXAEMW04cLuh9exhHohG5t4RzIDeITda/SVGyg4bPS+lDQ
5m7WDj5sVPcBQOHVOYmTvZAPJEgYDy2qEbhmgQJQ8prsjoq6NCDmtUzSj1uw8Ujzd2TxtyfvWDpI
v7mHyMAfT84R9EUt1NOcqHfc0m38YuYoP6m8DskH3REHe+Gowol0VwDdVn7M11mdZAFgGl0sXv1Q
N1ZlV8cWxGkb7FJ21OR3yjMjegSbK+/UZaKDblLi1HzpTmfkW6ZcTjrpyivSK7jKYgwmXeFP4NtE
n0TpcN1JcGYV4G9a6M8eTKtnQFOeDcVmbK8NacnpfaGo0gyLbwz5/rRpQAJy2g2NVYfpypmcAZSk
EUQQLeZY2twWPmDKbrRZ7Ey8l95N3WzfXkHjsCdgzlAA8zFVTDPmaE3ULldzI0NAIx8pP4yfkUS+
cPqJna0sPX1S03+v+1ntBnf4q+jBrqFbBWrd++P5nhIKPR/dG9Qf4xFJLL/tUKc5wiphxfAPuBPq
3YPUdvOI/VgqQhOsQkbOQ3HYlc0a22OJzjjzeHRuC36MT9oBIQIg8fUTeM1vX7L5p+GfrTf4JmF4
q36qacbsFucu6r+R2UGhm0Z/z7U+jcj5afh2f6+KjyJBiZsJB7DQgz7SzpjC8hXyJd63ekQNlQI5
Kpo2wJUjFtJQJPAqZW2UbacRDLJponXyfu2/WlA+zusWTlli/+ve06k5ObKC5/qGHPKVzMfolwnZ
s9G03W0Cm0RsemBLyIRVvyphcUXHl6uoUlVzJAyMIbmnWwPY311FQCSQ8LlqnSKFMBMxc4QvUtMc
ubZNYNB+VIMaxvW415I3us+G9FLM+HkOdKb7i6NZbQoWkUd1ttPtGzZIgK9q1knpdGbh3HpknvtQ
2qxGaxojeakyYs/zWZ50sl5mU/oioBcfVenxXw0SfGiLy0cAbeekS4PPqXJJwaqQXnEukLA1NUru
to4O4qZHEZRdJn3upLOqEvjbVn7hYptWtf1O1hS+OpgLPT62xDGSnZVuYEDCmbr/txdJIPV8hglu
ZQ0nx673ISI3oRR/zOaPC5cCrm9xsUiokJ5Le4Lp7RnTTKMhYQdOJlw4blvdenrEBRfQYbFh6xsd
c/kng/moZQNbkaXGXlOaXwO8IE65paeC+pp/yFEuj6w+r1zaupdydAg67QnVXtUSJIBvvGY5T5kX
z/0r+FVN9wk08Q0OsVwJIv8yv10QbTDZF+HRjR4vZi3z1HPbrwr0UmR0S+JSwJa5kZM2ztvyGKQu
iSFadMCp30oxttKJ3qViuIeybX0xfreJYhQCFe7NCKnJD1om9TQPUDSJXwg7huxP6I5gChUnVFhO
SwxIoxfM3KBsyt5lGn2mjEbMUSM+59ts4hrZj6nuD2Hu5mrn+/Ks6oZ9NXZ6bDeof5MmnOj2MEMR
9MOvLcXmMtQ/msWCImpS3Ql2llN6FcnH/JrYV5VWGIXzfrPpcdjZtT2elXtBbyhhcC9neCUTYNZi
7wZ76vhyRbZvVZwZg7Watd0p3vnPuTXUXvg4xKNZ/q9ZGqnMtsHqB8BoFMV1sc+OCRiBPRbmg8F8
BkgScAdP5jqZ1RrbmIluXvSmEdgwOZYn9RxxW3ewDYWjZ/d6Keg477wOp9YSC9gFzeqzZoQe4TxL
jXzQoIU1GW5aVbyo9VeBEp50fRUqcjdQpIJgEd6p7JkV6s+mPr64SZ6HF3mFvU6TYVGQ41yzaGS3
4JN241nTQypuf8mESdVrjAsuoZPC/k+9aQl2sRyZU4FPeoT5C+L6kMLD2wYS6qK9ye8qKilE4AcZ
NTs7kjSn7sAGEsYJ258fl441Cp6M/mKQvmXSebb3z5QaTjpkATUxzed/O93kTZc7gSAuDupGUApd
b2y6c80DnlE2SXkdsx1c5DMT1MURhLVC/Ns4yvTyw+xgHo0szBBNJTm9TfUBnXSYyviDOO2MkLSt
ExkNhNS7FuaefML0tREbEgAOJc5IXZM1IShcVhn4/ARvXuWRBHh03LvCr8/IxKQLOcvdFi3FBgzt
bSiRTsZ7pPg8UTSSmXhuM4YQ+R9ej0/N9tDWSsvp3uz7mKqoZiTFNdq6wn2bu+paNRjsfWww2OJn
tmHnV5gQEeyW83DRFfT0xtM+WFnm+3OFdkJGC1tyt41i12kRETCTaLVuUKmL9f1mF/prflPFHf9t
xWUBZuDjMfMzKcqvFizXwKNea8zVq7Ea4OKpkvamEk3ksrcVL5lRW8jXmeAfjC8o5mGGpSf25Pe4
2Tpaw8VXcdgfCb4+LeOma3PMCqTVzS9IBJiivIkFAKG94N/MQ8t7Fpo+wDWaid4ntx72aLnne/S/
oRKMI/hMHg/CZT69mfQZce2iCzMDhHEc8flFCpjXcMNiM+E5fbRQfRZbCz0Ox69/qsS9/8W/1v4V
x1YMwuw0wkQOGmNR7I+qypLCsP6/wVF/icRY/MqVvLE4xHQt5lbAYVNR7/1EzXsCdepslD71SGf6
X0/S7N/7U2zVd12dqOf53rLNApRYWW3VLcVCg/jJK/vn5nziXRCYXw6+cvblQXyrLDa6PqJ/Uz6K
nRqSGdmjCs6Z0G04sw15voSAC6OBIhgGdluuO7PbeT3jwTzgNP0hMN30cd8tmHecNnI4Uy2u2ZH/
tEmKn0k365C1XhStLNT5E0f6+2C8cJRtVReeiMNFroVi4JLDqVO1aF7hjOD7Bh9AcdkMuO/Bsx7J
MXUWEYbkzv1WJQcAruyy61mnj+IqADt+A7yh56eBMMTG/1gneb/KIvSpp8W9fyMy9pIB3hCjoBPJ
Doe60YRP1qYTMhjfrclC/SMCh5MH9qE9Qv4CmeHgBwoVQFIkzwMREqlwmnfKYEDMNqspwyDjtwqo
XLm93J2EvG2HloO0TM8V9VtlwOAXDpyxZ5KB6sgmjeBqLjTMAYkdwHcIinFpbuqaJv7DPC+tNCQX
mMxro1Tbs8uhER++b02X8eC8/+h+KIe/XY0tFWCesuLdbrHNqYmnkoPAONbFMhyxdGBaiGFa54yQ
BQGxPvXoQfAgUnDUJmo1jF31kz0z2/ZOvoutE/Q9KJ5Rhrv4BQqZrbX1gxu97Wu4H8vjGBMK+ViZ
8ZpN2qi5AS7V4QkBpntHQ43KLeaUTrzONFFtSt13JDOlO9XlJP/rdMFq7ij4EtYjGchCIc/bejoo
qN90HeQYMnZCYxTEfJ7/FB6Nan4O4TH1Thko2SCm81Aa8QbcmzC0JcZXXEwCbJDiK/tSX0FSNI++
aqYE3o5o59ZkNYtFPF/UtYQLhnlbzi9brpMORz6m8eBNu+/65hQATTjwb7SD+b9x0tYRjB2FyQ6u
m2i7Q1xeHzizcTLRPtWw7bOCuwl+5AbzRM+1j5e7eSwe1rHrzWxdxz6UOWkkcUjzyshLoa8XBmnT
Gw2peI1m2WGeudTQNbGWQLAa9RU9yY+yexG8WYEShGcdI3cWu/ma8p8YTMaoB/Ev1O2i+cu09bKk
wT9h7aE6IGwevC4gyjegwA8kK8rDiOeqBIiESS8B9XfKsXGiakjkqq9W2VwCBZL2STtj88q5tXf9
U5T9z/n+zVCTyCt73eUFnnKXtNE0bhMtkO3Maj+GTFJK+TorWBvBlpdnC0+o1gV4e6KeS6Y+46Ls
nD6STMgpJN2WV98ilGp8q40/qGqxZorET6N0/P3lLmWXQIs4FYLYnF7Kva/IvuJu59/iPzP1Rpdq
TsFvtGuCfqWOkmDZ3X1S71ChFn5PZ6kM6Ujb8C2fB/BhmYGq7gd+lAs40IydZzkfk5c++SbeUB2/
ubZ0Ilp9XYhNoiS7neM5bu+Wi7GJmoFYuimSmw5SnDdP1iL2wbZw+/Uw3DqfOKVpZGejcQULQkuv
ssChKQGpu6YdB/B24t03jQzqAsueMUThWSBaauBsP86GA0NHXu6mUzUEHIHBMdDNpXpfsymeiS8e
w0K6eqxJJbNSmQvtmh2VABcXDsCZzOnx+EWyajIXVuKv4aCDzyJ8HQ/af1i+MQ+K9T4xzRlLBSos
MwxY2MKnozCZK/Ht4x/IzGiqrx4KLXKDmMwHQmCMAf6iordY7kKLFjGS9CvDm5enKoIPzZLvVeWg
BYEIxxBNDXbAOYkTtT85YcgVQtgSTvI70yL9yMkVdQwIfclktjropSRfatb7Iebkv6eHH/rBQFJF
eeDqGR+SpuixX/+MSmo3qMaP5qBIgMpWfhUNtk7Ta7L9bAyQb5G9ckOK/AQm0ovB4Q1tUnQCPZqE
Fmpu9mLvel2fZBNpTnrS+Pi2apG1Er0whWPJ7DFWh3LK/E6hZlGDxALPBzwgnOBZ+tcWUiYqzaLn
V+9eCvGKai9ooQl3EYpzyFqCjw+nKn9L9YA5fQPQF3+dlTP6eTpgjexjYrQfqxLSY+AwSf/8UkBW
hDTAddCcQ5AuDs9Mx7inE7CnE91KIlpldaJbpoWTxigBeS905DjV9p/gJlSUs4wRcQtEZugWMqes
mNUswntCR7hKHaQ53Iul9UV7eZ1+Y3R43Nu5h/JfMAxvgG3/AuMsuxreToujM3pnlPU3i8v+Xagd
kAx7WlwbQEHN0f+cGwuxMou+WGgKV49I3T831xsbZdplW/TIExTzwIO+FcCL7+FFJeg9K6FrxvAx
QwTCZa1CtI+5YW2RXHceJILxxLf3A4VhJT+F51TZP6HRYHS9U1JzsuK3vBuWd4KOH/R5ypBtw+Yu
/bmnSFG88+xmDg/F/epzK2/HGJthOWQbDDxF+6ZOXD2EjXYPdb3/djjLZ1QDbzBF+hFQ7pSWFB2i
AJJGPl14HBRdeZ7jRyGiicCWjVx9Q3yV6h6vxweNjfPjLrUXAa4DWale8VW7GO7RRADtEVYH36Hk
nNJr6Vr387VUYcowLQFd+Ev0x249o9teKhy5/1adm+RmbeTcauhe+F8aNuqEjVv3tPNab2yCkU1t
9vbNtwn4HDIQ2Vq0SQXJucrppmCgChYWTT9VcXQpKL6+dhVcpqKyqC0UmUqWMWrbgwC/2pT1Jgfb
MmZG1IzyZ/ykCNSMUjLMdSEb9HPXjJSd8B+s14iG2NuE+pivys3oldT3z27Bs9TaUFsalgen3H/V
lzlj18qvoirdxPbTipFAIUvVHJ2EunSYwGhMHTRDK7WbkqT7K+9/EL6mb3c/fr4bA4RuIGbWC3gY
mbSnZjRFIuL1apy2bRjZc3XcUaNVct0T4NA3/t+F8uvubP0lUnh9IdHFC4gYOgmF/otFbGjE+7T4
jrPB6dN+Ndyqlnfnb6hoKVHleLL5jDn9f6kuvzt94GxtZKaJavUHqDIjvrCthnaT7D+QCf3K7P68
g0naAsM75Cpri9mEEYsFXHBGK2MQA2PyaaJnRFSx4YaifM5m1y+rpGeb3gYga5MnEzEcKFlsB0WJ
qIw7qZYoxkc6gm7B+SiQy3p0KZIsAwC19D8geBPtdUxPHCBxmVy8WWPit6GAujzYta/9R4TrGKDQ
vfme7m1Kunexbp8mWTvjhFcB/CDgwudhqStvYjg/PcGJBDWhhcTcYue0yu8takLShXVkAHBc8CsK
6lOgj4fVGlb4gRJeN0leUyEg2iJywSCLvNqXbLK8O99m1iX28LkJ23d1UGpOiayl9e3Lpzb3QgZ+
z79LTiA6M8AWp89Bg9l0q+9ePDkW0hmImmAlwFhYNojU0apqfDRiz/RFJLVOqQLohi/u41KQF8je
wPGx+rPl49sadLP73a9xTzP+jwInYzHpkBBZTQBoG1SVUVbP0Ufy7YOsBqY/zUgJxANZNEs+lyQi
4YkcIj6jRjtfxtAu8eytS8+5QmiDR/CS2bKHSt7wR6Jwuj9JNISjjaZPawKxsKhSMcmT8MPTIDmv
QuWMhkaNj/ZrKGBYgMq03ReAvu0FcxQhu+Fs7TRqwVzB55xu+myTWB/8y7lW/ZpRA5bYl3ridNNZ
ZnTleVS/ngnHMQc5Rof+sW9HAU+uMbg65mULTravJ0/Iu5hhZZS2vEwAefgPRMMYSG16KrNPssK9
eOtr2pg+MzjWLSoU+zLoaK773ybpnvfU/E3gZZeJNKE1RoiuCWLrc5Ypo2MR6FnDN5h4/mCKbPaL
vzEldtA2uxWxEgjegAh58y9t04fVHdBACIPkrZyw5U/C0LGyRD/73vdZvJSNqHojnwbWJC6g3Sx3
/HIfb2ECc3txTtEhjgTITWG/aEYm+msU4gt8nPCmskX+s/y6VUTwmyxvy8RcfzAJrNDF9s97/oF6
5x4LQiFNnWAIPlMYpXKfNGB1UWRsqSQB4YRJY2WIClCLSs1o8XdLk1IhrNdJk4iv0dwrI8yCbQNF
8vxzBwkqTRax7KPwbWhCu7OvwhFEz/lsWtJRijNxeiHxUSlI83C8E5vl8XEaQ1NbO0hjJ8rlGBlZ
K+L+1Ovq7oGM++Yy4wobqSUwEIh1ziyjJUH6zD/m5VjjUUT1Ce2Ue/92/F8evmXusDXZA5QXxEZ9
OcndoHJ0BLXTe1Z9ej8HDdnl/fyDcxKhkWAAGdghXMxIB6AgLRAiZ/n/xQISTYCaWYAlOnYD8WPb
jRS2Ypxx7BMdnsrk5XRNG+S+2vwlIsLQ7V4j/aMVAEkJHG5Xi1EU0hS2Bn/Jff0SReSXdvRh14Qk
vje4PK/J4m0uOePgc5sbXhJFl5nkTMrX2UtFP+RrdFWvk02BtMarzRS1wMwYqb7oX7FOzqRC0DMD
z6u9Btw/Dmrqm3ZBOqdJu2n/TN51rYiW0KPtijMpfyUgbzr4Bxra3o3MFYd3guzURTq7btfmAyBk
sWYWNvJBV5JVmya+isiwgp30Quep3f2AAP439OlSpwEd5dyJjUY/XRgynD3nvKF+Lq+ttNZqQA3c
ancXuC/X5C7fQQPHOp83hy0iJ/bdW2ijCkKaQLa68trny72Kx8IPdd9NrcIDPBRCqyZC2naq/mvj
QsmyUVi6unHzCPDd6FH8L7AHmR8hnB+20ZohQj5+8ZCLopdvsk7D3M2ukvAxO4prBe1G0/+Q/92k
xIj/mztwlb68lX0t2nOV2XqV3Ro41pc/OEmwNXvu9rcc5gqw6uid/ObVE7uT+OpB6QeJo28VMTX4
dL+ERy4txWIfEn8qs6CJEoIrUYN2oVSIjISRpdfL3E+4kov6kaJZDS5Y2ERi2qlWgQVRsUs/rwCt
MIYNJr4Og4du6RdGVjDfFWdA2k1aEDgXytvp060Oy6fypSZftoneXqIkEsCxzgWTTfupqhC96mLw
g0Q2MFtISiwMRFgb6UeEcUprtkgzb1OcBrySkcBIOALwn6dwFLIyqUOz+X1OQDif4Vwlu88LEEGF
H+0gbkxlSp/lGB/zzCOdfuKbX9oPSBK8+iwysqglAw8kG8gKY5d6yT5TRI+Tm7V8Has2qmefU+Uj
LL/bmpDmaeI4DRhPKXnF7Hytao6Xi+OJeeiGD7ZG/eccGjMjs2bG3b0XSgsKpmm2YN89D9Oih1Yy
BQGgz5RJb+vSpHZPaZP/sqE32AQ4yOKqfywttClc5dq+NEcRQS3AEmFpsz2oQibnD8NB7KbSat5O
lgE+lvpG+dH1XSkfWSYyr3HwDcepwz4+NA8TjK+zWGmempjUDNmw3suxSadqU+nvcpneEAF+HZu/
zUllxnbRapTgPh785WTZFFd1N0Ee/RlPr+uGkZ6lLLoaLTIPL/RYrykO7nrzmgd+McKEQIdhR3Jd
Hgq6IHw1QymWq2w80DZ2h1mLilyHzPdFCWkzuAQ5Pfo+Q3KdW2IfkoHFdcogtmNwwX+xEv6806oJ
jkss07OTGx/Euk4sZR4mP9NotFSLombMcoTm3QEhVacBj/kib3m9pm0CIP5UmE+pDyAyMIPOUDWu
nURoFO9YkUJp7D1el7GwiHpprWRWZTLyURXMskGLYHl0t1mmuCv8I+a8huz6EkuFz7qNvEoFx1J5
arQgNOP9kGA2Zd/S5wKRx49RfUylAelym1fHamH0ZPtkD3vm3yk8bHfuYwhkYJSeikuLgzDCGLOo
l0uumzOsCnVKc7vALKbHPCDPbBxeTD6q4OV4bEubuyF5Iz0PBzyV0Vtu8hQrVu41y1UO+5eOsZob
za45zlNkbyuK9Hnv+7emjhWucpG66XFfUzQbo+HY5YrAqs5fR41TUiz4TCLCM96i52/Ccm5BK8da
/yC9tZzZj0HnbUVRjmeM+17seNqW6da0ATw9bIjbc1HRbXzJVBweGaNm0ffBEwoPzcEVTBP0JrqK
doTsg8kAItS63PDWNuK8g8DhOT4epgqeNQQe58l1n98OGg+Ew/S6/ot8s1J57/BgeUnG8N6fXhdS
DTnTI4Cxks58jVseTb+IB8fkF0DoZQNAcRWKo+NpOVbJSgxbT8eeD75qlbdpaOUY00lt+iyHi4sg
2D7XtizZcvfytNBj+DIbTl915jkxeifP0ZH73woFqzxO6gGAiy1ShFQLPmy5c1zvhcjpuBtWznsL
e8GiA2x7kBXxJigzZHb/niSsJYAujW3WI8L3j3SvCuA1u9XCoArsbc025YjI+thSG0WMzMigZhZZ
QND5yn+yguNFGh7EI8sJ+8SOmQ7qUigOCA/6pjtELN/XTgA+BRJhB6+zzbKy9hEuc2XY4shH8gtN
E4+34/z8mtusccVVQRDQXq7n6LmbvCfIeecE4rTPIjiH7TFFYktJqXpIIC2HyxOxptYNagt/9FB8
R1kSbD9Jyi4Go+Y59NJiQP7Euwqg4nPBxi9ejNT8P+WYvCIaS4m+qYcXnov6diaCq2/6LdOzp4OL
GH1w9T5A/9AuUXFoESOdq/AycBdQ5IfMdkBhKsCWasM+56DE+Nsj1QztylnFTWaKyG8NB87ZfpQc
b5zjBMZZTlZHY/GS70ju6hBCfIH7dKWtgZ+c9PWIbspEvhnjQvUMoAUWFVf1iGy4BifuWb5pggi1
44RWmtBYsdOT1YKTKWKqRyeJtF2FzIhtBMtpgg/AAvTd6mCldXxfNcuFVqCiuzr3hAsgQVzSs2XB
mgKXHrtiGuC+zqyLbUkFPRzTIpWvfJwXwlihzgOupjitU696/Y8EO4sHxwbAHgEkTbreRTVaA4Gb
H3IDe0N+wHP88fvzgrlsMxSVtKarOenmhK0yFDTd04lHTCfGL4HXccCrQIB0fMS0AYmNeCHKxU+1
+2nM/LQ6hgn6D7vebAtvToKeg0lylHrOCfLaRSN3Dy/zVqluK9HYT5A6M8BHyQj+I/+19LhwOZ3n
K6718+0dTlZPHkuIGPTXZZK8cevkULi5ktNqUMcM2iOEDYJ5WnjbIbb3zmoqMooISHg63QrphEto
sZsYJFbBvG6wkFiiJJIf0VxLesHzrvWSJv2t0nngLHt9Z30f9P8uOtg4DvvTVdjOH1rLNmm9Vsr1
XcMFo80rWH0lwbQZdpYM/tdT/A8tqPc3OjbI6lA812ll3wMA53FUMd/GhI+3V/WljLHc+OUzP78R
UBVwLNoG2q03VZLW2NT6xz/R4O2AmuoTcepsqKBovi7Ey61dviob21equvX6yI/WghOfKa3hLex0
lp7NtcwqIImSTQlXRHHaV9Xh0f0cCpf/ZE6nNRNJYVXkO+jjND/R801Y07I1DPHs17r60Q6Dyqpk
rXLA0RBCsl41/DPB4kXuPQnppetaxgV9gF0RactagMd4JAL7fwmsozhLz4G1l3vUSvKwCjiIHHfk
oQN6txsHSv8oD1oZCnJkuDnLgMqGnCZJa/nEXgEiIxQKc8sTWk50uOgGTYqhYcP7PfFbTVZR4txQ
O0NBAL6gSFlQQ8ditS4bRgTlgoqTjJzHVL843NIkRhdsFvBFHA6ksN21MVL27L/L3s7d5cLw4QDC
Hhm4Es6mnGRy8/qcTluAojcbzFVWed3ehlGc9E9heWyOVWgmeefl+KZ5aNBuC+9ughoG38czeIX3
uIGY7FNicJVscObtsF3Iuaro4QnHRkiMlkpTkzT2aJiwDeYgQ/w5H8K6yOMEBje0AL++ucBkzjJt
cI00nPvFIKh+8DOM4eu20xGL/nrhRyq9Pz+s/XfOwLVVggzhmWiImnF6cT/OZsv2aPZyelt86RLT
ywN7u+lExyDZvzlYFsE1QCb1FKloplESkGnznSkYkKr2UEjTrfTf2v+KM0XfsqamqpNLAA54yFKI
TPvpiVC/hbPCGShFRAR/Se1orpCnXdURSGkxMG8XDpaQxPHqQy60bdAjXNtthOEnwsV9/+dhbiPa
+VW956C4JSpsGyQ5P73hk5SzKPyA6w/viFnFUhofmfxKnLWi+yUof0z86zIU3+saWS/MbDigQZYa
/Ak/IImCVc6AayWIudfAZxlb/cOfT8HaBkn0EnAzB9I9yIGfahM9W5XVFxRoTPl4WlLdNlQDRId9
EWzKhQ6NTCX3Z3ks1NkhQY913nx+vUC7Rp0+ec7z5Oz4aMk0vPlhDhJHmBBO1qz69us2mfhWxPY6
Mg016iH0tNaJCtpzrjM2M8m1LdaKkRerzgvFOidM9P8tfe9FJjE9YwrmoLQJEL+zcFKGAtqULma2
nRNIuhP6+SqhpkK0x4l281oNocqRBgXmk35eG17iIMj8rBsCZC1ExZHCrKEAI/WweSSzZLQMnYzs
B+0Y8ChA7k/FPWyfrfW9QXxyjWIDa2a0MM0/kdrDPdGnW43YwwnvgKZe9XCwIJqwMO4jGvoquNXI
EIyk8rfuiIGCWNCrWM+JiBXu1DBHuVB5N2HxfRcX6FEZve2R/2XQjl+Y9Ci9qfnkHAasrkmxT8ZV
KsV0q+jTZGMeG6MLoPme19XluixqDRDE8L54L05D8/A1Gak9cLYmmxRczybZem+rSXBV8TmVLEv1
ivFK5/obU7hnXFvvW+C5NJ2rZhnDCkSFUC12d5SWSj+gC0DSyOXtgSpjYOfvrgqnSkjYNjZSeteg
A1hvBxjMg4LSMWDiUtvyXPHZfdkSS6KFpmVvZmUDuyrd/ttDY064eYcdYVQ1DpHESdiXEOP9RFkA
k3AVlhVd6FUIcI/LXrc8k2J4xqiTbDvlgv27qtCPzp0wz2gO0gNEXM8DddxMo5Wyak7gtDEioEhM
BtKZBR6lb0tnMaNoe6EV7E0V56FiSwJDSMXJv2CoHagOsSJuz/+YVJgVeAj8KATPksiZlwXln2XE
hnCNdnhMxtXciI+UlZnYKO1MrGdd/d4ZVN9L5RoKpzXAIxSDw0S+qDEP1mwHUBUiDHHdh608HEU8
sDuUHc5LLxmvtMY3rYnS8S0nedzZGqvdm9CMDULsG9Qy3uZk7zemtV44gXHMCWuhBE0L/gku6dpj
Nt/oR/VdYWUiXRpLtIMJRDlz2MxEFkdK0GlFpxa5nj25t7WvDGO71mTHkGbVR41JB87xKlEepKvN
c1PnZ57sWX0lPOQuDoFFoqW5N+scV9KY7vr9uveE0grzFV8qYbajwA5O2SsNUdkzNgqXbwaSw2Uz
HdbNV5ZfKk2YCitmG6mGXlyOlPj1GKz7UD0k3KR3lKbYbzQIdC46q2PF8f8oJ2NfHiNzKXh49LV9
r3wTSbbY7zKlchQcY1ZfmIESjmJfxaHGP2jhwt18K0dgq9SIbr1tHcTFI9mzxtv/rmnipbghVfLu
mSJQhdgndEunhya+cwpsvYiOd5pw7Er2ACF6GjHrIknrjwmf3OD6LesG608rRwIoZg3xtbSSRYnZ
YDcK0it3x3KMIWwVR6bu9Kwf3ROhpK6hJKPBH8TwbB21nKk47BIzzFnvDtR/aEmWcMwUDL0pPiw2
r2nEVKJxGcFLpYqk/MFMYF9S4GWBQbY5gcEWRW+/NY3rkVYU9u3F6nuCkVGnwfsEAit9hJgHII9H
/GmM4/cEMjyYh+QmpNuXpP7qYKhhUZemvcH7IfSEn17YEiFP0+NLrz5WuoA6HO92wBSQk2rPD5/W
A5Ht1Noc6SduOZrM+bavz7y1px/kfSsrmFCWCHx5/+pQv5s+Glt6w/OpEQkB+UcG4cncetixKPDd
95lznKwL6qYjS7fwLXFiaARplnFOCuLBg71mLHRJZsfget73jt1YU7n788gdiS1rB4JAePm02o/O
KukHE6RG5BihBuchkbIh0NstSoPYwSUjMHzbVBbNtkDmAeH4JZVoVEv3aJUK1XDD5CHSoFK896rV
CjjIpzjXth92Ry4eKZoqNMis0Tljui2NbwVpqIEJIVnjuX49IIh/KGEW2ZQaq8rAHdu/Ha2Na7ZV
X68p6K8eDTL+yrvTGja/mBewpFwXVUeEtKCRhIRK6OpADmsddHL3i3lejzRg11rurfIQlpesdsA+
aY2JN6axL/qvD6hpKMXzGBxguMJQTxCI8WK3dogQi76cEANtfwlhaiGeTdHYEHYHkuiSNrsmDJi9
KYOSdeh6sQlYxAc6XCTAAqnKNYKdei8ksxCm+M2PUgOozfIpybkXqvUd3TIUUShpR5fvy3P8DShN
VykRMvRKm8JMnuuPMd8CD8k4TwDHMQ6PrHFl+0yHRl5IYqNUpQULa2gbrBUYIaZLqPuuLHX+ysnq
7iG03fLZ8R16OGfU9kk/FVAV1C7U3/aiWblBJe6adP3jcygOOrQoPHVdGU0ichouvfHNbUM6emnh
ShIqXqWwcY0eNB/5n/HfkG9ThgNsm2MF53EPKN3EFNhRrfDL4sPBGbHrEoKve4OpWcC7lpClcNWe
mZhpi1jBisxeWtrCfsrgcRLQxHvikyVoQ+TkxlbwaXneELFUbXfQLBCdd6Le3ntU5lHf2zCwKCOH
Lt3OImKuY8KDUifUJpoiR3Ps/ZJ7Q9RQCkFpSlS5hVuD1HCKpVClBdDx5uPYeLxR00x8U9LwccRD
mwjzGJ1s/MXLotWdPB3sgLM3NHgG8wAKmir6iValJzdn2VVFBLlmsZZb3nDbHLXunLsRh6rEM+mn
2+V9ViQx4+4oh6MwrvAKgrXLaYnVFqK86UpzwzUOnTncpDn0thjKfWJiDNNTlXm2BM3s8wyXEeeM
ltEV3wVsuYw7YsLzOU9F7LIkQFl0GMHypmYpSQUZi3ig1siy7QdAbGBNdPUan1Rdd0/qgVAAEwxI
8UyHWbOAsR9JjX1U+ruMXyWH2Kxb8nkMu6lxPLz80dwNACboY+rFBXcxxvOTf3Q61669nubdqC8H
UhRRR88QWKFTB6BpU7NjjzPlbl9QOhZ0JdBaNRtmyVpOPqoFo/HtmdAMHSlu/Nx8XcyADjERSKrw
AkxSSMf96Ryp6B7rZVNzDLkErGETQ7HNCDnlHweNO2YNyiaZ4JKtuJrY4XWKQCYhOZJFMhR7UxnQ
fgKXIjROrtz+fhBIVCa/2WH1Vv16kq0hl444lTYhLbjpg4KymloeRo+V/P9cnlMbKIVFezm2hrMB
E94FiKpO7408aHjLfMCQwazVdct2x9Vs6qMLDHfKTPnPPhx8i8YauTQjUMU2zL5KSU+RLPuvA+a9
ssslSMZAD2MSLUha2h/6d7PXguS5ocgIl5oVUTKybV+checSl6sj5ADA2ozDdo8GbZVhkHsxGzuf
EFsxu7hntlSgGEdCwaDHNtD4zOEAC1L61k8IW6l6Ux4JkY6CRGKS9kwhIK5WT//WCL0YQl8/CClQ
cNIapf3PQ+q5gP/4U79pg6pH/Ymq+MBAt/ThfLjOgPp6eTfHyd00SoOoX2GiqkoGVufIzIQA8xQo
/iKDe0gGCHNs7a8T/NZscMpFAzvz7Bnblg+QRVEHRkIFAOmcmX2b9n08+b7YSc88T+mAS2ALc0xx
M+XrmId62dRPA7kzeELu7jh8bc7hUVfhnD5e0dmDIwvhztcO1RBxHZukdkRQzz5BDA4XeFOjaaGZ
QluKDAAc6xr4/7gm90r9s8Rgfp1au0bHCTuvZ7eIuPLICSL8kJbA0x1eh4R72uh3h0pRQUrNAU37
DL8mnJVKEFLB7cDfzGjqKQklRwHvWjYFCK2e6E1rdyOLHoqqcWCX6rba4MuFF2hFVyz+EQKgTLen
WCupH0AyqibCMI+pjIj0gqiEiqklQoNBJN7/MvJ9aIJfw6kHdJ5D8epiGCwM/7ce7GYJ9F5hSsGB
eL3xM6PT1nUWLtEZNP4hG7Uy7/iKntQjZZr7vmhyjyQHpAddev4rC+V+jWsKqkjcp/EKF0qKyQol
CwSddwEWLjg5/3BzE3cRy8LnJkw8g+5bFhnRlVTc2IA96p1FiFvnoEB70puBsLzufaizskZ5bpgK
x81vJpeqNyHpgPzsW1DfrHjd287ntsiKdY+YCpnbLTvyaCMJeI9XVvsZ+/jrZfyG+uGad4ke5rNv
pciS4aBvHDu7WRxSyVDugR4V8iYlhR+vRso8UpB+Cbr3ptmKtn2LA5Yhw1bX9vxrYjvww1OuszKb
t0m3DTYrOnRYEQWZZ9XjYfqrtW4KXGmef4yB9SKXy5bBAIYy5OWT20/HVzm89dRkYU/27+hbFQZW
xN8dzcNp2IXmxG/+4qQ+FLguI4cIhtI2goJNVqdwuAjx+1n9b48KVJ/R9cy3+gGXYNLJXgM3OFaX
LlnezJrmSShq1nUrRgthUUewzXeEdvcGpl5ud/XVSEehUlrkjJX1hJKVc8NVa8EoBsj62ubyIhPr
0ObqNpv2Tp2+QfeekgBsZCBdT4mzEOTV2Xmb7fWIsjxN3HmwMcXQqVst8OkMH1OAiMs6EtUk+lk3
rvY5f58tvrrmC5CXwNCkOlFovgb6qzaa10YtFpr4I2vGeX/gd/Uh7D3hb0fg/IblGhNr/Plg2eoU
EYnVztHH125vZ3S/3MoXYqcoidizwUMrux5pQ66IpOVwoUJof8GNZSvTC24LdBvNntEt7mYhAHod
1mfqnNDUOP9shElC7eFyRCYX/Q1so1O5nZfYK/QFpv6+pW1fczYkZU0NXs1WXuAiaxRdY9r6IUDd
7B/H6fcH1F3XycslVPDyZ3kDw/F/zzZ+DKsSEVTEC2zPtCUvlvRqfkDyVvsriYfMNw8n5+RsT441
QWBqPi8x6jIqR2MjtiTzakgTv7WbzOVSuKlWgQvgBrTK1uykX0wGHwDWnOLIpk43GL6gNFmz8KLd
iE7u3xwJW7w+DvUy2CmIA7T24zGVQsXMtzkQV1iMJWfMKUNC1pBv3a6bt2aV2Np6UiUkdGAXyGDj
gRCJW7XqL2b1fn7pe1PVs0QgKXAhVfp3hCkbY1FF8omCK61JY4F9axZmmcTTpSEiEbeGi1w7qu98
k1mjlpfSYaZkcok55NKA/eJg3cEqnVnwFt3hOhuVpQ11JJpHw0gmbXxxvqDJsEQZN5RfU1WCvlsE
zTpCtY8qgeIzvKpeszfHn2Ok3a0hfSpwzBK1wzIjWXlh9Rn9u9W74j7IHpneIZVuv86wBAY+9iCX
To8zGv2reBYPeJgLDCVZUOBwwKjSn/l5a/pk3oU3bmcMdSF3Qz6cQVzcEgX/6lPZKBNJxRpWRXgF
F3kr+4ehxHOOxWcvzpviGCndjlOWTMndB2xUdWtdfXpI7YbDWAi3OyKRN6avc2mZP/pki5RxoYRZ
rNxpHVUZFXD4+xJyj3bhhlZ3oC4y9eB2uiRvk89PUgWRtU69TdHTr9j61U8CDiUEnbgQIleXF8gQ
ddUbs9tfajV6jILeKikYW4H5VvilXHGZJLUp9o8jN5tuoxUNSLKx5gang7DM85yMt3g/W5uJTsNc
k4b1meBcRdziU3QbX4ox1txkXXEfReymeKwAklrCdxo4/2V9JBE/PNopgyHk6ngMO9/6EIQdtDWt
sMkJoKvvDyD9stwUXN/NTUT3IdJZZCX8UwP7aySQcYts1C8R/872fAK6S7E9u78M/9wbhT0QMLOm
QYrM6zY8v+b49BZgR6ZeO1IkUd6UXlKR4V+itrJJr0ryoV1By/CB6BGmH0MPGseAZlNFGzjKWDw5
PFMIUwIVcPzm2pIzfzOxEVlLXww5PmZWQKEtX7OztoCK5FK6PQThMIYjVqfhWAIZCyFuqb8JrliO
fW8hRiQ1uJ5ri6xINMCZC6acBIWLg5nh55TTlKdcmLsH/Eah4JL6hyTC7EuD7uMgtB6m98oXEsOk
blSUlGi7JqxPs3mcDR3oN5FmPGv8DbnMn1NJtE4lH2TeRUl0JSNTwrcjcW9tH8LxzByJ/RJ9AqCG
41srjq1awvy/nEJLtd52mfN0L+iherEXWJIyqbE4VepvY3mMEuwgNNAyGhOTr2MwvTTfv7YWvNux
3RT8PXl5DSbFGhti8l1HueITAYAIL3GwQaElOMn3gFdyihJbqrlD5MGp7/PS9TzENxAjytb7MvlJ
9IOMp3G10ePQDm/eKQTzHXgiY1gisxTzdIftzea1BgyDsCxyj1CIwYm4klbfHl6bXPKhO6z4D8hZ
/U5zrC3amy3Svx/YXH/YZsZ8PbFWx1HSwxyaQ7Ya9eAw/zKMWC95MCh+2jSqN+AwZSDBK3AW8Okm
KMEWjuTUyQ0wGmo9VuOiSYSPhW1Z3BGe1zB7vgfqdsEljSgEccWcJh5Q6DqXPYyjwe8xYAhV85qW
UzwFHuONViXMseMkXZaLqPaE3eUfDdB20q/Gavz5Bp4/zVNSgL6w8raofJ0pLNpD7rsCu81fJGDI
VcmmXvJcW1sTPTsJ6qj+zZnHVW3qFcRRrQ4J4qGY5SLKC2gY+VuZiyTeHZbO6bqIPTb/9SV/n0zI
UdadO8//QDFt0jRFIZP+qBFvBf2myTj25GOSyzwL44MhRC3+tVMPBNvS3eqWV9UxXFqUzAuIzsKf
YmE6P+TWGliq/6NyyLh5MbKxF/lwJC+9KvcamNdlg20t445hLZNof59zpBvW3Ll066h1WICmUQby
0dfxMdLqMlzSigQEQDFCX8H5qixzb3e+pNywnAWPX6yM8LnEOdZuneBH0zmAnB4MdbpbnLEyaoI9
yvLA0Uqfb2q8NQqLz38Se9fgfuYM5FqbSh5xS0GJTBs2JdP+BSthRfTCwXtIq4rmXx3usVPRm3NR
sVUUzbzkT+Nl+5dmXh1analo1FAQp6Y777p7qyvQpIQK+8iGK8vBMHRYAVFh08LRRkZQFDsgnjN1
S6rr0CaFanVnzKk2P2vNv2/TxY2BwwW153RvsnG9pz6qYs6BdJXvIkqY6IBpqnbyW/nW2nupmiDq
rmJW/1K+AcTjPPY51lGhWcmYAEo1FzQDq2yHtwqVSrwIVDC4lvV/0/2LbwVr+iUNyhYrlNiZUBPt
PcGY+YPCtJQDZbUhY4xv2Otg9UiTjo9PnaSKVE3KhbkV4Rz5leMjbuTDPFo/jdRU7oLyKEdjGs+l
oKnpAuaUCHXZj0sVl0z7yL2X+5HsrRYoBGGJ3W/qI+/xdE2gLdLtCiXh/2o5C2Xf8ZaaMzvL1+t1
XIryel/gJZLvXhvV3dukbRrAg/Xrq5JFpoXDu4zr1GVUt3W/1BUSkwEuXwvsNS7KPAX2ltlaV/MC
FscIay3LHW35HbVyJw264ZE8YzN6bRzGBRIdo3iUpuzC/7M8tL1FuKxyPXfZCpBi9h7ucoDHM6WE
3zILCOcVHyIg7yb2aTMT504sZkDqfVByfEFR3vzv2f4w9QV+DANxvWPP3TVh3V+uVs+PMD53IFq6
FIrxOV/RZaZlVvTAQHg55lx2cqvgIWPUf9TazDfgsrXAClZ9RkToqQdkmt/zA75BFNR3IwNw2eHH
QhE3PqPPZ1gYRn6vDIra3zO6dwJwSZWXebfGQnQuG3+bPIB9kS4yeTqbjZXLWtM/zkZ30koZky9S
qNbqWwdeD8/abSag2Ew50ZugYS/zT1jCg2P8f9n7oQERP55RnnPox/aTJhv82JFZO2xAVijNWZ11
6iLHqvXx5xMML2YfuuTpz10NR0GxH/WkMbMCR3d8qD/DEDyIGP9E0dOIqLmvl7+m2F1TUYzfPdo7
RUVdXM4DF/MvlSw+JdAqfB/XPEdUzXlplC3d26kca49OinZz68Jr7esa72Kw7Icw7+a264PXOt2k
RLObjMVPsljtvYV79ECJOgouHHqk1ZKeAdjw7a6Ky4+xc96tCxkktQK34yAqokv683WUln3P26rf
yjENLWQUwZ9xPcSWeqNnTLI8MlqkcjaIWXdMPoaTRI0k/YIUeQlHyR7c2r5W2Mg3DYkyzlAB10b9
71zscynkDpk5mAsySuksbuymeNINWRUvbxwKbuLjOMC3errj3NPH5MKgCJZzqwfl/D6ZbOB04+Ej
+OugZRmY1NE0nNYqNmcJOgK3UxrKrjDqAfAcVYZa0RYNulZvTPBpuvvBqfYBRLAuXw14EKjJI6+D
umGP7FKYoZOPdrBjOs92b/D19C7SZBaZ3XI6+cbEVLiLKhUMMeIysN0+oB5zDPPJyNbQAsWnO2tw
7RBupODmzA7qF642Iulxh/3Ghe2ZRcV+Y4Ed0M9hWS7Pj+hZUQIOzhOqV8j3FThFSVKhW42vXqZD
lR4kwzkrUTUN8M41h1A+hn4cfHOKuJ8AErbbWdmoqR0W2SgJXSnqw65reSxn1twdB5gtrc6ZzOXn
HeFVrVD4VMK4bmH4eUpgb1/6gfSzQz4efBVFdGx9inXB2hCu881k4hmVvJ+cXOaPwVyH6PqyIr45
oxdEUHEQFfFedDCpPifRX1x/HsS9Riu5WCfFSQD7/3+9efF1hdrwvukV0KY+GluzDxmhKc2LoFiS
J3Nm8n11tLxJ5dCzNk6ig0VFnylH4k4OlAyLYvFZAcBn9Ac+VwAxpLTZayKexbyCV0/XRBH/8Xo4
8hH0Qh/qtI/bfZxNbRwCEn++ow9R4DJ5OdUDz6LKfCViIR+mnwXKqitYlDiHE7DKGiFaumP/Nn88
7/1j2VANqrTtJnsY9woGtIB6xRA3KE+mPvsSnygkCtepw9T9e45xEUJKQ9QyBKiweR/dB7j72aE5
jFrf6jktbHU5X6NxEB12I976tqGhpuUxwjcLSfuWcJHXaxKLtTpm8czbNiNfTufxtBJTOm09w1hM
dUBRAqCA/ROaxNeWLc9j3rv0NFlLyKjtUQiLRG8i/ZhA2wUNJi2NRsEW5xtWfu+JZCnohd8Gl1DI
ubdRLbgaTnBOdVWvHP0px7pqIRiHMKZJXCsWMI96W2fN0FIaBLd7jP5BfAVxk7/tva28v6IrVgby
3SPT5XwgOwX3T8XCNIQeMKOjxrN1r2xDgA08R1jMV7wih3hX25t7fUXokL8Fk87VjBEh9FLhRqk9
L7Xuwzn6Qtnau3QdNZbm5IkraYgM1ZSRLj1xsJEh8n0888t6vO9NIx7dvC3qUXa9FZFN23a4Yafs
/s+ju77an/lWd/CiP+0A4s7N0gS4qQ10V5nZa1v57vFUJEJoju+IgS3HPQwgbpOwpfpLVqqP7eJc
4zkBS0XSdqpOb6C2Z+eBrzupL71nUOqlu33ARyi90my/x8gn3N7N/M5qM0rNfFBsaBZLKpqnXJbI
Emq/tOJm3cvRjw+gesBm0IW5C2oDIK5sTC8fn4yTg3ZBTGj1/+etIHIhQOL50DgjQJ/sT/0cB83M
OBrfseC9wq/84TGRQdlnu6PCswKzHyORjA2CO/PYbLo6/+7g4m1XUfC9Y+vCZs2Ye0rUxg5E1qnw
S21SAhkL66T6pS8/F8pN8tThIIuYZRML/yhyA54oBv4oUi6z7o9jDVd87RnBvhtgRnXplIKWkmu3
JjL9LWxSrpUCJ2zdkO19XUaZL3wn2FvC3EzeLqSPXgFbXqe0qMIe09ZgYB40SjsgqX8E3UwWLq7I
DTS3A4KDIN2KAs1MQX3r9+nwrqj2xxoQ8tWbk2m1h6d+2saaU62E1R+rbTqoHhbrAZi5wtIHKTev
SdBLhM8UkG0/rEJ+FwPXjJCRuRxSs+nfjDfqhLCQFxi2CjG3RVzEY3ZEW6bsk8x7jRBQePUDeLp2
88K4+0IEDS47tYbdXPtkzwDBvFxOLqGjNyp4Z7VZoJw3agGgIE8YaZoxTPna6HPOyRyXkAjHLNaG
MEefHYl6DzozFBM0WWZt4W9YNXjLyoxQoQIbLYLKDOoD4Dv7Uh2FP1Gzf/vu7NnG8znt0l+bSii1
OxIlAbIxr5NtoZiAAGOcIJyrJlEwX9/dIlKDkYIuCvYW8YRpHvWVLV/Jxyo+k6jGM95jsFN0REgT
BSYBpdS1hgxm2hdToc52nUEg802mBjYcbSDsn0LtqLu58lX20aoMotM761HzuoZMt2ZNx2liydzV
qIDeE7QvxDBCGO2EFBANMMXdFEwD0jKPqgrzBf7PgSPF/RyYGG304meCPFjZJCX6PgznUVUnFH3d
vF82QzbHpvYj8aVBJ1QWTb5H5+W//6oEy/vgJnfvX6yBzgK8eUYbZlxJN24DtIFfptOJDmjVJcDI
6q+/7nYdYlIIuB3r2H5V8gybsYZek9rAwILjPMkig+sXoyCXsFM5quNSBSFBEAs+Y5jwWdU+5GMe
v7ZH3rv9jdxtuML7IBdk2+NPnPVUfLuRYV0EUgK5g07pTUrfBXHKnIfpf4yEaZZZGEu0lUQCS22e
nGLaQg0MsIjGfIJMYr1/i+JlWNiGPEx5wXPMxHA6/GyGJEwMyaX13VNSYa4iecVEY0RGOfIjClJy
N34tZPKoudaAsCAU1D9zf7xebDjUTA8FXpKOfUWPLYelHo9+ukSG1mPHv8nlqjf0Q5UmfGZ+3dtt
xtWxbVAplSGXaqK/ui2gaTeoCcnG01UbYHZTgc6GC9xAIARWx746dI2iuqFN13b2Mwj4ZtBnOQNr
ixpwOFcRXVtc5J6IjUrgs1spubQuoPwo6yWFmtdPyBmfnLk7sWmDI0etQq8l2d6AV72rSbEB0xcP
oiziJLw2HZPKjsSo5c6WdeMUkZIpsBt7A0VGAW2ARz99+8h8d+a2V7Qk/8KPOEwI1F/9JpzaNRap
cUHT8KtJsCApfzlwBlWCAz7sUCQ8nVhlPo4kwvnuv8VCbDD1l6hN2kxnS9Fdp7Hr2W/E4KYDU1fz
ypVTTlVKdhJjE47PNazlfWjuP9xxyzewOd670aoISpsYg+w3b2mTxlrhCjdy+TZvEwX8QacDiScp
JoeJK5q5Laqq1qiYd5adwv8fWMOCBBAC5VdnUnVb8PE3fVqcfVt6LXMLIT5gs+lTmBDc8oNmpOaP
EYsTqp39x/zSIY0NsaTGp6ycqEBHWXp59LznZBDt7MZcZq0x0fogk7ZckmNsfurINwaXTHG+6jTG
jOYKxuocW8o3zZ36dewDe1NA19EoZn7WIKH/NIYx/xOV8thMbMX7Vbe8dVN8mCJvap8nChwKFMvt
D2SPI1xl+qStFzA6oKu83TO3UDUSBsdNliPr1Lqi+k8kEA9rPmGVxt5Myq1SilcTHYORFNUyKAnd
k/b5rw1wZFJ0BqQbEpSgfp2oCGhV/OLulbYQggLTmmgjkjjRVe1C096y2Kxn9c6Bmu4mfnfQIa4J
y7C7hSiv3CrkAMAxdWNdtd8VfHHf3H2eo0o6QLYjpDeUFDw8Lo1rwG9gYOWs1tLmefkcj/eKTQhl
kbUctS6LkmPLjOHYi1eh9DOt6gp63JS0yxfmgbocdjiPxaIUoGzCdgweHHivV8kMIE3wsMvOdwhu
pBBQWc+XPRoWgWTAKt58myLGLDQky6upISXZdELOWzvf7vFbAIFkBEGeekpHrg3VPjivelmKPXBK
dpXQWJlVp3PIesiCoAubvrpOBM9Nz5vaVN11h4fpQOZTCZOpfgpHrLb80kwoMkn01zAqTfb2a+Yz
8jIjH0yplDFr3pYspa7lVhvTI4sHwf9keO5DXXdp0kU0kAbB/S0OJssSIvJ68Aj5csUfuzb/o4U8
bBMv9fPTeA0D2s+uyVSrvUYjB2NicOtqXaTnW4azMCdbRHFE+jFTWQLw7jjyDd96yYQISDPG2KAF
bMu0kOIoYiP7t0mEdTJYqaClXxqvZHJfAcVYUCm8aLorbgWdyHmRcdmlUzgJ3Gjc8UCtzNd6gZzV
SAvDDlwCig5TfzmdTk+p29d9hBgLMU7bYxylSqYGzK5Y9DU/3iYtWG4RV9nOzsReAVcq6wUKP985
hu/AB8REGZtgf4iMjwP3dzTHnjiOgbMAEpZU7tdC5n21OSnWRu0u7Op1AnfeBCf+mhoKfOmPJj0z
y88fWJskCiXfbNASwaW/tF4E8c5klc4kEI00KF90SQ2q37kY8ebh7Z4ylbbzTHtKLqX2ONzx7ZlO
2/Nu1LcvG50E0m0mII9igHMmdTF95a8ukB3czZW6omrIzDSKkcgmDslUIDYNxlkEt3ACbZQCj8vR
sHWqiO/Y69p0m61f4TRr34sY8ZtUYcrAj9EgxZ0+jOlVYJuCxwxCfsw5Jo2pEC+QixWXf2rUl0sG
ENAdBxfv7UvCXotChwAoIdpTZJXL0zjEggmvmkdnjrLN+3R8dqkHYjFBliLjavs2sF50hTO3qDOd
blZyC4/7gvJQKvmscpEKortSW+5U7OpiTI5GmR7ck+AGGuiDgn96A5BUeDrpu/omsJW4U0sLCvA0
/cjFxpjLxL7b/Z3hAI1wC7Sq3OxTl3aV08WXTOqwWyZ3RtGXhppO6kg1G1GGlFTxrO67VSm/StZ3
4ocR9F7LDi6uYrkSjPOkhNZVDuw1py3JuFBOEs3P708GpT7Q3vTz/GT5nF6A3C+nJ1AgkJ+wQSR8
djIcTY9bbQBA8FMTk8UunxiGLYsB9pzPbqAZdzgP/pB68mM+O2KAKOEd5iMkogl80jrOdemIUdgS
wV+B6b1fbW91CDSkxs+Q4fe2ytrb5u4zQaKfL5v88QkT1IllYBnwcbbYd6EpAl03Qw+qmorBGpn6
GSepBsBFMUg1EAL/0/JivJFnv9gqqnzNj69Pp5soCBiFYHbqINXIx6FFSKue1UZAv39TveNAmfBF
tjjv9N7xydorRZlfC6Rucz6Evqy4xVN/kfLzRffNpqmXqv+psLe/kVDY171TIFMhMh42osKuEsAE
Hd1988tFr+o9J71Ug1a2T7m0WP9b3Q8eM3drAkaa9jPP89LLrJQstZfzu650G21EH31x/bHKTA4C
hUVbMTwBaTL84For3gHtWMZ8hVVtEnRcv3uCNfQDYH4vZNgzfDLmzEe454wxJvfIOZHDpzZoSgLs
DWns9RGYxLxMR2mCybNs+Dwg1BhHTijoYvM2xSc/9jEAYmMT7+DMWM+0C1Jj5qo6OQIPyZtI1Fw5
g1k0vFNC+TIVTAa7ZB+O/tsrAtKm9y+HsmdRHr2J8MifPu/rSj0RUTod19eBph/ZXUqwyTRXuchK
A4PYiJVOwasIXR3tC8Cx0KJnquTxQWt1PbuoWGtROJT7pM4zmyUT+pjl7R4ZLZ3Oz2FPjiHZeXtc
sZXhSjn1Hgc0eF6b+kBYV7jyt7gQ0jT06SUIjQOWg4Y4NDmN/mQ1P2Ylpw7EAfZy7pw/+pmta3iZ
OgGqAVSeUsFxCDrkQcwoqaCZ3eW4ffwXX1iXpcT0njm9dURbFhR0WF/0UrinEfokHelduf8W0v+e
Me4DSUI64raIoSo4cveDMB1M3LOWBg/XiAIoDubdR7uqDDeTLddekezmNzcx6p9bPX4TBXcY6TLe
ZLqRvTLtkAJeLH7tYGqJ9MOkZHFFpG1yh0ZZ1t4JLpGJMj0UkGQQs9kM84hjl0l1+cIvybj3fqpx
PvaU1zZ7RhYQRNZO7OsRL6jEbi5CcZYEHVyAy3uZODa0Oz6dY/+yoHbqpiGiC0voRK+f7YlG7C8o
1lxHhU3MM9iNlc9d5r/OZLiItiYc50ES5c/jR4WzIZN9ZNouTtLEqUtBrRFuXcg4C3VFKio08xfk
oLpriEukzGDmeeTBeJCrpCsKLV389lzAn5z+XiGLDMjRF/SmpmgA0NOi0uGU4YUpX6ZfbMxi4ihv
1RD1h+Qvw63QW3+Pa86Hgqjg4M1+nldkPOhXsYu1k1u6nGcE6PD1UuRYmHLxC0jHuGDK+Y+9ohb2
D+LvrxDZCd3TXJuySts3AgCOfgBfiADUiN3DpbWon0izmj5155XUFDteMzUQ/sIsXKmbGq1e1RPX
aaC0iiaVPCpBr9JMUkxJzJ4sTkUru6Wpv3sqay925zmPoTSv9JrChdq73710veLB81J+TUqqtFwS
y8Pugr0QtM1kW7QnrZT1ch7j18OZzOyxYsxGTh/ZTCAB/et6kl3osGa1ohn+nJUom247InPXMyBB
Au4PSek5vqLAUGwH578gCOcGQxk26ujDUhHoXsWwcq76oDPCbq+7F3oBQqPB08o9PiGYXuuIQO3I
tnNUIFmxUhD1v1fNoLm5n/0KkFYk6w7AOfbJroUmFbMm4jwOyZb/SodXlpfPZNRGehoMZChH9VyD
m3DPys93hmYIGJADw/nuvRD7xGg8l2Je3//YZBy6YkgVm0eufW5rm8a5FmwolSrL3iWM1qKMngbg
FTEJtiuoM9dkMkqf3QxzyDgDX5Xuus7lxGtSOWnzdsVT2RTZ3UkfUhVc66WLudwNGzCI8BgauUPK
L3ALOe6Bl1OjprMqrXO26IV5Puwz5dQHod57RzgOEnJM6/u0jUQd6zd+gEzxP1FSQd8UK0QQ2yWe
nAFTFzYrEohRMbmz1HeYh1CPza+gADsD6GbYpEsB/a6yUO4eM70AKLm+kD4mbVPPpw4S2BMtZno6
If2fpVoP77fFieLAqoHpWlWZPvhHN3oKBWRpZ8FiPioZpLfzGzjPNo2j8EzM2V6sLn1kPZHSRPVA
0WBcmoHJMYmQv+tnBtEll4OYbkGQ1Y/nJ187wNq1TVCAu9cAXmgR/v2vnnocGf27Gff+edrYnzFe
NdfUP/iGy4oW9SEzzFjKzY8h6uezhCHxDKilOZ//Imtll37ywTfVUfVWhTIhCh1moWSOsF6Chiwj
An2DZ0GnAungbF8MMB3hsL9RwnE2HhIw59Si8d7+e5nHQxbNs0kukkij5xvJA9Onsvy0F+00dDgv
Fb9JN8S1iz5MxiXHySp8ISylg4X2TJVEnh1KuDn4fjv/a70lTVTijI7g658r76U8Q5ihoYI0lQMt
fC8vflhguw1vJU+/JYG7Ui8N7GThNYoYrxTbYJwQp1Eon8nuQNREWNqo/n267kxYNb5zcvTM+dwn
RnjKXpsVGjTkh+YglekNNVPfT1g2xYX7hqMZkk9osqLPStA7AvNrdbb+c5wpDRm5B+fHShDVseuL
wev+JMCtHxE/FxdiPB597FUb+n2jlOnHoHvgpLLCHoWY7a75MmGWDCkEeSqbLz+Sj8JR8uUOF+Q4
80nj1SwYvoLFEjtxh712XsPG7P5Zt6+ASZ2MvWObLxIF/7aQ4+FLHu4kfB0jpWoNo19RddmIXxoB
UAYgiiUdZJ583PRedD+w0hBlaPa56Mvyhm+72u1mFtA1cRC/nZDukmFvhAkNZpUm/4S22tT8fXN+
vP9N+47b8XNx4CRwFTF5qeVqJp+vvr3Hskc/LNqyv7rDgH3wExO4wF9XtRX5iAJmaDOod1dwxFLT
h1eScOr34KW0plVrO535sV6MrPf+E7e+M0o8TgbThN8Q9puRkssCA8BGdkUXKUFlKt9v9O3pqjZO
Dov1/BHqBCUHrehNVZ9ek6ih5CIbhqd1RYOoCRGgVwu710EeNqz+IIjYpbUpXtJ+TSRSHzdIEyx4
BZbREps9ROgNRfZec/GlIMFKgrJEC4OdqKslNqOEWYmln2E45qGOcTAKfW95zgcceBhiUeBpJ3uT
jQtLT12DmymfO52KiVZcF+EWPcslnwuz5eYZtA4jjJv2c8Upx5/5QKnt3Zkp7k/cAMIg31uGtov1
FC31jP3Q7gOfvyeYAIRVgnDepL1fdu1UoBkDkGZuXvFAUnLFUqQ+jt4FHwFmLIkNQkA04yIbinia
0t0lb6rurUmF6zPx9gnZdgqrIRPtWkH6g17CAjs98Lmq43IxmwAnw0VHJjBWLEn6TDavjPLRTNTr
P48bHmRD1UqKgIxQbnTOXQQ61V13japIj0D2W1YO7r9dw58fpuT39j7XOg0XIThmPBdE1zeZBAEU
Zuyc1qLe21OHuRcpRluyXWelgSUCI0+iEG7abp1aMtyLQN/Ei3Akg3AfloNIjd3dThaLoN9Pp1+s
n1i1r+iFzFvE+972QwB0D7K/6qd58AftiMYFLYS0S7nHtA/Nwfx4yU+U0qKb/oi3DX3J19AzsQuL
8jHeDgzYUtS8fNAJrIxakuSRRemwyAZiEtmTUUUwxlPI8J8mi0Jbot/42Hxu7flneIzBbbsMSaha
mGh3IcyUOqafWlOhhUsAsI5VSdmU3FxIQSVdpwFhVDjwB0CzO8TEdDbgb6yAZadI3KQzkV7CdZTe
F2SaHb9zTsseXd7uMpjAzEtkRFw52EmBgXstUaaLFkkdt3PbvjPe/GnzXwsqczaUGCqVQHDAQqw0
paaWQjBHtCBNsbNeiktW35RfILZBY/Q5HKeBMPoKHWXDOZW+BlxlF6Svolz8qL5TOXajEQbkX0Ud
SfQwopKG/8UBG8DWjZyD5eYnVHjboYJbTLd4lSwy+z2j0D2tx+kItxQUApr5TuItNBIZoe6RWSTs
PLP1jdtTPJZ3wDaA5BMDZjLkYA2WzaJPI871r4lYkZkA1w0CrqtWvodhxMtTHbMZWwf8gD0fUXWl
dTwuwXMan90CvNpTh6b1pVq3Eibv8IuaA3R/eSgb9SfSpqZ2A1qk3jiINBs8YixX0YQ8am/QCZtD
Qy9W/8ZAbfo5IrCQneM2DWMcDqRQlgZIkeYCKQ/dX4hJ8gBpP+BXgkUWavfn48bFUWjzPdUINPf+
pRNJBccQFoOEOC7RVkoCJRlIU89YVJ/g5tepIt57a1s7DOMXZIaVuqkUZLB3/+DCmHzGDRpm5o5C
MbNr3UHDvUL1/FESjoVStQgEmg2Kg3scRxW2KqTcCnr9x6jrHFA+CIpmGorFL208/DzDZVzl5s+T
BzudEnMUKeeE8NiNcoatBoPQ8nFzqgiBhv1TifYGVZawOYePvHDDRD0FRV5Yb6Ss42U3PmOqv3iz
Y+ktbMYpixAbUN9lD4fIca+DuqCbtsdBA9+weMRoijTlov3ON0uJoSx6QO//SEk20QBoY0O87M2b
kDr8ycjPGYfl03BaeZz09OGmOhT/1r0qZs562ak7tik1R2MWii2aSoJMdgWEtA9uQN0uebLaWGtb
RaV6PnC2lG22pWQ5vKgvKspm/tiMWnGTVLrTTUJF39ltHma8khWcv9eMoZJag/3Ra6f/Q2ItyW8a
dGRPQHLWbR9jNj5n+1E1dkS88MWgWkRgfaoHtmRt+fwbEGec2/ptyucs2ltzfwPtwWfRWuZ3/y1p
Q/p2FJRvRScgBa7qYiYvObZufHhaRkZ7h4DdrSVl0H0iPVfCt1XUNOxqXgZbVTKBClztdgmL1lEd
hzl6YtVsHAIlLM6Nak/9M9SOuP9jgJSJUeCsAFHj8CSxmLBzSBdJrODZp0naIqA2pcXAukz2BgXr
rBOROSObLixbV1XtafX/et0/Vpre2SknCGujaztvuG87b+8QVo5oWoTHoFu1nzEScyRBnuazexWd
kUmuvgvbCbMlog+UkWd3rTbNJoq0pMr/hYGEgD0y+40F6xSI+YOGb5KDnwzCDvAdjstUqCqnT/UW
J6siXGTYvJT1TfQKr46aE8R6tFg+kezmXK7/RO3qgikktzIpjcxWFbHlBLgr2heoBQXRb+lXOl4W
+EnLKiylh3ySpU/FuXCzXQNnqF/Znk905Al1YsyVq+qJNtG9LQY/aw5+XweDP60kaPNgxb4spkfV
C+K0GHWnxagEvAYTc0juwKJB24PJNAvoegARL2XfSo+LM3o9dNbJCYHbGSQ5Jjy4eWYzUZ/rVGaC
e2FrgAhIRnev0qONn+m+elumo5f1uB76QpmzfFoq0FQJ/SO3GI/euRrZOObtSU8CPLnToKQqes2s
pnqk4OJyvLy73Zd3SjRKi5tvDjs8JqzGzK1049/SY0Z0ShO1TZtTZB9nJgzuBy9K/lhlGfxwhDQN
pvw1sJRp0TM8KTy9GNG7SydKeXFl14GaqQGjDc6txYvXym4PDORxDsihcHXsEA1F+5IMSrCSsH3R
uowf/6EOyBP7hB3kH6z3PVKEt9WcWZn3FTDqeBcP8e2ooQPdP0Ge6+hW9Dpiz0NG+ywhhz89wNeu
ycTqiCJIXMP/WoAKDAmh/tS4HFhfQ+eQoZyuJllf4o029Sup0QlTBbHXjO9EwkPuBrBcVCDnx6cK
fOu39McglFEDsFaVPLowU/iaCmNczxjFQtrGswbKD5Q61Bho+Mjm6+cyof3Zx4NMnVPpnTmwyvbR
yg3PHiAhgAnklebgyhQff6kNack2w3UH28tXHryPMyFF/TGJFEdyLjNMmHdknW2E8iApqEnK18Dd
Ig4qGNf6l+rTdLiwsdsJVozCDVP6K6ajIB5+qwPVr0uCRzTsPhIwAkH/18FWFgwF6tS8T7PuJNgK
ZFNFUfQvDRfazAsCd2JFHSht1ssqeUgmoCS4XLgfQU+hoyP23ByqHUlfDoEsQLMNUl7Cbuei1P8e
TgojYJsR4laNq3F482P8yD/XYyoDbtBGeWUn/tXJ9wDa+iqfbqYZuc12a7Ps99LtSvprLeV3Ywqx
PJWoCFswPyfFheu97JERgJtKuTGKAvalQMHmMwOjNPVF5pm+5IeB/hKGqEw3JKo5Owe4UDEte9KH
CCakP9CMBhNiLVr6yDB+3IDGMlKxefzpIIHMWrXpdthbAwTiPvNQQAdDjE4NLKN95ZzUnlbHPVF/
Kj3C9l1KM1Uos9v/OUGRM0UFpdm/LrRetMAtom0tLKpqoJpYI9ENgzJd/OJVPjL/mAJlK7dqUyW+
VezU04RLxb2CfOydVuIFc9IdRHAXoPdX4V+2VGaz2CfSGj42fdhUuPyTDsiy+rZsB7e63xPPHqAh
Z5a7OqqZcXe4alKz+up602EdDwMwb+0RuZn/15y6fcpKEWduDdykCB0lAVVvZzuAJ9CU0QaBT2ei
vwAWJwp7PfFBtt6oxdJ4/cSmryGXUJjFSV2NesxZK6Q7Hngt7PBarccyAulZYPFNUG0SIGWjhxHz
VyeSTHryzSzoT0Tfs+tt5O3Pu0P9WnoptM0GU3tdAk2i+EfUoZ7icDPHFg567O6y0E0KmT/F4YH/
YgzEPgtxEiOUVwK0bNeNg+orLoDcTw/0jKdhAV9qtrLrku+4/lvUfTGAVg+/rbnyh129GsTuv+8z
LTBqVmU6Sbsfmgtv/aG1w9+xq9nrunoY9/qwMkDTucaZwDdB0i0dFzgEjotRpDfcBfz6UGGx5pwn
ZzKtQL8W3gr6iu1fWT3VKKNaEIktgV2CTaBbkugqxYeTg6qmB/Gl2nvU9H4JtA9B3MYV4UdNT8nU
VG7N5+8ZlyS+yN96CbZtDqfZ3PWrMdsqOjmy0ckET6bowTi61YZ3ZSLwHGal3B7QPxKq7j94uL3u
4krUhA/byKQzaenIxdrhbXc+TkQAacrSdyNrXnfwpjXm+g7UDdfTg5wA9qmFHPJIcfs90oHlqHmM
eWmswqgs3LP2ml2ryW26oBgFW6lc45USeE1crwFVclcywYL/6raBZGhH2DudjnenHiBgSC7WJAt8
IJqTb/NFLEMI6gilCjs0DQVD1YH73O4QtOkx2yBE8KYXQVw2xvRLTgrmXk1tbjfl7ebCcyraQWSl
U4XzBu4e7AtxXCROf3gSyoSY5Iy168iIPB6WDS9K9nWcZg8bcZVtk3XJ6D4wUrgwSOdmiGLRtQW4
Xz/IqOQAB1/DIlagjGv1RCHhFXcmAEqGRDzo/RrvUw/6URKhE5owP5/xoSv8anoI9RJJ1KAPoHQA
1dXCeYLBjjyvoqRKUVyx1ie5eiRHgJlu3QrF9uU4WlM0nPetkzNEhKrC2q/Ho0f2bMIjteaJoWUU
YJRoQWn5MtqjzG7OGhETC/M3ne52ShJKf91yb8xYbHwkiehaEFBstfhyQp/tvk5mEAx1r/vxuU0M
LxzSGWBSkCkoIbvq6tXgmZ+Lb/RbX3RnKnC3SHZmn0OLyHWB4r5tOLQigkW07Eup5SFQUmVDAWue
trD+R4y1YEdoX/sV2BVw8JemEQGoyxTrq7txNTj1T6v7IigmbTwvTp1JKmxIiNIpuaMsvhVm9sF6
cnSfyvTBOm4EIuUbUPAAWmqT0RV3WM4h22v8FaWCz5XfaAEAQdLwzeP45DnylBOGE+ywD3EWzEVI
nler4nQ6KY89b5JqRQKKCnzOrGzYPELQxVPkmrwXlUmD++/OIo3nub9HqSYKKZ/W00jOdctoPIut
/Hyc4r95pHJ7RG0YVaaJvC1h0oaujHhVVL9upS9kq38HqW1ex1UDPcqDZsreQkpVRXbGwLxVyplk
+QS6KwhWPDBYo/RoVl5iHuIcib+8uMDMRvLva7Ly5litPmx3or84gcmjkCyxoSxzCHfTVErNDTDh
XP3DRS+SiLHrXcYQsnRX36/ea7sYSWQPYpMN4kaa8/wcaHXQor38TqGgw58s6bTsqTz/5wrfdEVG
AYCtdjhj1FWvVjT9UufePfqapTYnxgkJ8EUEIQlt5jdqRYsDZ4nUog5Mcm+EXdbWvB87A/ShFrCU
Uo/wDpU9+NRIWlrgTAeZ74EqSPnenWebSVM0MPEVA8kHslUg9pzDZ8lV1NS+1wz2akjX3PVQr7Gt
B55wApvSM0XeRL8kmc4dAmHXwBAWpkB+js6/IVQcqn7wxanotolWvROpYH1poVodUsB5cUyQk3Nw
fZvfkr/gwhOEBkzfWQN6L2KxIyXdkPEQ5gxroiULjOAFSpc8TMWU5xvCa4UlFiOP1/62TtASoFuC
Rknda9nphqDOPwhVMmNaNADq14OKB7kc3DPchltqFSi34DoUqylZVVJHw0rghS8tP3AbEvNBegHf
EiJ2D4C+8mcTZKPOpcGXiD3jMrJkU1Ia6Q4DVLAEH3MzpSMvazx1RBlhLc4Ivx/lBz2k9KqoocFH
I8lc/SRFdOS06PLBJh0D9OAFX6z90FM3YhEBdJiSJGi+lr/3bEFHdi1q3LvxR9NkEbtxEosOumtr
n+4lV3nNjz25iyYih/76fmtsL/Sg6i/daP5xP7KQ9EhOT6xVYvL2VjjWckHUbEATq5ysdUvS7SJa
Jo3LWYhHcunhIn2nLoxQ9SLM8WxVLJupM45soEepYhhka99haN4Gcnss5JVnp/AUP/zJrvxyQEgk
dbUEOQ9WQAjiuSvn8wYZ1+HjRtG8N1GChmFYBgzQWkJegHYxKRpoSuLqA3x8nma2H/T/Fk5nDlrR
/dBnRrb7yUXPSWMiZssfiV/F4cz8cF6ualwL6SEahPaSjAUgiULvkIuaMSnA2fCwoI9KRo0PyLJL
V4mzgzoBFXw4HleH0L0yCnXSMpqs7W+TgNZTPJ7sUpCdzVqsLBLSH2QOr3Nsg11F/iVhR6wrVbWA
kTCparvb1xATQAP4I8o1T8bnosqoFOzk8Y6rIx/lWqhJ2A1hUNCO1fDdm8WACybt+cGjDkPstqFJ
RLjT64yOXr5zDjQpwL/Y1J5as4Kv1iB2M1TkJ0TfIRFE35IYiFjvY2Qvby/48rKBvLx0afNkfmXj
gVWVDz0mF9jCgrsxSqKxbxr+6Ms+kUA20XnlDnzpN/goBL9mPIi52nrHjvofrPhv52dsCCHNayv5
m2WfeQseiTl7j7kSvtq2E+F51lMIWsLfyS8COyPWpk0/sCqTktm0lU02I6WtO53uKhAzY6xf5tsI
fhm6vbT1+wV9WaLpuKJacHhZxczxgnW/XnB9AzJ2MrZuX44LgrDzIJLKjvrydxeM9b8ShIMakk0E
Qzn9OVopnV5SqjwU6YjDHWhAusqb9iTtTdtgUQSr0Y0KJAEcq4Tlq844EJ/l56w/0ibA0bbaPLG7
wZwLVzaGwNKJGKbwTch5LK0mAToEeJf1by88mKuMQllRbgNH9eVrOYZFzxoA8cQrVm1I/CzVebaL
PztLg32njXfKv7hGJSIpkcbrQgiaKcUvIIxSZeHFDMh5NLjGyEqVunq7isjDvXnhDYDMoXSD3qI9
7uklMJwE/wymmZxfoxM54M/Oijtrb9C3G4nFWjJppSKPF0ZUt+/a/cj/hJOYmHiFIEV88vXZVaOt
2h73D5kkWa05PklVNSo9adoVY0BuFIlFruhzCG4OE2SuBrERNWMsPDQTYkPmNYwp0MzcN5cSPq3i
Vi2IQr+lb5zmmOa83zH7+04g6BjqpLyTT3Y5ReLGV/0gbLrkYlISTHGJQkGtDx+MafLRx04cZQ9z
mnPrYlLqx7VVjhYeqakARY+vixDkB80xg/QW6UmwerKSZly+4N1QOC/dDVv5ztuWuLi+XE720AXe
HXeTxLHX+7pc7T/ytqNPAi/B8GLMFV8CL6pgq1uWQevQBVWbkzyES71tJoTYufOrbslYe37xBdfQ
DeNaqcFKdz9udrFh6UR+1jhu6tvUrQLI5zg2OOeu+Yd+H12s91h8ak/rkO1FbQa4q7oePvnL6mvA
CroZ5xeISg6X6M6C5SkkE4FmEObuG3B7vsid+OFf0ks2I1Vk1fI3QVGKDPRvXbYtQwLCEszt8xbK
IlBZF0vj3t5PvCDxRbdy15rGSusm+L7qE0eaKrSmM7GO90Qgk03vgpQGCqYQqFWzqSQxQc+k9jWI
+JhHEc1nwJLGSiHNHYqDWKOtzu/hFW4kilMT3Fup0t7mezuiRGMJGhxvyLg+FhTV49epiVh9z7co
NzyxQMTg1ngOElrAoaVO+hBuj9m7OPHGMAvkVvZvFi8FEBtJ4X8pVpACAVBICJyMy3RBHIf1VeEw
i5LgkgGBinOdSEvwFjrBDEl+edjsOttijfwfPRNT89Qw+bflJq1b+tSsYSPzjtRNJgqqHiY1xxfc
5fULA8EWaY3s/ZSMmmfd1+GpfcXo35f6Egbi8rWWTSVjoMEDQWWVP/6ydwgOyTNaAgnjLK0V5sfu
qvLcHVAgjJC6/+H0p6fsq23vvdV0enAOAErZR2tUxNYeIdHh96sQj2tq1uRTslJB9jOFqe1lyHQu
s/yeNrJsne2azViqnqsZvdNHU2x15vKvsJl1Rox7aJeTkzK4vYv9scAB3HfPEO1tHcN6kf67rHVz
xSQeM9QjTPVlf2UYhyPlcHVVOnA6LFfLnypGoSMhf2Q8MSQ6Cagz/d52jszyoq0gVScws81Gr6mf
Qfas05bX6R5wJrPLj7aBuG4w7sefUglp84AM5SBL4r+yAyppBZSzIdKrsfqjOxieHTr4e/D4bc8r
KGPEdLM+IcKNu6JFZYI8hI/lVjGDxH+G9BsJ0wdCasWxWKtm9f91/aV4np0wuAvM4W71sVDfbADB
Kmnx84FM2Y0ZgOErVLICly1Aa9JnHedPI1kq0OhVK7AM5BY5wAk5jcGLs08wOmvCqa4VAWJOQGQ/
aETqZkOy9gBLsYCHsCoNx8YyGhWlXgHb5ZSEosx1FvY2rHGu9+XtYI+H5SI9wWKr5vaI4N6W9x4R
7XzuxPHnQlDrfYIYZPURX1wniu7Lc5fLd+amrpirgM22SmWwxfUdG1sI5ZVZyWdo51GjvldNJS7P
82PJlmka1dR+hMyZgEKpUWab7LoV/8jYhs/MYl6cSPt4wM3S3Z6Drmpj3gSLzIJKzqAuO0FQaxna
0n1WCAKZYRxchTRS9JxxTZoc+oWCCu+KWd+CConq3NczrCvWOywGw53SOu9t/l5OVC7n+KiiOvC1
S13hWBk6XqEcBjGaEtGpKjIm5lbmOqojOjQEIIyCHIRUs80yp1vCQMWu7kvMVoYc7ZJLLirfWJ8y
cvL81GvMrMZyi1aCgV+OkZxAcEbWkqTer5cU6RiQONMBpKnwlXxE3VPSj6RqSEriOBh6c46g4ERc
Kgmv31FmMouGRfd5FZGJ/yLst2N6BmMlTgaggaTFI6yKQVUHgYEQ31i/+m3GvJZJ5yeaWT5iAJwl
eaJP8ScvVpntHWxZEfgLge9cqcStwjNcDUVPCWBnMgplzvQbFqPEupxuRkwzLsCMru+BXHuIdYWY
RrIwWx/hDuaXJX5HLf2uNPKjEQqOYRHMJ96Jc6fJavXqOZ2QK1gSiQBV4KNYqkFJw99fq2Rnx5sw
YkBbQvJtvkWw56IurjzDd0ZxXnJddfNthf4l/7NKnuRlaxqcGqZwiTXUujpOF0/npA2UojKbVLAp
iH9O1QEKGiviALauH48DEGFcmI1fvI8wE2q5+TE6PqGnqsSzEf5FiGxGE1dfSGimDLNWqrW+avI1
uZdw1qTLxjm+Zjtd27C1rrRkzZ8WuwNaAO81F9V6AVD06jwTp7xj99xkOr6TxebrQOuQTAai+3b8
QCH5pv2zWkuKVqbL8UCcmt/eHLIC/P/Ar6WnZwsqx3j7AIAuwkrjOZxUj418fAoe+UCIoNNYMbt6
R6MM4G+6DBkpeR5mdKAyzG/bOVXBLGOun9W7Puz2aMcdmZzN8nyrs2FKmYGMw+qo16KtAiYNTACu
ELJgZcbNHRAk885qxONMDqgUnWt1Yesj0SBjdGRoHzzeAC9ZIkc37K9u37l+pYxQn5rdqGrSO0ss
3JhxY2Cimn8LMohRHnRxZjL3GOeudIpin3BVzUsicJD8PEDy5c9123Uj4HQgy+6VXuhosoife9s3
zomI2wuGR5zSdeGAA37jMH07BkO8SNdbmNaFVXyPGCR+BURLl5O1ID7w8cA7eLsbE/45571uHNQ1
58BScLsz6AoSP/Lq186tTb+tuFS10xuu79xwoHm9JoeQ2/QXDUlGqJ4ZlqGK+Jx3e0EMSLmbkpjZ
N3sw8bpy0xw4J0yLTIwkHguQblxy1yOQBmILWrrdtL9IPy1nv43vO4sH4ZWnJW2kWHdhKHBpdvfF
XlFhdkEnXcAS56zaSwCs/mh8BGlKwWk8Z91o8djrwyh2nUPzRQpix8f5UvTVyCxndkR59sKDoIh+
2fLNtlNQiw2C5j2BkZGCIkpFh7Nms42H/cnz3UUAmmQvuDF2yqFOOWjEk1Zxh7IRAPoG0fb9dpDt
r/P3qrnsXVaZgQ0AerH+iUTR7rJxCFmltKz0PEb3nkQS/ju98CcRw7Izs/m43H6WjVMK03W97XBg
8bXDJ1rGscbkQtoPQOK1km5yh4AQZQ8TOC00AvEuZIX6FcqEz51G3KMoyATSQGQJplxObC5vBxXf
flNkSYgxnJdxTyd8G2Fed2DmGxT0H8M5PW5Q42OvZKVRCvjOuVuIkFlabE6atwFKa+onTxxteNnk
DLMPRgNT2BNMxUvt+sVM15OwAROSGAq1o85BZ3zovKtGkF9MOobINY/5XmxmGjlgeAbh1GgP4/zo
UEv01LwxcSUEG5RTOyGz0oZX8yMHDe/Hk3Zeh41s1bKHK12GvEgvgwkBxhUwJi6oQrX/kWUo0ML1
vV+tqZX58viAJI5137uw5Ux8RPdhXtQfdygFzf6IoUvh3HQjo4eRQ2LvBPncIftiYMA/e0beDQ/z
bldEU48izCmuUsZ3xgWjXLi8Ebfb9FtD9Nr+WfnMOs0hGj9Tvh53qSd6fMQkGjiNs4C91Ux7rXkm
nkRYB0dL+PoMbKR2/XMTC1Oqaq4m8W+L1n5wBBaESvqUoXEBy15nGOVjVr1SjYTB3pvii2zMOOoD
3X+q7JPt0TWo3bIfjT7ZWePOzoBg7NcBCBdCGOr8+5iTQcSvvmoYr1A/oltS4tAiwVNGBO3vPoi/
Sc96UxbGrrQDJ0XF3h0+ptaiAyN29ZwD8rn941NJxZT4zvflbkO99J1jm/ktexg1SmPkldiZS/ZT
oawI3d4lSWKMDuH7HjC9txI0k4x/OkcKytM4e4QjE2M2wZ2ul7YUgU+zEkfKH4uOug1NFADMfAOM
/y2RWfRVG1yPMDqvsK4egz/4sEdS/BePXAMvvYCP8gjACOgLxbNtnDI5843PTIvueTn2MXXOoTFn
czL8YZGH4ghKw7cNbNuzBYil1ipgwhVu5tsNJbfAn/gp/lPlEf4SOalOSJ4T6ggNEpu70lcwNp6t
yo23xPMjjBasAOl26DBwzO13jYPtAQsTgrurs1J1Qq16A6m7MVIxVQqN/72Ee6c1ruvQOWvBGYsB
wmZcasvhPzZ9q6KaPCqOdskFbm5swDw62r78rk0dG9oYsouPkG/899BYMtIMBti4cQGv9kR3GQH6
rUk/Rzh9Ola9X4CxLeW2QFq8WSx2WzwLa/JF7qy8pa0sV331mdX11FcHJdc8838m0NV2Gj9aZqvF
x8BVxrqpAv/N6IIRyMwZDmcNaskjNe2yakcAe4+506qdBpAN1W67+kBjFE1NYrOpaaWLLWt0PAZt
zrD95/ZIcaaspuz0yccRtrpZAS+eIUgOuTP7YMXjBsravfM92JSs4nYmH6+pCxSBqET3pUw4WpK0
bix/HrpT5W2HOiZBTBKih+yOMBAc9GeItQ6K6qLA48qpWz9LsfcX2Ob39L+BHP6uGckL+meBIQiq
1Xjt1M0KCxF4GgyY76XbwyKTLQqL8DAvDg5L428Pb0vzb072Vj9R3keNJZXaIR5OfpspZXlvClE+
dnjBotbeKyrBfNo4e5hZ1hT7mNWHbjhZd5QF4N/cgJcKXVTC1bRVnpFGefaA9AuL98llEDA2M5Rl
49Y3vg9kiGcQScY/KB3wgPxZ7PrMzuE7Hnq+QcDB/SZe9vJKXX4gzAXanDJQkSunkMRNs0NSXO8w
N3uSUS6Or0HQHV5dswZ8YBOoszC52ppecmxLbP5eNzfRu4NXu4jq1F7fA50fkIG0VHQap2xfYEol
tCh53i6HZNTUMibtumSPT36H5FT4i/aNjreJq9wJoLhNBpUvAH8KPBEKcoO+nPq68N6hqUdfAmj5
4IU93C6B2wF+lUhnPuDACJNCj3k7h+TV3yJdDRcLRjLF+z+VDa5de4UhgKOeVf2bZ2bOAffiu4Tg
3z7ickg7L8lPqzA8s7DzUQodPPLlQR1QXBPmnFs22BVkFegSLFrMsqaczPub8Ug5ypoZUCaY4WWX
PYzbhIrgcVIiuX/cnbyp7/EC0KXQ1nbXbLfyU/1t16fQJoVn0eDM79nmLPk9+WlVvQq5cI4FnCU/
rf8gU5WL7v3HjyCqgvey92YS7YePi/RgpmnNOjc+QEu5CnCc6d8vouu9D8mPzn8Yx+4pq+Dq8ssJ
ENc7GAOOYzYz7d4K9cAOFapi5flQ0qOD6pMHht0GFCzhotIhgU3XyHWky8oQPtr4x0Q69HKkx6jE
ubBA08O2B5DgQ2Ei9Zrp4HqEBq9d/kntIlsu6BugFvOnrtMLtguhfMiNhfrjSwce35BFtknI0mB6
fZCbNQtfnBwWtRRgZpAiY5Pf9tBwm9pBcpywZ1yB3QYKYL9M65ePnZdgBMMKOs5pv82vRtyqQ+nq
PiDbRXhcjOAhJQ+XiRFwFDZ1sZK16jPlnibSA3YfJkf9QZIoVgbY58cMu3S/Y66Zd2TGtQrvS+m0
JaC5sSvebtZw0PDgsPnL0cMygOmOH7+wUo+QHps5I0/SSgGE5FlPN3PVu8NypTth6v+aDY9Wjftq
0hBzfZo8JEDELdDiISvcUxLDgx86YA2U34eriC5fApI2IhqJEEYJfoVFHrXxJ5RgtPX9cxZbE27M
hhQSsVju8sOdQxRiFjSDywkjoWb/+0KlCoA9HUfv5T87vqEqObKyxI1qQwm7XnElAqpulbYhXbA3
KDepFGnWm4ltKrrR7EKxBgaWlP3Up3wFJAIbaTNH8807wh03f8ASVJ/Zxjwdk5+muXnT2dlDfzZf
PM4FGVf7812XE6b3d5hZL+62iiB9Dke/pC0253aOTIGu4HWyYWYTUfO1azGtdvAgsRUADKey0PD8
vvOuO1ZW/PWaZi0hPDjnUWqZPQtlESgL0PxqWBJX5ksoJYmUkicfxfO7Fiu7Li//g80b8MvPnfn3
yEakHEdnjKGR5lk2inkFQqbVft4hd2DsFvtx3xzvMRk+ZQZF4RFOIJqzy3xHXgJVCSpQ1TUM+0bO
vyg9RhSH6/98IDxKJgBj37MGrsFyC8XuUzC9yT02n7kTbMi5B2cS7i6Vg9W7GgF1RlWOfTQfyCSt
O8peGuqdR8Bobz2rajIQOIP1Kpuvdt4DYGyxNEDqbvuYuWMpHg4WwUv42Q+UiT3mkui7THbqKRz1
IGpnkikB3ChbWc+7RgTcAuZuiYT2Ozqwfxrh4BmuDRJCOWwIxY1OzykPpOeA5sZ7p3HbdLH7mw9u
1Z/KeARtFd0S17H0zOeFDX1ZhMrNt3dmPD3NsXYlW1vZDpG+m3lpD1Fk6rJxqbxaORztoBn5VQZx
RUFBQGTXtQtUfzpGm36wq1v0u1KAGbzF98Ov/bkY3At0JLOFxJ0e9q9aEYGdUJ7DKVAGAcvADdbc
kTrCYgxVo/SZgVYVSoDedk8BBKsgV3caQFkoncxBjytNCZ5ZqflZC+S7OqRttkEm36ivoT9AO8fQ
3qnbGdnmIVafMVaa+n1eEjhjGga2L/fPRsDTCxuYm0kmji7LIvtoA4K4UeFd/qT0/dBtpReTKDJK
yLd2k0jE3KtCnKyoxtTFsC0LqnMDM44uvDc9ThO2/YXYPakdtY/OauQ+VW4x4FWfZQU+KIvckKuw
5CxIrgeAkPbnwMCysZAsngsiv3JE2WEQmC2xNbGjqD90CkNugx0J9GlKzalD/ptgLznfxKe7502/
vWaKPlBfRRIcrTkktLGTux8iPqhMrLewgi9N5WDCXmPOela41km+xUl5el4R8QXn8IPSmC5ccO9l
NlqWJsOrsQQCL+c3574ABu0F5MXY1R+JOmDYzx6RuTAIIW4g+lXC94HOYb1vfF4O9wTiNxR/hYgL
o0iPoIwmiiVAJFpQB0jwwiMutHKsA4zCIRWWbvdERsUfHWMJKFWDNGCLWRtSg6AHYnEhnDGLrRtj
BKeHiuiq7rl6t6u6PTtslYxESoBuPHmRzLqeCgLxqySia9YFVwsMbJhMDuw/r01FXl/Gk2oBixki
jTWNkiZp7H9NCmWMztwqLaeym3sBvKbqQoUDMSbBoh+ofAPu6epiEFj6gYSDnh57WObL7uNHHRN/
YBRnTCPysSXwkSVXqb0kX1KyiapHWMmNuCFtFXW96No2Nxhiuvb/Ot06f/xLgT4CijU5vN4WCMS1
uNHN+byU81AjX6vwM7QsmJh6su+0ZSkwzu3F8iTYhfogLzdoF0vPs6X+UaXUZwsjHgFrKmTXmlxb
B7QyaOXzQoZIscsnV4CdcQk9ExfJFYidyxZsdiBC1bL+tnVaMEIEdh0zcgOghNsIh2XaU0Ycw1XF
PptCHXc0zU8FE55CT8yPCwHDSdiFNZTW1/l7YrJWc9DNu9KDxL0Q3BbDdq2mRdzWUI7kCxz/k9YF
d/qpwDScCYzFasAVLSqjfgdZ+MQsZlgXctS4+4mzuaOgwdaGT7khxPY3ZiAU/HDBAAAOJNDlQQXX
omZyQzHCYcNIX06rwDAozBw8SVpVGfa/7tl+95amsipyR+C3blXpffcSGQ0nsnNquvB6IthnUBPE
a/v7gzoueV02FYE/azZNam5gy60KN1XtBzfHlwmToOT6Nz5FgiPHSXxqHkX3r308Iy0l+pfvr3IQ
zX4Ho74qm0xYucLovDhIMwfLKM/1ettEC/ilJNCeXTfWJWLobVxDpxPJeNUbbvIJDX8RTndCUl0O
rICavmqGUTw4WcXdXBVBJHeXInOeTbalFbeQwpjua1gmjb1Vb7pR6rSVvrZnotC/cvwbTUoS+LKe
Cll+sBxfMPxpaSkwkoJ2mCWic7qtl3Bg4Sv37xXkZzsHA1LyLM+mVgY6UJ9QVlo+M1MO58lMed2Z
m3vqvDjwWRghLhc0glu4PhuwLhmKg6xSUrkb1mf6Hz4X1DjgQBqf7k9+1Jb81dijyHtbe9VtIw2X
JUiprjtHf2WvwPspKhv3ucEQD3Mh3N0ByA9vx/i0/NKQRxsoQw0viAIgZMt+hxnvjS/yxF0ZM0oe
4VzGsPmZ5L9v5P7vLMjnye4JFNLB3WsjB5Gip997BhBDJzWamM5yBXHvbmgH44LTVokrOFCK1XfZ
nla1FIMxLS6/KvfuEV1Gk8qiL9Mbi1zY868rM5Z9LXUI+jgeSdivEWye2yQe5yHnuaQmGFa3U+6o
euasDyeppyv+tSl6SF3de0mLDRo3yCsfEXiSIYmZ6LE+/OSAYH6OnqzMpOyB78SWKDAYzy+l/3Pe
3IbDQHhnnD6owOk7r2jhOzdbplxVentSIwzhKdk+TRw1EgfhXYO5ABTVVt1VHipgkZkrKy/cBEun
zBfNYxxpQWNufM78XqkyiCUJ6r/jR2Jq5lEsElvHs2OGupu0PCJ300jZj70bqxYTuNmur87pYnDr
DQb5kRuVoUIr3fyc/zdC/FH9pcn5M/bgTrEkxYgfIaQOcZ4T2nX7opbeO5S9LrAFw3H5WrH4JUD+
mCkkTboW9kqfgM1Llszusooz2Ucx+dxgYizydseeuZirkGfWM0T5Zvd1xy9asK+05JcAji+rUHJU
EonYrf7Tmy3iRTa/u3v5QHQjKzQhfG4cR9q6iSuKjX/cZ3AbS4IDEtawivhfswqUB3nYi3yGyoI/
lKak51t1Wq398yHK888c6W0w466xrxomUed4K04s1RKoj50BEaAGsyGothCqO8cfSXV7zusvZdGn
tZSJHY1Aq4c2sux8p7/mTy3hjHwTPRe6RywditqAnFiJps+XtkOVslKeccqt/1P/wTP+KULCyM7O
5xQ7tqBImXyiINrzWwT/H28ZHvJf4vmK58KaULDOeHNbw29Rtvsmmern0TML1tN5D8/lxJo0IyvG
PiRmZ36Ot0HMtriw7gsSGPfOZcgHRC+NJVJfu6UPIWtG9Pz9W6uxGYQZJ1CWl00wVyOdlV1/FBB7
VWhqFHYkQMH38+I3iTdOBi1Oz5s832MxiKhbIOzDLY5R94ChP0h5hMSDspHR6J8X3UIj3WeQhySH
SWurJU5zyPR0Q9B5BATnsfNN2h07UkTjT2XdW9PLrX7w9qBt6iKf0wPW345Lu+b5aqHiu1UsJP6j
dHImKjfsKsT19d88SoY4EJ3br18TIcFngC29AuIg7IKIZrTogIdD35diJYFPzXIUhTDcXudi93ZD
OVsR34JrWqszhUF2arNJ4kBmodfzMVGbToh8PTXfXhSGPp+I7DZ0whvVfpK348U8E/wyPSH5mV2i
RPQR2COFFFtcAHwbOFZiA5jc2O3Wv53B3KwwRyw9097wzbnaZJ1EnCoSlw/iSm8blnby/svksG3g
H1lTFfyykZFDPuJFKVs0GuRidpSWF7WwSSpFCXAgMd0jg4jd9E46OOOQqKT/721prSHrL2Rk9dJq
sDkyTRfOnDAx+sKLuhXx+0dFy1KgBKij/v6aIrD/Mod3nRsSgoIEnuIfVLSD5FTNYOFZLjL7kV+8
MdaG6SliYctoCzz/RXe7AojK1CqUX74wz05GSQltSZ68BmLJhdxy50RddIRGZ7fRKxJ6g4UNNP3z
EEzsvp4nUaZ5FXGu0QRFhuaugSb6l5x8v6mpfU5LAt7a7Jj7ySRkd2AOVws8DDLaQHWJRT6YQ0J4
BHVMX3GZ2AgoLCCqFhAkinl85QzLdn39VjGwa/U08huBkk76+2Vtr09Ju6ypRldJG3QVuud20Knu
lmrr6b8AjVrXeiuUnzwbEs/nxOVdk708jGVubOrIsih53fVkJAUZqOo0ODge38za0NgLGoizohsv
Od9sN3bK3xn39LzSgQy3MMhFZy7iKICXNn90RePFxh8OErotsEXZHLuvvH3VycH69Vk7i4g9vpGn
hHp9KwrCbGlKoStf6lmApBLEcdlhoQq6ur3mZ6Hie/yK/7fy8dvJZs4Uz0hIeT6Ole72bBJqO5t5
XjpPX4SgtVS2neGUJsTsiqPvt8olImPKn1gSSW8Oi4/rq5EpO8l9KEMsR+tT4C/U+GZK0GxJ6/Hk
N0OYABLMHovv6nagypplQgMVJwHbY6mHkDQRwWZ29WKqxHdEKDnDJfmhVYNECmU+h8xDP9bVDPNM
BW7IPwnQIMZrie+bDmC1Tb33syrT8ubMx4VDcjXFuzskX9SUNJQfRfNwVMpN3Hg5zH4Aa03jFK2Q
vyACBZwOewWa0ID/4XPyZiYf3FzTe4DkfD5xMHxkkO3ab8GuyhDIHHXEhHWdnXgQLi9cA5L3XVQg
/LAy5EyRbEKac53zr5cPsB7ir+1KYgIlAN5tXrcIu/dPJTjv/NDz5T6E/mhBdgtW6uM22ChUdSnQ
nHmrFtJ3pCLEhl80qRd6w/VYR7LpjBJI566Q9l1RE/eCeHAYCYqAk+Gu93EXvxM/2pF6PbGZfaxG
Ipibk7f6qfpky/zGqGNaWGBKWfKoDzNTPajNjjQ3908Irg0srTlUBFRzVtofNqCm7Jb7N7U0Pm9w
XR/1v1Bl0iZku3/p6Sblxoi4UlSaXkrqqzk3FhBtcmpfjQEfXVh69YLEtWvl281omVGWumE6NQ0w
gZR3jXwXWfXbucijbPKI831Nmx5J00cvAoNb5UXTt8FUJXiIKm+m21kHBvTxnoGsRq2w0Pjj2Ci9
rN6wQYBRAc8DeGajfS9CIKYGhKV0wwlzocYOFTTSXjdUm/kF3xnPEiAVzGDiGNzKT7xr2oTrRPcV
BvyWOfJh+V6eVMzJymr+scaU6dfaSazpNmrTypBIhQptc5vGUB2C8bjqZ+3Q5tLq6+0lEMij6UUJ
vIjqXdNOCpAy1BiUYjtddp1D0suHmmzIqW6D3CUE9t/X5fKYptYDe4pmSZiwmIE/0Vff8dErJ6mm
iMNR7H/IJXJ0CvCg2WcIvp8qVHoRyQT6oIvaRbnbttmFbROOTC2lQUVeZ2E8F3+9w4lhp7NDsLTa
uzGOdu0+8LUpcRqtfFNZiAskPeLP6lG1CUBX4hC+EKzZi0ESnzVK97P5ScvMKBZO5QGOJlVukGHg
+nL6V+gIp8+vsoxKMVYfBtYIhQlDuFbutEAgcfduQegP1OMVw5ZLXrDEWVNFDWEbZ+8jltX8ZFFb
/sG3cf+9Hd3o8n0A2Jt3/G68yLN2YdhFDT0ckOQ4FdcGnSAFsiK/kfcpLIG6/QPpQbg7wclez3YH
8Db6rz/LrUl7z5angIRqf+WSbTJQQ08lkUstaW4aNTTo45IuGx2qeDd8Bx64esnHFTBLW9+wXRtV
HhiKYqnvVX7f6ZVXgdSVRTwHdMEXohNZjDFAx8k6aR24IhaBO+/i0ATjZxuIHGlIp2sRJps7Hm3s
xRhLvM0dRn+ui+evXarhXCDMNfF9C/NBH71UjqgHEqtvFaJhx0VAQNkuxWNLUqS7UzvjCUDe0Qpy
aweqxlIuVnlz8Qd7FZJKBHgux7VqDDp0c3h4AOl3Q9GzltrHm16zKCUCnYmYnLR/9UUlW526+cDj
Db2SQXJYd8uFm98PRxEdUOI1dNGhZulsYgcVxAvgyRF6GVFmLVedc7ydMpz49b+yBAhwPxMG+rKi
/vNQFBLfgS8IBO+qr9wtO95kA0jiLmCXNa9+PeDneIY7wk6VAVcGSuGE0jk4+/V10gEOofua2oCv
M+1S+KAm0Opfc/Uv8Uq4e1f9hwkgsC62WjbVpaSLp+ayOhBJzpJf0Rcs25JBGPO/Z+jeHHNZiYiH
axIz3o+lEqIc7HBnJihB6OFuhcFode6DJgJJZL5560uKlSuG9Ps+Fpv4yPKpJyReSp7lPkAR0zhJ
l1D5zYrwHf+zz9O9TkZjb3VVt+IM9UZm+aYN53UJmLLiPs8oNQvfWtZTho5rfFtwXfp8NthFr9Yp
CV7zMp5sbelsGGnT2WvzCx8dMykqmPlAMWmLwQjsBy/MBnIcY5SwEEJN0QcsARUIoPwroVxTOdt3
WXShPHC3pnLFGQP3gYq6khuMxom/KXG/pFNeBUpv3AXBeM/MjhCRrNhK5H6g5u72tBktZGcd/1HT
UnsVzVoqr399etD/lr9+y7PL1gAlnqAhrgrqsYkYtVEl2TDXnyf3ljRvPVlBNR9cPvqvyUEbtjfj
3Bv3Z5Gaogqu4G9PilsJMy2keGIwlH+RJ17oo2QnKH+SF6SlDecjlFL26UQYWPxFS6qFMskIG3xz
DVlGPVkYE/CZDpjEybY6U/FgKa+HXtZOb2OXQa3Ln0AHznMlGGagM61FrQ3VrfF00YfVrkz0ICvV
nd82wyWzzy2cccnMmhXumghIBG1FBNvvRdrGYD3acAwxAK4Jv1NawGsnsX4h8jpqFnkIQUGpTnCp
Rrr5aa1BFXsrtBmpySQU4Sj7mrrVaUYjT+b9ZQPb4hAtBLrCGi1IIJJGQUGU3alQozm2p9rze0Zj
U9TfNhukf4Rs8q0hyFWF6ujDQidRxc/9Po9cFeSrB2CxCiyInhJLmpv9dRKRSzKhW498JU1XeAPA
kn6kYSifN6/q6gZjVap9YHJySYAaeF8U3hiQNhj/bJS9g3qniCQVSMwRXP5Q1EOlmuF1g/3BVW5H
DQ65p0TYEmpjdcMEmeqp4UXEC2ou1Do4VS03YqweiLELdr9YZkWTHS7DIWXvY5A9MBMQbOPKehy4
lRUuNpJLdx+vsfJHRL4j6IvH469iPPBYpGoMt6kwucWLka2i2grow8yt9KtnkqoZ+vl3iFeElzU+
zdKyYI0iNgkQ5ECj0RkBsdSiQcYzbIbXQ8S43pEhIzSONkA50pqwXCnken4SrHIl7gNEag7jJooL
xR0SMxQcHM2XMnZA4i1fM1/ELCKSo4kFhrDyuffGDGiUohBUQnpDZCJEietChB4ZSgPAmaLdiMUF
O65+fAbREiYKqS8x/p4QNtuDlL8EuGUFrUoApe9luTZCWZjhdv2OKoMzrANy7xAJVrrs963zR7Y7
Q0GFjWFP/ktX7oGXPVcUaGu4PN9aK5B8c8Q4QMmwA4POBcpDn+iys76axSncnTDWbiEvOw0VD3PG
1ZkIf2I4tCfS/aGc6zUoWnRPPy1iU1uzAF+4sygSIGs8mJVdCyiwEfp+7HzzdGmQ/ZXaLE1t9sJ/
rEqBaNcxdhLlSMOlakct4hYtlakZ4jtYbLG+T8dEtCORTIVmEuiej4PRiUvE/Rahcwbmkiq7+CTx
5buWuQ3HRpXxaixsDuzMX03nhufiTSKEjMDTamoOkJ7qwKgtKd1rZ51boPN2rIfqFwED37G/fUIU
Z7zsbBKn70exCBoVi17QsYFZAzQQA/Dyx9NENafxs7tTSlOdwbY9I/AgVv79737w1ktnkphac4+y
6bzwtjIx/fqsLNUQVeRXNeFx2Z2qsTTqYntuMq5TzY2FyQJOFE0xCL5A/9egNvTGh/q6QCchxRST
1VaehNlMYq797p8DABpGL7kidrsdIRaVFbUua66kaho8jF66VH+XCrwU0TV6KcyL2QMGZVovGLmj
zJbWwrL2PAeEBon6zNgb9D6EdqWG4ruQv9qYbdWtSPBnP36qtPUi+jjDj05ZRLrECYmgSRsq9hcF
RfN7Qpl59kR9RyaBPFfU/JYcVSj7CyLhwA8GCJPHEmS+3YryVoy76ScTxSc+C0AYdF6ZpbWEKsUQ
QC72smSsBbw7wvsV6nZgzm2VYz48TDJMc05m12eosBXRsu5WGNcWmAHgyHKa/J3NMwsMgVmkyxht
ICL+/J7kwkATcUYqI+sWs57d2t+LAniLblwZMrV/tzS85u3OqvBa0A+UNsWp2t77PkbXQic0d51e
ZmyFZdr15OD6GMAbJo1imbuyaP1yfM0AaPrZdQ5RgNUygZznjiJn1KCIo4En8EoFLAIaenZyd7bL
KudDeYam0EKOB81Gz1TDTISVwXJEoahoqhAZYRr8JvzLX2nZ1AFHFXyXafMwAOdI5XmN8SG9rkEv
Lfu36Qs4adP5nIgpxskedukaxvS6jT4LY5RzwLeRFO5hPSqHVF3rdRs6DqqCrKalnBfSxexM8K5u
64UCp0ek/IWZaGTHUGsv6k+av0BI3YgADZBVYzkaOSlJXMN/hhQJD5Yc6LoyHFsGW7WkSm10abzP
rsliN4tk0froEXpXKV+YVO6ThCCl3mHOemvMt2OE/Nx1xwZ8DY2yDzoPQZb6WilgF1Pl3J9AdX7x
+9iqq+EsLU2cKlJmcaZlaFZtCDWaMjXdqkXCQY4FwJ/rtYq9ExrXk5vPQsSPyvipKR43Tw3L1KKr
Jd1ukd3iJy87zxreOsVdyqGWmWGTQMob33CFcjo2U8LQUflpEbkitKurSAgsMdSFy8ZtV5uV59Vl
8AIObCw+yYBEnNP/T9tlGXVJVg5mMjDkBygyEyBXWRts5KsO3qTem9/pEB0IWYb+6M1JEnx68aD3
W+ihpeYtWJ106Y4H0CWP/lbpO0q1pZpBt+386a9nNEXcsogcRfLeATtE0fDOcCfLUGMaoRGPWK9P
hI3PRGbLEkDPu9tfGN76GcW6hmjGkU9DDAWAOH7drPOoJJO7zwBZocEvh8bWJINdAWho5nHF8JMS
Zgrj2rrUlzqeiP6ivUIBUA6VhBHqDgPfcsFsOXdRoEY3ivqpwd9x+5Lf220DB44v/4I3U9Szqd5H
YkAYzgBLXG7ZX8WH6ujcKDe3hLYNM0eVrfIo4E3TykZI4Yk17BHZ6zmy5VRq1d8RWK1SUaHbgN7h
d21fy74+rtgDl3V/jAf1CQZ0H/gUXt5I4JGVYDYC6dTSRx2mVK6OGU+iy2FVKb75+WnB55i1ATsa
21JvY17yAZMPofAaRqp7wjGrtDoSu1vH2fxkB+AMtthfelAbAZWJnawjYFOHAfBZaA6hS7VYIhCw
9I0eaaUbqYnbChkJFPhgJs08dZEo7/5vbKp5/qqZyI1uRmwAwyxvtA6RIYsvOiYPTsf4QgtjLv1b
ALmUM2eLGk4nm/7iiWxdx+n+M7CAv2FjFfA2FqkQwrNogUqSeYepDw63bh5FEYnDXd4daB7KBrEy
/f/XQ2glIRmJ/w9fVeS/jvvua4R8l6CbyNK51pa3+MSEkYQQifyy6BoO3BLzvqAk+OofmtOlx5Z4
Lba4I96iO1VWTCi/jO62axYIsYAVq9p551b8gnbGtUUBz6/R+1h7/i1mnphwWQaBsMn5ITEt7NbT
ZPJ8qScPz3rktZV3b2QCPF81+rJpykHcWuahbV/nQlPt4A0r//Zf+Zht+62bO1JEtV4CkVEDgbJ+
P4UR6OhzTDId8BSmAi3uQHV8SgfwL05sKDWKRz2sK0Czdpt3uvLKbLbPuyHgHP+GwpihGaNvCZAz
Ok2Cl6TOX5Dp/+eUqyd6B2k3fTsk7uPoGGT/kEofU7NQbYzswUVU2xOjOx4NFdx1XFM3MPvTrJi6
RXzcWYb+R21qO2fkt5J7YMrbrOKCIYLu3Jt06sbMWttLUmFjcIab5ApiK5/480yZQJL57UjkbbJf
kAcu00pScsY067X3YO3ro/tg7mhbWjqBRUW72KvOcv5JkjwQyXWDyX0DbdkilPtvckfr5YzxmBZm
dLA8iplZr/PreYzzuQF5YdQsJUS60byjIKDzMIlYNSgUlCRfo0zj5YH+WcrpH58YVubYFN/hib8i
jApGwi9pfn0AuQwfR/YJRY1/a4DdJRfd0d9xz3yYgVrX6HfjKROruqqnJMVpxU5x1gerYErSLevn
NmOJ7b5dkmFX+4u9xh9I04QP55Tzc4/o28d5XRreL6KP7oA1XtbLGpYgmYRPRrR4LB7NfoiAueHC
5DuI9Z38uxw+LZ9bE4ZAU7XkB0lScWdMk6mKCxtdoLQJIcf1V4ASp8uTtjISVfYnjQUhsL/x/W5g
Hq0jJlpPDoM+te4OoBt86xLYhJgUre9W0AKzNx+zwbYtIxMB+O5OMf5r1e0B1SmQ6Gtof+m551Rw
4+IH96KPFDSuDRaxWaCZkVHV+kVshD81YWAVzIv1RACZizCOvM3+wB0MafJuEv/3rhSTm237rnjU
JbZkUsmgu3/xp5QFxKxSULIa132jRwO2BLmbZF1qeBlKnnJklorw8t9KV722efMQtBoO/BpIA0v5
U0lQAsv3gjJzmctb8lImgAthzC7SO7U6chiZc8aR8cSVwjzCDFDUBSazM+WesBCtCkXPSYsZ8y0m
VgzvAgHKFyGMhyXE5ZI48kc+6/c77afpxr7zvVe9epILKSYp0nlhO9fg+i6g7LBPXjwIL2P/i0i/
IofK/sXvDt+NQ9f8UUA9FprKfBfJaskgrcFME1NrdEI2Fh31jpeluBsGAugmEt1PJTdAuE+loi7Q
kGM9W3v/A5v5ko8m2vwAfa4G/Liio37MAOHc4HBpSYt2tR2Nu7BboBeVP86i1rgKWuklq1haXGdo
M0Bga3/cLiesqNA8YE52NWankN+FcOze/1swUdJ07bLIm2mqV28CfEvigtUCJYFLufEzdbXBKHFO
PLHelVcEFHQ45IUl9f6Zf1Sl/LRWcE4DE8mPAjmzsv7cVoUMtdrj+J/yBcbX3n7CYu1o8fTJKr2l
5ZLNhZ83X0pnFS9f4yNVwKt+wPuHoiM+dKAHMcy18EeRgukwuiihaGAErxXEOtn7AvLCLcfCwLjc
J7QdMczDi1mTC/xxtyDyeUWDOTp+9YUgXkA2AdR+Iuu89UuJU9YoCZ0zzzdHTtvYFJr+Uqhr1gTP
gx4YivuGVsSGUKkRXUPVEfiKKwf7YtjbUE1Y3SDJhPAuQJFMZmdc8+TSWd+6P0gw/4GXLX4bO4wG
A24Qys2nweVqzkMvGJwY64vDm7z34C/FGQQZYd57mg1yvLnvJX0r4n58C5KWum+Uxh1AqtnleuNY
lAC+GthEj0Fe3JkVHC7NFnqhdCM3gaiTOv6USXnDoMN8Z4AUPqPkp9dB2sW1NuUp+3oO3W2FybgG
wL/SVoyP4pd+5/yFF0kecigXlFE/4uWXgC/MYKzN7msYeVepD/+/JD6riYXQsbeyB+8FjWcJRGdv
whn0fPDEShCOV0sI1Y0rqf4R6Qd3yHx+w2Q67gGqyfbrTiWi4e6bWBaTHfX8JBMnTMCZmayNnHKr
UMQr5Swa10dhg+RB50ViWEZYtZQC/r2WPMudSOV+lyEU8kj4CZmrB19r93vQa+vdbZ8O9lpWPuXq
oeReH1aREcF4t1cUf5DDxEeAD4JqVeRgVLuxAIl4ILvTz5dgNHGa7z52bfcA6fZ9kyQ1PtSZkmQH
IJPNlTOgUPKh+ngaHnGfbI2kSPXGm2DrxY6nLO8r1HvvHPtavaO1tiTP8houKFzcEEsvInWHRG+H
/f+L17lvL2vt2yamDGzv2GerPLcXAYQVq9DixdL1ft00Jum61DIsK7T+7k37QqL36+I2SAV08ohN
85RfRwidpToiOiCvdiiuNRZ7xp0elnpczCdM+rBlS7DEwBxYZysBLMhPAkr/MeM0Z2sZg3OZy4Ed
o6EPj6fqJe6lC7daQ3PVoEknTgVAeXqWtACoOiP6nm1LwuTEiwazHYnamLUoqNKClDIe9LjzVsxY
vHEvCYv6+eUfKpd5Gvvc5u2EoGoXNpk/K3Z97HWiT2gM/57fSZp9e7+Hw+AbzghOQZmOR+hnhcay
DkoNaV3feLg70/hvIlylPp7G6XGNdAVwEyaiEzybZFJOJT05a640v7gi+Flnr2DGkBz54Zwev5NE
IaRGfPAHxoniTNv8qibHlUWObq1BbdO5FsNJMSBY8d4WbndZBGIW996MVhV5+w7n044dEi5BYm4K
FBcSdmXWnPTyMMd0cnngr1bpiSLxP1KPeCxeURAdRxgeMFPfsCrsfWJn2roJtUywZtxLCkqAu2sH
kqnAiVG34tXUZhqwdAeZfv0mh1H7P+IcGK+OU9DbJ9MlQFpXvxXKHURxKBv8cqubltJH69KaJtLp
W59UpgLjHh3gY96lqzjAu7VmaGons7sozGNcB4sK6aXj4W3klxs3wt0Fj2MksS1VGH8i6oN0l/sl
0vxqtKnPtmi8d3FRva0baEjE9luN/MavXMrFByMGbeSEv1wdSVuJ43UIbmWR7NEVsbYFzY0Juy0x
EsdYM3OGorwZ9L+LkDMkXGDp3J+LPhfrwLyUUislTx3QcO4ufQu6YBax33U1/PjZtOJx7XBeABQR
cDLuRH5YHgPbOU2SheieNYGLJBSLsFk/eI8nYnIm+gto6MllTCC4ElhKym8VEOF0Q/UZLKmPHbuN
jloCRCXIE0tmjLbz1ExuGBOyyadTV9vkJa3CH+XClzaKm5FQ3ywI3ulDE3msqnSPw7d74r/HpEgu
erav+vbr5I+YkS9hVc6tT3o+OP5ps3EUAo68Qa+m7WOnCDffPZktAUTTupMwwhzmrCRmfAXE4KBU
n9N7rNuPUCpKDaNIi9G5zyWbaK1sIraPflDZ1l4R8ud08x7nZs6GV4iEhxAqUNfQBFoCYMfmr2KB
pKqnQqKUFTrG7yi/Ub5w1d6/73YSBQMBEgF9THFbFBsaiLyHyy+VJv5CW2EWokfzKHaBWZXDP3ju
/S7jbSRQvaU0lcgEgMaAV4lRMrX3SuwvWAhd/lp5hWZyW/TdUdcszR7mVIFnSFhI8qqRRWZisxSS
k+FY+4QGlS6wExh5OC6PtYq0SmtSCL5QvXQ18dPJNaPOncAD41+oy1JnJPeVsjXOWQT2t6Hhfg7m
qy4Y0nKUK1QSAnm11UbghdA5JCpHgNdZVgKPxSPNvDjMZymVrbRPRytb7YKlNNiswo8/+ClCpqTC
wjOHHe3WSW1H1b320AWv18NacStODnjcY+Qa83dDrLOWbOQNqNNbEfqSFg9HmG4/l81PXqyoe/k2
HRh6sNZsn/B61mSy7E/Clj/C8SOxvGrdR3nIm/BHDZi9WtP8oAwEig+yUEW9+7OEeN1VaiXZx84a
k0lhB+dsGWAtxyBbzVI+MEf9MdDihCxdnihATQI2vpqIWZw3wO3uX/JB+W7htP/2rjy3Qv7osEM/
qan7oI/7uXVmyeUySXZ93/caOYOzZ0Zfvfwspsk6cCU+rAXR7LnWojuVjF389qkP81yMRbJhIBhU
vDqOVxkxLN2RcG5Hnr0WYwRC32fgzZxY+qd9AkFDajPooLuOKcIBMRSKBsMlbYfR0Kz+RZ428MRC
1cXNQ1cc5dfzhRn38xljjA+lZ5/pD0m/EIHzTDqcm898yB/ssQ3nTmdMbwDZccHNIhM4utJi+hR0
4Nhg3ru+4kDEEdE5hjttIPV0p9sH3zhY8J2re2ZeoxZOKFFwya6Ewtl25RLy15snh0aTWf/iWg2G
FRoY/5A/3vyoOaJ3GTfLZjgX4bY77aFG5NBvIuWp3avuqbZTTU+iBiobCdsltrRoSRYXD8h4xA5D
0MO3/69rKXiQ9qz0tKP9L5Zur3rUp5U46bUbYMF1Y+lJwHRgyzoADFD8flPBCLh1//HqQT0IWBmI
8P9vZkKOApyH3P09urNete9vEZWQKIBv8BAdVEDI9yh2cIQ4OeSIdCvCse9lwMyhwRXfaN9gKH1Z
ir1Osz1IuMmW1vXg8jbLBQzcSAU7D9v/SZAqo80L5kCKQM7FrzVxCCQPZAFWz6ZdwX2sEk51Qktz
HfHH4z0dbYWHUSeWjN8tM0oDAGz78vajLHX2GWcNWxTq/pNqigZkO/agF4uDsB8BiSbrPw/ec0n6
gEnmvgNn87l0Qy9MVV/t7L0/fuimGNBRgvOGgQFzRoP6eTgNqa5YrUrNWCQuNtKShhyFXUKU0Pd9
A/ARjepHwXCEp8HmXqUDNlThI+0bwGo1mQOWAEwfjMoTUfjBsQ695RBqhg2avdEwi6vp1Eje1j4N
neTmpNNrE3xilXQcF/RFyfXPoVnCRUspBxdtgSZ7OJ9HkhEceA9po8gO/dRzGlQIHuxSrVfLi18O
/xnolN3/oeC+xtCu+3EWoZ3waUwF4OwJuB6admjVRdfAloiISIdCpEE8M1gb+5dky0z38Q80Wte9
Orc0XC2NzGk57wusjLru7JOd5owAAdK/EUZzfuxG9ro/+XdRYlkkOR8WllWXM0cT7rzXgBEaDBN2
riKz8BTOhbsHQBh3nIX+zGjX6HCbDsZey8/m4hxI0HACwRqgN5XCjXyGJprL/Pl8xR5vpImpWuIJ
tKH9qRV3KBsouGAqknzeXKPH3NaE0GR5VWkQQWIJcBa0ytH7z18Lc/KlQbkTsI7LKGt62mr0bVTd
MVNxBeIBhz5CfvmdXyB2VA0+EAfpt/kVawyAv8wy/IiSoHRDwiJ/rR/l10vZnsey3DuUVeKHOo0K
bE+FCmZ3bzulhQ2gNun5s/aqTuabKJoVSRZY6YEFtFflFDddW8WX/g1qZLQidEu/PpVy/itB43l7
5eHukHX1sloY3qAjcLzNk3yZMjM1qkvo6MNCNimms+N0ABS5HKHN5+u09KAMdUAQsBV8A9g9sThH
56LYnbdm6KTEJPb+1ItQzCaatnNec94JxuatST/p+lLgeXGIG8IdcJHVsWZyxylBb94kdBH9U8sv
G5DMvd75myq6tm5jpEtp5tNAuZCJM2PgluZrNl47PffKveptxizoDEP9AGSWCHru+jegxTDLm3Rz
g5x+vVspwXyloygWTSQIaVR9GkamrT/gOzdvJokp8v9mnB6iHhdy0SaVFB/MT0qOlZaAqJtnapAd
BmHtLy4EjGzw92E5bBEUiSc3r1hWrJAh3FS28WGcgXDdv+OykxAkYiyyDbArSS/eoDEahP5Tl0a4
o5nnUlFHoG4cG6FelpH0YKaH+kD/XVq9fU2oLsW3I+APQwsWtljeXTYKrGwnhORCsVwWdWwnwYS4
2qJKBhsOXutThFgU1sBBFGZmg3y95a3MYO5aO/wkZimOOywSestueMAJUbcRfExzdO4UBjr2K7kU
XISyJh3ZbtxP7yKtIKdTgyZj9/g1j0p1VY5fcyt4ycbJGvxwaWS1nWV2LOTNUVfBu5REjIZKf2HJ
i8Q8Dy2DFiPN8MapjxGIR8zH7Jl0GEYzfc0pqThKFptjV+y2l3LG980b5LtZ4UCiqXEzl5bei/Id
PRbU1ym9k2kQ/e+1mzD4VrI3UW/j+F294ElbCy06JU4TY1UBJ6AB/FeaW9JIoaKj8ze7VpU86Rfk
yCFPp/aya36z5jVoVbMZai4YJjlJPPwS7QUg8JOuSJABJuvQ67ypeGJeAKRZxNN5JcGb4eRXMjYZ
uxRTrpzBbR/xHQM/n1vw/LTajHLPbZFkzHvBX83SPzDjDqAJI0WpKG5Mvx+Gy8bqOyT17hDv9swn
z71DChekZXAlvjMIR6VMW25Ve7eTjy9ZrgsYnUy1yUeXbCzkWP8fY8QVFY0cbaA4iMUUU9LRART/
0u15OWcmkBOwbxHQhtNroDne8VTka6CVucayyNmvhuadTqrrwAJbIpyYzyfBXaPXxfuKMAFOIdgS
klWq28NmPKHk4WFodYPkFXq01BdxlIE3IMNCej8SipNKfxJ/45Slb6wouV0IY7LZQrbCDFaTwZ8j
v+yGxAlDQ1vPKTKPLcbqmJPHmT0NqLM+iuMPOYqiV4VjKbLmmdVD7EUcw20Xvh3z9cfmFjO1RYu9
MQniu3yAM3xA/xOOJ1rOm9FLaNbTuuNdICUB83UjbSjsdHRpuJS8VRGUbj+pb573Z4IphAsAoW6q
GPl6/0eei9bRMGdcByFIhV6WzJgwd9HaMconGCuPTYmnX0v4XMjj5RMoUeJmEOS16m1He43qSiqm
Dq+YKOj7myGXUoOzj2SD5C3eAYAfYtwL8AQH/y3pILQ/vNimsCWd2NcjKwvjlXalOGdy93S1tJLz
klHG86bf5SG8Ad7IumH1uuiOtE12g/B/GTAfKpRtdy6tAK3FVSLLDXfTyGP8pxBNTEzjIgvdbTQ0
9Wl8no9yX2hrlpTu0Yh0uVBes3THJjQxVMOgSbgwb1QZgkHmoOpvAKErYaJAWqKWNTL+WChoBGUB
6qntAjRyZgC/j+OunYWELiEdgIAoozEPf+olJUeo10nkgZ4VyLN87gkrIq2u5IeBhPSCwQ+fKLBT
W4ht+Ehbv8+6Lyi/zU+XoCHa08HyHwYmOcTtqOpbTQvUMDjeaephKFxdbxmxfQgdCr5PlDeHcM3n
D+pcQHGU2lpY/7e3eXRF+rZjw4xCVT727jpUsKsg1rpStJ8tSkn7d0jLhovyo7Yx6IcICebyB0hC
NABP3NV/VSKSlF9udJfM/BLkSKBUcz67q63KZy7RfP9b9TD3DqmZHPmWKoKyyC+QBR+Xf4z41I9H
QhGiQynz0VvbSlBl09mcLKYrtdowJ2OghQgdRLhUj5fE1W0HcK4n4ybJH1/f2FRH/L7w05APAxOE
gBcg9AUTgOxVxGwpndLAGKqdWN5mD0882/1bIDroGOjm2A2wMoR03jYYk08aBycpbDTpAfq+n3G5
OFWc9dPY+DyeD7btwuzq1j6uzqXMNRZSXgTZlto30IcjyQwgP0LEFu0A1FH+lWRyNsrrx9VU8NaA
jcF0C2b3VJIIowFBah6AM2WlD/05sdIWgETNe4AahnGnZBWVdZ8BsvSDDyEyXKP2r33Mf1FpIrN9
qT+AcXQbm92mvftacfIV7qX1MTSXeCxIZGiJyw93eFGAWXyikXTRlqhanhhqAA6PApxVv+4r+Y0x
OLfdcKPd5z/B8Vt8OECxQ0S3w7NpcOI0i1PZRxku0JSCWxO8I2s+J+vFj9Y20wKa9cToymo8/XJ4
l36qyWagjX6uYSSiENViTbrk5KfVh/aKWPBkNC7ZBvZnwhA0RfbjyF9NgaLgci6T9472YgPYV9IU
uybxI3CR6mhVqDJJXja9JiCEy9TlDpczt0GGlQcAWgpBK2i6S/Xitrp3wSOCsh7bmwtsv2Vw895F
VfboMhyGr/O+NKusotQkJoGSUv4ZzftJPlUXDgPJMDv7fQdfIxiw47toBqEwL9GMaJZsR/bx3TjO
QzGzzgf0XLCHRcXfKvgeWIOfMkgUGORCTAqOod+4j6aip7/MS1AnfICNopVdxp4vd6ZEvNe1feNr
W6Sd/GObvD6/QPDa0t5qf/Zk1rFHvic+YHZctMKWKYh+O04ZspS2ksDf9Gq87GFFAXfCDvSSGYzy
LB7RScNKRQmSRoF+6XdnaF/Lz0lC+RD/RNjQfDKAfCPjiuRwF7bEM72Tal4aLijqOY1/+Hi+8bf7
9WMYJTiQ7X0zYgX6aEs2qPaAsBDbpwPURdesF2JhVT49XoBtN3jXiWn0LEZYr+PXgx81pitDKJa3
8aMGkESfrsQ9HW1+Ny63yank/W/833nvQpBzV48lG4ZwyeZf9edpc2PIbkNswajJYzTlcq7kBrNu
57iQ+yMRpmlETssG9uYhv3wbySQLoksY5AZdpjyhcXUM1/XduyHeC5PkVVidcNbWk3JROgGJHTWc
oc2UOhznaW4wvmmJ0uq4pjtwJaVfOSEQSRyLL+4trC8jSndaUlSvWSWaoaykX8TSjVHxoqsYgEn/
idGMXWb7owKBOB0GUDk/wv+TSSGyTOSF/Hoywoe8Mg78hqEX8wt0EPjRgRvErzqpX2ZgUXtfUfiB
gouvRxFwM2Alw5v5lBvXP+hjim3QZ3zIrCtwk4xrPJWSJSPT3C+gtRaSYua3CgE2ybI1Yl8Vsa9M
l7AOh6hqDPtl/kOFPmXrBRcvf43s5muQPkKxn/6PhKmll+Q6CThhjPQitWjXBEkHxaWUPpJrJ1M2
eyqztGEp7cHMRFPTxkII0ZLno28L+40MAyQJgbGSiaXXzWn6RFElwdKip7PY02gnau7sqDXEFq42
aHyxUBmV9jJT60WADHkKUf5lxBho61imL+PeWyZXulSfLBkc9y4zEJZYv0r1JG5VxLkph7WtPaQO
u0wPzY4qvX6VWTz+S/LCEWmYHFUQEop4xAO7BpaMFV5IzLPrGppdoxWes4OZOqsZqoyZhNn9rSiI
usDZOetMB/7u2FBbV/jfsG+2kr2y423jLynXtOMlzuW+SeagdrvCPstO0E4uyeuMl/ncEeblaQDA
DUsSYfmjriQ67lw2I/IkGF8SWpZG1FRqYHJWrFVRgf9fE/iYwOcSFXtVK3crDZG3UmRu3xWN/l0t
FClGNrt8/fDsR7r4152Z8i/9VzH2601c/ephbJtYm8mfmjTwgL4xOOFSTxD76GaFVIZGWKwYj/65
0/BzW4lz6ncDkhdj+/+/4JZZ5nyNFgkVsGcTcuVLt1JJivYVj0xZRSB0TT/uGS+W03D9MpLgwcY2
wDFSuq5N5fsPa+WRcKcYRiy0r2p6k25v+hWhswHozkHO9fjUkFZHaTKD32LLI9OC+cRW2SaKJKQk
2Nj3U9NS4eFFnVb569vLYeA5eOhVjLi51VOwHVBiBhpc+4ynDYx9qFAx/n/kOt8bGTea9HT0i3X5
v719qGu2P0Q2NE9fhJlKaNboN7pmDaPSPelS8KepFSoD1rzlNzHn20Din4Dx6fQopUmK3NpFEhYd
Dl2jWST3wPVLtzm8Zxm3NirCdvlRwIJDGZBBDCu8b6ynrBN2T8lEdKRe53dHhpHJoGqi/B8bEtIJ
MXsmUSzMCQ/MKb90kRUbt/njZTOhdBaH9p205Qr4YggWkzFTuq9TsXilyMpg+v/eewA0wLeS9na9
xszvbIOjkLTFbxPJ9lS3bNjsCoC2WRj5kDBLJsTvEmE/L5mSV189ojmdWmSA321i69hYytSt3K1B
mMEHNZboFGsc9CPtVj8re62tO0MPzDuQnMaPs+Gxo1tv6kedhuLOP1KADiECyLYTneSQBb9wW7US
FkA91sMke9yhl72TlrqUHttwZqmfd0xzbGuWG4afPFBtWDjUb3EfsXYlX5/plC9zb5XUq0BHHYxf
Vqfi6wHPyfu7cGebxNkZb8q1IQfht2fplY1aQm0o6HPFgmx8DOP7lwXZHK3KV5IrPHhIGmX0I0ci
gxmN1o05ZMOdYoGQHF4XZQGZ82KIeg9b3IZtPl5BffKsyTc3T1TSCoSPrlzcWO6ULOIFHSBXawyw
4+ZgjCumvkgmYzDUIgj6f8ddMpnFoKM3Gtge/h7yGNBaTwdIzHhvy4H4P8zN5iF8W2m6uslAk02v
3QH6qaubyvtsuD8g36ttXf8Amu7f3iH4ozj1HmatxISvlzD3h0Np2DexHFmGurmFaMTDd6keBd2h
yTgMHUD8XCkzyY2BoFO2TY8evOg+v4Xhs9xd9CRVK1r4RctLZ8cxcFaZakvDtJRrdNJVwpn+H3gc
N0QIHYPJbWRoRyoJZ2rgerlCMg+wA2tuqe6jOVkqSoLBr8M3iNadLDLN2pGdyw3XGpN0wu+bYiL5
9+Sl2gc51rRhR9hDOjQ88gC/i5sfp6UNx/ixoKRjGYmIVjcYAVabd84H5AOQv4S2e3o+TFcUhzND
jGFGPrv4ahxI/qB86BIQEVCOOL0BurMWW8FATkBQvkYC7j9Bv/76LgO47fsSSqXVr1ZjK6amuO9N
QdVMhODwgbmMRXfpJvK72j1x3pgpOjX9rGaO5cGYSI1/pnQHJMrFT7FZuc1h6FyLeNLDp/83nniO
xHvauCT+95dwFHjQWJozyNyGESXwNej8yjOEDLZU0GcxDidUfxKeg717pUKP55g3+vFDU/mhNqI+
DU3WbKYSLlGISg5H+IOAdAsAoRvar/QHJ5+Nwhd0AB10614BqwV2X8YYOmOEhe98SFD4B5taPi/N
BeKi1FsyzA1SWS/tZMZSjQdlOM3VlFRNYqmCNsC23SS/xJ++UHVpOFtFl06Si/NlMR7kxipvyAxt
N1d8Xu+pFZQ6nTh8UjiuQOq+inL7kxywZ3+H8q6tBkBPcIcmm2O36iwbrDwYoZwYxVTmnvnYU2J7
qMtB+2hD+JsbBmgI04j8loLFtc4QD8/ajgNhznOBB9uh0UStSVh/cS+p5a46hJmvyREs1DDo06zc
ta89EL3o6xnsxpx5PLs4OsIfefOqbQkfoFLoJqSr+oPwPagld7cxX2O3c6a1QYwg7AkSpEtH9zJU
uxQ9815usrIxY1FTBT/B/IiBXQ7A+xpOaU4AET+/U/+czRNg61M4kUugCX1NrjTEyt14mujlVK5Q
karWifmtnqNwZEQbUgJKvMLRyGdHtSm44Aj/11H2Qd+OcunEWrMANtf/648tEkmOid2OPg6yBo+S
p+7HIKdY8AveNR3k5dH84EMXWw1qJE/Dq1va/PJnSOLg8oNptQYl4ovn5B9C7sRv8zqG/iqYa+t+
TofEj6Z6Kkp6jGw4s4hODdoeMYU2STit2V3Avgd4Jew47r+gccx79M8P9ZUeuf8yexsouo1KZd6B
agUOX0F++MH7SCIDbgxBExU+PLHyXnY9qEIceA3oZYQr4kB3Mh/kMI/zZJ7bQaHEPGEQYvA9nbHa
mke+pIbyVrBbJP1DvVeq/h5/bT5RhgAfmR2bWFhereTL20hNKef8bzqTfkx4cUEuVPxyySUHqK/S
4tWACxM+1SRPyZLRmP7HvbIqlKsHbn5ZxeL7SwHGK+HOVosP4BePv1XWDv8dD/91ExLzxn2ySwvp
FD3+rE55DMO7ZybA5+AUIrPVA7RhPGKS/qBfyARU4TPWMSj9501Ww/vRI2aX4oCFT3FCFdVb0/BW
+077kL89Cqo9lB+rYCm3417TRJR2G60OnQW4aRXbrqt81prQ/9JXM9P0bhV8YAA90vFdnh8wAq3a
lzfeyNSZs3Zk92N+b4fjLnLGrGpmg9KvWDKSHCF5rUwIq8fEs2q+oCtjXyDSUEt+jYGmpVypGlhO
bFwbGWDmlAqMsj+4Cz8vR/6cKGwTNN//8UQNNSQCnvkPFOz6rncPKhBajUpZKo7O6ecpvOdTYfFo
dHSAQySTEmZAikHhsIpSM3BOiyHQ/27AmzB30SVY8LR8zWhfbIcDjRm2fbmbFyxa8Ktk+FmNktAX
rK1GlC/zLlHcfHy7bbAVOgJClqa5jTDC1cZlIZ/BUaSqDGB3+wi92T6WufmWc3EkVAX0kdbEf1yA
QkCktEH/vgPOGFDcBzCNs8BUDlNml7zkTC7vORUTyYP9SLiQZ9NXorVFVt1g3Y7YRUL/PC/4HmX0
lu0Avf1AS2JROvYMfN/Bn4SUxX3u6+EQ79ad1wo/zdFv35YXqLUH02dO3I9CiSr8B8iWAeRwIjhD
1T5YZ9TIWz1rbOjWsDoSRQXcnfKY9nm3Y0g/Of/gkR/c4+ae8IZhF5X9jXxk0gPk2k0caunUCpNa
VsIfZwFdINeTHj3RhUvWiPIaEN0SwMu+LCuv5PqwtNqVVisgYIbKDZCtxVNqK1xRBlFiEyK2P5L1
+SOB+oD8Lv2ZYqji1txGxPftSbVCmmSPjV9CDaHUjRjOCPoXOGg8DlAvasVqe/PVqJgQNEvL9uBx
iN3bJrJLuq20+8oVbcy0Ed9hR2NqdhHZEopn+P9SqdXdF08syTxNI1Ls+EoJ2eeUgxhev5cqxDUS
HRzgNMDcsCMWPbXylr0HqDBqwK9CxoxlP+MVjZgNurwIQBVGqze8BahZIVwitDpYBHZO1gfVLSZ5
hH2LNKV0wkfNyrJx4QgVvXm8TMi3xKy5j+1PGHG5ZNexNQJ+41eq0ZWS/hbRAmGbg5w7KuqKR1sw
S6sYw/KUUsIf19ECyPW7ap6bh/qKRUYZkkEnPxfPIWQMbLRtgcYcZh/n2GusjN8mbrfym2bcdv2o
QZtv/S4mPRChGyvuODIjI/Jncy0ttBUmZ1i+DzJHIB4qqUuZS+CY/t88IBXaUEQ2lrvAvS12wwDZ
YmBVa2fwMMgKf5ilIaTaqryWmErou7qEUcNyr0GiyCNycNknvHEWbyN2TvxK52rsj7qeXqVep17Q
pZZYF3osmkBurGkALjT4Hcv3levteQd3j04qdTLvHi9/Ko5/K5zYC2hz5nSSw1Abw9I/j4qLysSj
L14KUDStWft5j+/PIQsBLBbiBcYceJabi2k8eTbFufV0MXFmsNDW6wDQIeM1lxzMVp3/qVBzqpj3
lLnAlmawR832ZYa/lA+IoZP9/QEDqrcrEy7t4BhHiN4Fnh0bWo/qyWD3jxJovI9tynnZcM8JudMT
CcDgMMrlGcfOlwrsOqXgkKJZUrBsfsNOMnv7W5USMYD+wYqgc26fkqQEfatkplUPugJ9cASudavY
V2x+wb4gZg0v1bA8RVH7b8br6Cj1TfhmyGLHSwJ034JujWNn53CECrqTuYaelvMM0GZmVb+gUvEz
296qLVJVQN0DFNuLC77JwM85BHpsPhekbC+MqvVI48bkN4FUoxPYBZPC8UOyF6vkYvnWhdGM5xFw
R+93LKmx5WBUgvCcpzkv7PyU7D8waTlFKrktn+myCC6ltVCJmbe1tvLeSQOs+lV0xy6VT9edG0Ks
xGZGeNizv70cfKzokgEHLToeuEwQFD5Nbo8eRFzFVa+TWPOLFI3KCt1ikXH4jKRTCXlfZ7vFTA0Q
voVW/G2j6/haIH6cDHAFs19IDuPUQ3zZ83Q1DQOT04vKaCGaaKI3GGJ7IFtxFyctSty0caJyHCAj
4PFMw/yj8fE1gOciYVIZ2NPMb+LAfhF/NxbPUaYAYr5VI7fSDclmEi8EMlaggMA5hfTxGwDPhoqn
nW0xdTnVLzkuZdQV5EwMJ+H4hehFXfX12DQlWBt3GpHwP1y6Um9DsCPrKx3tbU26rsnic32abRgg
+w4pmhpRRVGpoHzB7oZCj9EzA0LwSuf5LmhIAB9WTNojapnZRZj72rgjW2z2a33eL5Ty+q4E0NCd
uezs43xl35MCJZgTf4/cmQqHlFgihDEuDjpzmJ2FdJPBQkf94AZNbJrcVfkrV/gS5UyklazOnp6f
Frcao4dYcPiCY1CnQxghKt0Otgpwv70+1CBcY71T2xCwNP0Ltf8M8DISl8L+jE0TM5f6+sydcy7k
tEN6SHOFuPoMfj1kc3QGbR1li3mmITo/YK5QgRDhbLeGwfg2Eq9MzfGdp3rqtwG8eiTGaCDmbqZ/
kBCATJ1d5x7UH2XjLtufnnRlxL+9hD+2HyzMEJUJCdJxn8ELoY680+T2pBH6qDUoCJrseM4XQs9v
ylMHMAhjLg9IzvK/2GG4uxZTn1Det2PFbp7nXdFOnYpSzxLvlSDTsvUvcXvSl0czsPSbzZG3ClO9
HnoDpa1KVBr6K7zxYUimzZx0kemmlta7ClBKDeLZZ3myWqtLFybEq4Qf7gHWXWu63aaI0eh6iopa
kUKfFD7yNYQ5fby9x9kexGvFu0EQVv1jFsRbFLFs/ggDxFhIV46KuWND8m7iS6YSPYp2ZjlVWfFh
LIfBZJ4MjPDYr7ZeqX87zVk0c0+VKiGYUY0mJCx4cg8KJxW7rwnBxihjWsLIPisj6ReqGArr/Z0W
cisCrW9zGgvCmOASvgik8/eKB4T3DcG4zmIEPz0ngebPS1xOQAkR+43PlGwwBQc51jt9IdeOKRQa
iUbl0vaHB1uOjMCWIbkz3ZZcZqT/YcWt2h2ZlsfGpdhHeVuMlTslPy3C3anIVOqHxsQTIHSyF2/f
YcAwrUBfsTR6DR5LIcGlVaGM/ePJple2RD0gS7ms/Gh/tQHHu0W+3rJ+LLXMuYFPBrh7g0gBNKWJ
UR+JoLyqkehHwTUqVVeORhQYKEv7gcVXYYfhxOx7LGrurp6x/0Zj7Kd3LPUWkOxC3QT6KSVoVNzT
VEWH+Tdgfm1xj6/+2GR97oxJBMvm4iQmeytrhn5RMee5mNAYy3GB33EFavsoAvwjdkFrcMQt8xp3
036PRuPzi0kU19CKUasOJGVoW57qIxAGmE6d5ycgBdllHoVrc0Xi7ldVoAb3FzPEGmiJuKkHppXu
mGsX/KDBhXqdUcY/5shJqZrrK8Q+ZMYrayI=
`protect end_protected

