

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZqI7Lq/aGyAcoaejBEIk07VX9jYIkvdeTPQu9dSbDEADopcPNa+0k8THWemULZmXocovtHBV2sQ+
UG9Mr3L0hg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
R4vPs+jPUBq40hDi8U6b9avbUk2Eb50U4A+mDDli/Y0olyqpMjS2bHK8VDjTVAFuQ+H3qih0cQYm
+ik1m47VLNMfNDfRLbftE2okRK8Kx81MRcEafr+7z29VxyL2KSwmOKbcDCEkIT1VX5y+96x7q9/g
O5zX1cVuj6hrFncQjBI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RHGRLed4zRtfx3HaMZFysMR3Ua1JohlSUQn/uIq0QNaCK2P96ztDgqQoqe6ZQ11betfsHTRFzq/1
66ClFz6QxXME/fh2KrrXSgUZxYxwfstEZlyOThrSfu+qzCsdk0R654q7wyvVT8+Lni3RuXc5nFXx
raCVZl6qLm50r3EadUq562wDBW7iVkrMp3OgccKyJyw39sT1Jc+0IkzHuHqjKA44tfGTOOSTHNUj
YgsyeZCJS72pabS90ZfprHyjsELB7Bxw/M9/XLEV7l1LP+SCDJFvOP5dNLZDBmwYIJ5OoU7247Tk
wYu3m6ZFZNnTwWGI9SAZJyiXILRa8hVZPL9TSA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OU7rNiePgxinwm/ruLBNeniAmTTLdwPhOZ1i35IGtDWXtaPoMnsPLRF6vnJo1xeYUES1MIlBqaG4
FUeyfrnBl3ofk5rfTbxL16dBcEtA8Z/duJARcLCIBD/J+xf2VlSqIo8dG9Ww8/L9pBTHpNAObSOU
o17xArTTrLfHWXZRGfRwuRpGlTLTYOMvS1AGhQcPbXjHrlijOoz3XigDVsnyGbHfkSgOlGBCnyDS
TPebi8IC8YIl88ieW+lqTL6jl+3DZ55iTfCJKbFt/HrE1Uou1l+60xI/9h9XhrNzE5ANic5eFmyC
tdncsHEBtx+UfZhyFrHV8z72yZoLCX2rOJ+IJA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GUoHfgebfwQKNkw122kR1rRfB4ZFf7/0xjFIvV3auOQ9RcZO2jgecvvtUAn3nocoMNPW1jFFZW0u
xgkVDSrwVJrMR/obpu7gqo1n1FD2E5BpOJV2Gwso9aZGhgTdfd0mINfCxPi4lxUYuTw1vd+iNkBH
peC7j2xzDHSu6o2S58c=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lW3oa+bS7VSdBch0q4Lk4kIel2MxeXNlqo+JkBKYCThE5vtBv3Mob32tRj6s2h8BAos9XGsKRu0r
zWpu3cgAnv8lYIL4/UPBP9T+caGqWHHoGULrLn4zuybUvPzfGPj+ANXGfPXBomTO48UgPFWBnBA2
3vlOjCiOyKLMQAUrg8RqpfdYfcnwHxk8ebrE+lZJf6NCQtrqGu/EnH7PYFH/8MSQa6yey02fLQ2J
HenzdGNam7fu3z20gETHgePuewowRrJu5bEZOzlor2RrSnb0hcSbcO4/KSA9EcbmjzBMjE5uRYAM
1y+0t4rNGr+0XAjpp8m6B8lGF+m1jIGYMJ55eQ==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AYjoOGO5c2rCxRUY5RbgjfKwpMKJQrCDGPu9wzqv2ZhoT9Trod7xJlCnzNNU4kNJPTgmDf05Bkoo
EvR1hgWeTmTgCGdy7Qci0Z0L3pdxnOg9i69qsJO1qAW46sOYPeZHpvATo3irsreTIyOEcblYRdLh
Raj2T02eEhljrx1UdWXHwIq6kJGwbPaiMRXRJewJ75w53lF3nNUwTYgttUbm/hKuK4MTBvyDWlHF
UReBw5kEbERTaRF91+HNJUeoBgfLIgVhtPzX3Yzqy4fl1PxZ0BzAGNRQWfLI4TBSyl64znmxdzaS
+wcpSJ3OHZL4sBSIwGqpZ8UuNr53DWWwkd5lqw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_11", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
F93W5rP9wRsskpVAtvm9VhlFJY5TOuivcFKT2bVYmeqxn925TMU0N0nDRJZmC+O7NbtC0kbL9Hfv
iPaQAjkvtWKCEafU216A83pjNwYVINq3GbStXAtCrvf3KbYJMQPnr6FzKWLa0RlmEqf2z1LRIJMY
cR3LKzziLGgP+oQLz6W3siXeoyqxsbDm+dasSbu2YxzGAvkTos4kX2slGrQzxYSQogS6j/MzVgIk
Vhsm3BYDbtVT5TsiHGfRfi137tS2Q9o11KN44GT+JYigwORe+GyKi5xjI6kGPl1N1DK12TlRGsgC
Wq2YWMn2ABYXE2F8mkwPOJqSaaAR0S5MMCjkaQ==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EO2KlFB8vWgjeXvua8SEZL2APl0WfdPtqoF/0VTjBDZhkKh8T7GBS9tSSrCin7kHRBUGF6hOUPK2
V0JQtp4yW7c3oVbMN2ePIV7UdtkAszA2lMqOqeKJbWn0TfxRWL5adG+jGlhhYEbaT6tkCGPbbtbk
y5Kew5kT3RyGP8Rb0tim3cGvqi2BdBxqdc5Sb+Vyj0havZUyZo1AsjuLnNukDIYIrPCtqOY22MTp
VlNOr/u23OIMx+xx7Z4aOvZacPCxfg662ljyHetf5a0wu31WI6zf/69lkXq1iWJtHgEJn2iDpIWs
bSWDEtGgKAFHGKVAoc0vIGP3aPG6DIsqRyQ90Q==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967968)
`protect data_block
g+/zY5eCfOcGMzGb96U+wytPoD4CHZv/+wp2Ig3baN9soImfBUchpOff9xtgmXnr2u9wbjNkZmCG
11rLIPpM6U947MQDthHIljMQRJc9NuIUjcxiBR7o0yDOBzVY6tVShKrQWe5SAQAPxZbbL4BeBCm8
7XjIDyhjLkE60haG16X3rN4HWSpqB6iLHCGQSAnO5Kpo5htnVArqiml6nnhRJiMik36YlNz89Hwm
Lk1ssCRJ170w+XooIUzgV8AWYlfpVgeqKU9Un/RHlce1t3K9C1UXSU8abqYJxOXcOzZno2wo/sPI
0uIJf85n2K2qrMxGfNmxbhA6xHOJsWhTG1aPAgISW1XYqWMRFNAteKMarVyNQHcrtsbrK/2AMpc9
Rs6PtsDqAb8D5s2jr/AwUFgosycdJ6FB71vcMxlVUgOdcuU6s8qRBSYnWrhQKivjRBPyCEh+FvzY
Cc6kcovEUiU7cFQ998udFbrIiZoihYZbTLlp9Ql9taUzblYcAuEbOqcpg91fRMn4rmdQUUhUUJM1
y39bNoXZk2y1dAw9e2kQ343/1GVvR+N6tmT7ckcBW8ONmChpvt/qGrP3A12p82HfgTEm3vfv0Ovz
aIp7lufCdddULEolyajvtgF886lFJl9L0bUYoST1mQ1v4xXF/0lTNV6hUdPJCV+ASGe1roTybChG
9nW6977nBDF+/iip5O7Es/e7FSEDRylvwN0Mxw77DX+xMBJQZ3bUqwGcu4rSlUPZLonoKvwQ+yUu
FpHpuL5BGV7Joz4X1V+vm7RH+XLdBjj8IcVx30wgyXGjw+yxKqz468rRE72ot0fhJ8kkMqsaGhPy
/OrOzRTIXU0GuA5lVSt/XZ9M4HQ21qZc2PmmFR4CHKaT2zwnu42U/XXGrekXDHi1Prn+EcqN503+
K2ynN7mcZvesyzwL2XiF6lcvcHvCcZZgXsmrVuk/faLQt+NHqo7orUuDEaKcWcsHDYJi/34PKfPg
/Ad0Dd94yZhMW02SI1ks0bpCyzsbUsQ2il+9oHHIzBZvl0oqExxQfrdH9RuTqXKVY1TNN8h7QGP6
JymyR010CAqUyIR+dTJ8olkmLZ6GyAJ40He8hezsOigP0Kf/gSw+hzDxoC4so459PIpvfPvpy0B5
R3QZJqOWhpoQjuKSYLZZVEh70x6ZZLY9kGfvzClX2GadbO/Pb6dkEI0E0XGWaZZqgPcKOrhotLBK
2DJx3JY5nxLv6YO+sMJTIkYM+Ly0BOUcxakRRxW5DS1ElHoRCu36BX3LvABk4WlLrPkPju3XfXU7
6yN4+XkiO6ixA3fzJ/R2axt84O/KOzm5Anp78Tf5JokL5qe/fANquWW4g3/1Bi0lk5WZT0JL7yrb
agLaqvGr1RKM9TyFoB34Fv8DBTFJP056pbCOqYBjru1lJgwvtNhT5xYca6G7WoSyAN15/QRMOLCj
feig+wBhu8lHVF8iqa2uZRShihkRUJeBK8YiDFBM6Aqu8I94L+fqJB+sH4PxOPzsaJK4fBpoxmwe
OiUrLKbggCmsPs3fl2yqFbOXX0+sudOSojfBp+cBt37nLPT8wntO/ZLN5MymWmYgNTV1QUr4vEyO
g8bd52QwR4HPp4YieZtbVX+li9v/pLHtEUWzctcbslJEKoafO4A6drDZZP51ETFYHq0s9Ifw8Drr
MaNM5RqyUbZ77taNE0a64hjOkzn2XSCBxhzd7Hxkcv3pPgQHXkyYZHfSaz+FZYo66TYKO5VSc6Ix
ts7+l2pdQW64m8sMoYtRqpYtO6Q4kfQuFhjXtlkGBHNFjwd7TLEGaoWE5wnIP707/ANwN4cIwGPP
KkDsYXh2IADh3mCHT2M+hhhcXr7PxX+8A5LGYHtfh28mX3Ym0qayxWaOz3nuKXqd8tGFGEqnmAMc
QXGk8XC/S5uhOAS6w5WL5G76Hfsz0kB8o8LzasAsB6/LCVuR39TF5G9f5GAJ16pm67kGA7Yy96r/
M5JCDDMSHO2VGonYMTgdamOt0vTTxIJiKY5bohH3VX6MsHwCX+3IMxiPc4RBZzUw6rStOYBTKmKF
wM0vYS/SHTYJmrQy0yDA/dRYpTroc6/aQT7X8x7k2LeKPB8IQ0SYDyDPZ48DPBjryoYHbFusHovg
ff3AnPBrMaFzzHFG8dfJfr0tIM6jSEUXhk+SFXYAKnnAmkWJCHneYTZgBPjEuYgfWh1tOIql25Qg
/J5BSnBeDKUIBmNMCldCJILAKSRBr0Qj9Ohzd+P+h1giaygULwjJow2iLBwrZcbNmmGa1S69zB5A
ScKZfQRVrnDMgYevyOKE0oSgUkz+Q36/8ysCJuG4RlZVu7yDO8ZBVTidTYcDVja25HUE/34Eu9zV
B65z2i74c8lknwq4xMiUaVgG4IDNXBxy+BaRL0bLl+CzPYQKt7gShenB3hV00/cM+ovZSzB+qb6E
V+kw7xYhqoR4Opl2vmEB96oAf7lqxbuKbNfFLhRAP5s+qShJ3WOsUOxymCw35wME9xqChDCUJC1m
BQc20VgAuJjDRtg3QMWOFMiOZ6BDT5VrlDEbJ0bs9AAaLnUmp1km5GTfbXhIHqr5zs5IZr0l5pYg
eBb5lCn0IeytZymApjY1ZivM5qnE4qNQz8AJRtYCNgTsOuFAHq6CCajKwfeWn4njcvoqjNqtRWZQ
xKk2GxZSpJoIVEsLm5ZHPp1H/LAfOtKoXwLMTG0cUEMf/kAvhiGvRCOoqt+8aSwx+MS7GzY6X9bN
ym5kydobp75F/jHy4SKw5RC61EHyymzac7TYawyA0aCVgCbciYrEFnFZNir/qRRfQqQa/571x3GJ
J4UGFkMwSL6oonoRU4OEMPYGXa9rccwi3lAITtBG/HUN3JpVdujn2vUxY3zDlfBRVDEgpcRb/fiR
uPvV5jQtfUaFQcVRSi1afOfpKZzHqPe/NOZW0az7ZtrEMHM2xnNxpbddDGKFRdFyXKOv2Qw1LQXJ
eU7XgcK+k14zOVEF4zEDWBEpUcg4D2zTHFhq1smZyW3x8cHVog3af0/naKjl6NYNId/Utrw4MYdh
boefRpUL2siy6oL7YuCAi/VAMI+YJcyxS4p2ldWhQ/JtzA9mc45VEr2BU+7CmcHgnMSRXulu4ofQ
LDvgyOBfNk2GXX92OYCzDBzKrBGKEVcQn6Sn89gug7z2LbnKVoqS5mV5uYVV9ygdsf7fWoj7RpNR
XuTVnyNn6rUbu+A9ZEeQQQeGgPcaYzYXjQZ+wUEVIZBg4CVDrxhUkRbpHVBuho8o3HCwrB/MBwb2
t1FjmG6R/dnDUURa0m9a8K9wJD897NhqXwnE0TukqSANnBP6cx/XCVTT1UMygWj0TBFVAImDE9WS
z3zN8zZaeScrzyzItSx8jBDvtBkfo1vzt1JLR081xElbYoHPG5bcYcjpPnXKXWl4V3VAWAN/4/5o
Ub78vQGm9JJ2e6YWLGDPcCu4FO1FS+YvvuSGhqV4DMd3BuEr6kSGwwXTecAqauQGY2p8S7BVnwCW
bCaDV95LiesCT+gfbzOp5LD2Qj8JtYYGLNxXjSUr6QMo4ZaYFIBFXKyXoYcxX9ZyLhRJVAeVLCMA
96kxkghpi3IzIi7fV3n0rzMfPZpDsWhGLz47ZVpG//vyqbCkPzUVZL0WO3cM/UTnhkxh1N/WT6yI
JgPGvGU/YQurcRkp5U6cfnn6Odxe8H93hr0ki2WIZkRu48jSrCLVukcUceazTO9A/zPW78pmtnVL
QchGSg/jZ7eGFZxPoOD7ijE4xKwGGOMgVDoiyNljFKSsAyi3kQ99O3spzHJz9o9LCkWyT71aCg4L
vEw1ZJ9w/dArI9+VONTxcb6cHcBFZYGNXVosHAyvXFmaI7M1pkNYHv2lsqgTSPF7n64GHtsF3Os1
34S4Thjak7C3Fabtije6CaPno7QsJl4VqOw+51e0QVGzIqloVJ0m6Di8itqA5XXr6b0KDXAn6mie
xrPyFq0V4f3ot7XptFrngYNcu7fynWolQy3AJJb8YWACWBVsWglQRystdjnq2DFutCVs3TUu2zXv
iohvzXF9zpRQUoWibodnHVwn8V0Oyg2JIOIpadXtNa+yhWHP0CJugGTzZc4KpsLE9N57dGxKhApI
KmifiE9+WGaKLDQv62uZFg8qZnXkNSo0TUBUetnz8imtK4WW3gP0c4BtsDK3uNAJxH7VtFPqnetO
Fx/qImOwVQoRQqmSasdNaigO8H06ZPP8AOND01mRd9iTFETcewxm1P8GbYixuedyJ0G2hiv7pZFx
0WRuOotcmJaNJz6E7P9MxyiQt+wW/53KJdiJpCh6cr4JiCxutQ9NNYdV5NAOGnAGmYqmh8nGCDyq
bASbuAUc4F/DsMpnalxvAzQ/U/GoTKoF/gcvo4p2UJIZbf/x2MIfmgKobOsYPxPCe5r9Ccm/cCkX
9AOm112RmmVrRF47FeCIMaQ1RWYkSRBuRHEBACk/Hni2d6GaLBeS2xTXwOboxhcsaHGqBaytVy4g
dgaWS2BijsiyH7fxeXZQNg3z3WE3FMYYfvzqP3JuzpmrfrBxUanV45G3DDj+m5O7bpjb6zQi1IAo
MF0LFBaLgOOG4AL8J52LE5F++xSTxSUF55odGq6LadAzJsu1QuVi8W3S6sB5PC7Eq7SNeboKwMQU
DFBvI4eTkT9k/bsnxkw352oYxEjC2N7qo1N+m+pd86laJfnOGcjAgmnC4i67xGHN3ZqbOl5HU41X
P5YlnW/1oMVoes9kYvK5bG8ZfbABIkN11Nz+JUe0POQFUpY0t5pBJP4viM+LVpLtLgKSdBGVDfi8
QjOIVp6dQrlBSJNXUwwhTFZ8QxQUOcP7T01JKNiEUf4Qhszp1i/LC4jX/3VBtpQdDE6Bnp0USpmm
3wFnbR5ndw05/V7U/uL+LpMVUb+0ILPGv/KzfOCZ9auMBch07nUhALUAU/DuJgZ6owC5Di9XZ1Zc
EZTwbzfIEzxSbYRNlBf8YBjS7GqbGhoHQ9jKpW6bavrmn3HDl3davCwjmKaeVb4LdBH4yOjNnoOR
TMFqR232Ua9S/faui0IgPEJSFF5HD5Wq5mGHw+qd5GnSsFlAFZFtAo543bAq2wz2PgNnm1apZqW4
MlB/6Udgo1RvTI4RCULgBmqWs7yp2XwHoNEviFTSi6hjC4y9QSBuaBydGR3qCeJDSauJmgvz1ERh
OhvSzsO8gDZEk8cFY7KqbQRlDk624X+uZS8w0Tn0d4QcId/uLVL1kr1AzCwREsOb8Operf7bC09/
dLJtsKPMtac9YSGv1DDo0tPaogxnzfnxcqic5vVGNXXqy3VIA7/SA0MCGzx1u4Va9MIgH23yHDtt
8DezqyXqUB/YtZxgswuUkrswx4nN9vw87e5a0s/H17RWcChwvqk1yEgtmErdr1+zsKZm19Ji88td
9Ry1MSRDj/uhg6ytP3IRTIUb3yVCHWx3dOvDp8n7rjMcoq9QfnfwWv7Ree8P0qdmxgvvfXxOyFhb
D/krB0fzQuN4gHDPw36CfgBVnN+AhOCFIyCkkSzhFNzfCzTkOWjva4VTYB3k1oSjsqwGeIqfT4B5
mHwhDPrEnCrU40vX1pnqrBf2qMNhSvEcTOVHg3U0m+pqF/pTimYSuznGGynbMcfi3Cf6q2HwABOz
mt8IH8FJFp/jJyOHgvYu4ix6u2YymjBqSUSmVzSG3hxu62qx25ML6dolJSzaTx9Dnb3bP7L+gk8t
F/UoP3imGqA3rj59a5DvV45W/gO2J+fNG9aN6neGuS7NfltrRXvF4ilXihOVcPckbdS4jkQ9A6AB
moLLql9pD+6na2f+c1wzyAJi6VTqFxAOlUlpwMWNVvmZggmD7vAwp6XoPI3mn/eEOmrZqEkds5cu
3Pc2I8mqQFwcDkqkKKhTKS9F5rfELR2CVlVvVTJ19w0FpJm0u84zvAJd/dioZJ80ECnoCKCLVDOU
yUEUzF0MMk06WHgunX92BD19vri9YiQ2OB+Uljl9Yu5PPHov8U82i7jj5TpnyU+/uOFkz6eZ845b
TEq1f4xYxG9xl1uq+iLmnhyq6/YWockyTzje3WaueUQLfz3srYoXMpKeA3/niqhxbjyaYQzPVxDd
Mk5/DHjY7UqwAOe8+z687Rejog+tgS5Xg+nhPF7M7Y3eBlLsN5Cf6rDYoauILbfuls2PmN3SjWZW
vJiJ2+0vzuNLX1e2sVT9ocQ9X4jHAYR61eitHrO4prZRcXxysqbx2NRogDyNYollTBSyxeB/eHLL
WpNDcTx6+gRBgnbSx7A/6TghgF2DpcJ+bgVySPKKVTGn2Q1xsbuK7oFHBeXGeXRbNfRNvp7OicIG
Uq4vV5oUh0JfZwcA41uyaqYnrO/XNU7pwr+oRQquFAhMXIyLzVOFnOtMrjizsL/jjOKW1+Bpk2fQ
R2NAT1LUF81bZCqLMH3afX9DkFlyM82nT+nsl+FXJP0vAfQb7ZdW81tWqwBD6hQWE5RW9cAQaG9x
+n7+uZ5sMcJBZmR+fCEJ7q4ms2Lm+MVp7PZBoTnVPqlfVMK62n+jJoXFgrsAgIpiZj7J4wjd/8Hg
Y4XWCtEnHQIlevgLCNjp2gLdsqR4gHP15LeyqQqjEZILERb+IdULDHZA+yuNfszYKVh4X1e935a8
ZtVFynr1gcZapsV08b0obzyLPIg3TfsB6LB/V67sXR+Zsnwe5+xUXNKldeeQIgq8m/sUv5H5auTR
KiZIHlQTkztY7Dzhh7gexlU37gy/LArDM6+U3Vykg9V02uJQ8tAjIWmyzYLw8nskEosA9VLEqWzC
G/AyXBS9/J5kHP22nAhz13CaSdlEEASi10g0RavALuszJ5yxQru0Z5ozWYPtlFKKDIjgHkxjWNsN
hOW/iBGnhmCXmwEgB3aOE7wh/sW9Gze27l9SnlbdDs8tAmQnBZ6Jgpo/O39u3xRXNVELm9bzREFS
1N7WJy0qq9KHj6iYH3o/oGMeXKSvyNgOpNSgVnI3DZkeKvwiONgqUDLkLcxPl0/8EW0MGo6ZdWa/
PCgrqHaDQNmhrZJaBtANxTxnrqtkT7NVGTZNdnz2V/4IvpRqBxHWElQVKXvV7lUp06KaEiTTTUni
WrS33Vr2ogGjqk4zZ9EV7YPdhk7LtWS03E647Gfvys/xcXei02C2Y9o321hxAKFo8IgsRr0oug82
EH5f3dKDP9u/nfA+LZzDvGoprV2SHwl/TfFuYjMbQ9nxTtyUAXyekTcIdbUWa3Z797D4lbwdtsrP
cTLS1aKeG0mA3J5/QPjq8x6YpP8HpnbpmVGURSfVjMTHXcnXu/3ZFC6KDbBNpSr0O/YA3jxqXdXF
BMTTYI2y9vfp6Kj7X7fQdf7CFqYSS1q0QeuyHrNHK1Tizl9LuLDH0OH55fHhC/pHkA93d2dvK+fT
G+UI9VZl9YoxLUY77F3ikmdgKWm0t/OnbLSguLsjsVTjCoPmrNozmi0cHU/PYtA+GwsUX+f5M0F1
vmDyjT9rBcohjhNaUn54DahDlueahYV1o0iupOiesJskIoVBn6EDuJK5znSswikiH0/vOm2iptaC
oapkR4liJKmg2rR5sIwVceb7RmLoFgSA171+N6KD1brq38L0K3xxlE+uTHHEm/tFF7qgWjaWmHhT
y0uHrj5gf288z8h61v37LKjIGNmNfOjtdFfViLBJimD3PS3JEUupP0l0R/e4o27aXQst0UZioCwE
Jq774NnfF3yeYpYVA5Q3E70X8ZC+yKcza7G50u0Rq4V7gY7QmmqAqq7Qbi8W/xcaMqqYUaIBCa2H
9v0KgbkgfkLrvSm82BbQ+vkAco/2W4jIqHchzmjjDfI9FyQ4EF+h3H0QbGhDmFTT3nxpI2M2fGuz
QiX/Nl2/uV2kbeOPlkFOnicZjoVHU7VSy3B5V0UpVwZ7WMKlNXYgrh7kpbu22uiuvf/PlKoAYr15
CCQOVhIrR9LFaElbuQlr5mAKwsowi7WE6/Psdc4z/AVkIPPFhrWYwUnK9e1ResHZ/X+W6q550V8V
5tMEdIqCdQdhPMOKFpMFmnigr2AZyQhB537ssHAwKnAPhmSw7QluukJB/nTW9f+J8F+sEvIJIf1t
R6UoVne81oG4nAVzfImmXWpSQJ76ieTbIkXMhnVpMKkkjNzWpjs7+YpT/7Sb7AlYN0viTCqDCXVB
qJhIYfkrmGnzverYybab7UA4rn7Sop5wb28vls4giCoswDgmcu931jO5+BaV8mKxXyjRujqw5F7i
e9LxCqVzCjvharYRGjI3lk8Ez4qdqmYrH5jZVA8o3Ko63nUl4iqOYyVk/egHcZ7rIV0e4ULsaZDi
vE1u8kms1bp+JXrokwZU71A7XdeBu8Cave2pLPTeTCfyejjhx+rffOzJR1PC95MELGqtbB9OESD8
oWXwjQJr2tswFqi1/L3fHHVOMlQS0/BrE5KrP4fo0HMO/EH3/IviwEBPBELuGrgBf9DxD/lr1N8H
7fbTNbVwxra0i+9yGsy4Q1EyLwzyF26gg3bRu0ozT398ckZnsuTRLeuFalExB/4xLYdeoej61knL
D15nsgJEQisgXS7vlYTw1aBUZO7T28hfgEWYiFUVp0X5l47tz8jf+bTHcV90VCqnR2bdBA+swxIU
ttNT5MYAO0t6TIuS71k00dgwI1qix3j8MtMoyyJ8olD9L22a9uZ73eKm/64XkGIytowTThNSEXzV
RON4yM+Ez425tdkPEyLl+/apBdjp0xxJpYs4GpypIjBei88TVlizY8Et768IlT8HMX3dDZz4/BBU
evY+Z0U5ep3ZLt0jj9dgrC9YkUaRBPyWISyixI8OlgXOGM+15uULV28LV1e6trJcAVObrERH+8fm
6SAek/Eh6k91WeFAAvjMs6hw78GVV40+kQm7Ov8S3qZ7wgePfFM+fVR4XE6k8b9KJUYW+iLJmvrH
+xvIMbzLc9HyU2p9YqaFRmqIf7MJN3p8mUx0E8zQc0lG3fZVMaKKhRK3M02ihtgQm5yGkaVwklY2
XI8ntgFwkvlaTolkqBjbWoa+s/HgGELj4CPBAGXDUzDbipEzxz+3vPKtnZeqsBJbpkmp5s9dTaI6
JXVffg6uBvdTPpJ1ki7ypKB9I0Y4zD8wYIN57iU9HZ4eRZPVmYHJWXTgUcBshbXz78HmsEjLxuz+
6vmwdnTRYVytBthZcF3djn/uCIPyUNIJNOm6w+E6pHQ40xip8G+1MZNinj9yfe5pW5zcO5OUOcHa
v/N7VxgMsGeOGPp7oNd0eyKj0icIsWApBTEm5K2rcPAF5eD54KKPWaj98uOWJBL3khfQRgk7Q+UC
UBcfEdii7FEmQ0RP0IH0d6rxbeI48eo61WK8iqpsv2E6p3wkLZgJbZf3VIQBbxeamBHZzrwlKDpy
NhMjTsaUQvU1i0SKbiaoZOY2K7ZGVIkoJmnEZVCOaRj0aSETRC8U1qRUPbyP2AEDKnuSnMW7Hb11
8XHBUvhLBmQw9E5a+UJl57+gtr3rHj/s4Njc0gnaxMiKla70aSRmOl/vkyZ+WU/Ci5CMzCGkmWGw
fdcrGNgNdzQLug8v+EmWA5B5twEomdQGxRYABtu02Cb6yEQYuZiFi+pudlwIw8qj+UsgmIP+akOl
79TRstj48t1MMT5AxWsEGmE+sA5GSz/0BKLmcdbdMmK7+7xZmQ4lVE/ZdZb9xQlvb6jMacmw/Yq6
p/xGlx7evsoMK7KIE+sd8N8eJKSGl9WfwV+pPSXXAs4ZMuIBsqXvu+DuKeQUEYUyXU+TetYIlSLM
IJikgXJttEtZG9v3Jkrbz3zmxAPWRf66wkYm/Rf4iZx5FIsp/A/iMCa+Mwv51utVVkyOFPIVsT91
/YEwgAEt8pq6yICTwnU24NzL16vU0StZDDoIZ8ODdI0s/69z8FcnlY3+jOGgzVMSgPxQI0iRZzon
R59Td1nRV/ynrMmpIee6T4UqL0YXYX180YsUlBHu2Pzi7QSX2lDmRhLhQ8fICEuv/jmHkVtGtVmC
gD23We6ob9iJXguWmLoI3aErYewo2qCC9whBIM2JkApyEhqGbxh0uYtT2OWhsZ95jxEEEOoPrIx6
KLFC4gg6YhVXXDJSMJKQIBSTI4DUTOGqRdhyuyYlD4ghn/6IuyBJfRgBWRn9C8o4F89NwPpZJ7PU
uUte0SgoZKWZBmQtVAuVlrKTxAzxGXAwFF//aP7WJ2RIBBOeB0zf9tTscelouWTHSaOJb6MourMH
8D8ADeDred+oH/H9cl1bIH640stFAoBLitw2k8stMdh8iP0OpUglJm6l96N/XfGgH4bDD6vnJVlT
DVn3wjBttskTPgdB2LcxfgAwMUPn+hWOvUFMX8/omWSGmxfx7AfXZav6lW1wHLtw4lZK9R3+my4U
IJ52mVjOIks6xBGthg6bJK71/uXa9M/9tDzHpgLClZryG+4N+Qc0BY+mhb/J7lp1QVDOdQs/oLM3
ECBlHwRJGxIAbp5fU36Y4znWeCVJM9ExnBeqlym/53Rsdq9kXk8YwWwfUOJA1w58TCfRkXtrHPto
iQG+J7CTtONn+p7gLtQTLh27PdsXDKhkAmNGe7ISZ9V1MkUIEh3EpR/WfUzLRp4Sq3C92GHB88X2
RkHJkLgBvZqQmtm6HQAIdD699smcp4P1UUphv8P00dY2VAudxggn64xNW1uWDJH40zqcHhUHsEQM
r3ouhw7EIDPprmYHceideZNvMPiNC4tYsiMWe5PBTfI5M9IlCdhsnKG1AbC6vzGmlxfGCx8iDcW+
Cp49Xh4Yss0FLo4+EAJWoXSm0K78+08i2K7EvK60q1OWgLiAW7oo6rkDJmGJsrJ81iTViNZXFtb3
tmqboLEOVZm/lbSlG+C2EbTYCSDb6h9MSJBqh/Sie1DoPeanJfvMFCTKeWEX870DjJEPBCg1tMwN
4mSau+xPZrkxStkqh1zlHATmTfbaid7e9301QnoHs0ybi5ei7AIAVC9hoEJlJs0XSA/gq4+nDmBR
aqnz9P3ttym+l1/ih8QA6WxI/7+mVhCkCslclgcx8QJKEYxHfAZQiP3WbilZ6U7Vz7zLt7I/+E/p
J+12htHDpsi9VX1DUx128qobnXqa4/O22tSxTtpryuzSRvw1fYgX/P17TdUeiQXWs1+Ta4M8lKDy
q77aRsTBdK9f/aERvIftP4CGiHjLw9VoVUuzFacadAPawLQEx2r59HkdAs5waq0vhnH9EOQw+zpB
fSgxWLElYGLlwl4V8qto7XdMCT3vhSvNrYxDbkTLTp1lzFmYYwIpQfz9Je3sn1bPtbf6QjfLbb2l
9KQCCxG7X3OztJVRIYRoGU4EAdOvMSTewwOSI6mRtEeIFRqs6BkjV3eRDDh94IoNTeqJAzB/j8gT
0NMJwQCwU4251L1gcI89gyu4WR7U31NYBtDHdZCvH4ZlkH4TxwCd8DGS6AvZtmOsmZIhdzjmluEJ
vnIjzIVP5pWdaPd4ZxSckdSqhvb6SA/If1o35d9YrV60Jpz6nHNIJVt9JJ5t3bWaVPjTxJ7edSJs
/rOZhMAlsk6/i4h7+QJaojUVtDVWuvXsVvy5TZQDQz/33vtBdnt4j/caCtwzlrLr61ATSs11XC+U
sxp985A5cxtM0bY/Y7nbOvbh90Ex67RGGeWBiH0QAUZQuQmUJOkzR9n7ed+eZjELpOLFLSV054n2
oJweXg/TjY46SKmXfvZ78Qwhbl7kWTZMZ2/hZiDrdePAlcIquuNxGRxv4RTfOh9bUtGWU0VYfg/A
eqmrk9c2jW0JJ5GQDKaS22IdHEo7GXuoKV5vt4Hil+GYK+V8bUbAvmB/bRw/Yp/EHCuV2HdjOVUl
kBcSK/6B3ceF0alcWpW73JG+C3Kz8ubmaIWW+oo+OYT5skr/kBuPvAAQU5iGmnj+7GdpvRtxN8NB
IzPZ5+1oyHIgLwpGjiltXvt6cANchWLuTk0yk6XJYGk8W8GmT+UnZmUP1ol9U21INV4BCsirz7UJ
6Vz4NBr+5HXVBVcqdfUfgQuC46fL5PUVVl9fbKJ8KW+rOkwb2uCjh67F5O8YdirqbTn2n8ASDvLR
3EKWcmxa/4cyFl9WlAhYUEsE7Axv2EnelbV/3n9rsceEaF5Z9S8xrXfLIcrEN16/9qBOWZ0Gjvg+
fmv4W175POzwx+Rf3Tobr+OOisj0LlrlG2eLTpU2pc3WWxEfNfkfTKIff6rzmCw92yb9b+QwBDu1
g/a6uMP9aJ/iIHZ7FXzIktLf2SIrLs7avldLhmkLX12HIrf+DPCtKDLDwXc3tut1xnu+ktYK3PF7
fymsr9EVBjkQQeKkUwIz1HYAkl5eg6e5Mv66qGZfAO5NgirhOI+wedwUw+IKv5efl4g//FpSsO9+
4lnXJEIbbtIZvJSB/pJJm/O06LitHf3IEroH6RNKA+jtkBdEz1lhYOViRE2ReiQzKJjNK7wWGesb
3mPgtrHVciRdPiMCiHjnna0ZyGHpg6h93Jv9F1VtRSWsZ/ZFQTtWukLP8nnfqMp+nEQa0JiPkXZT
NnDTmuSchwA3+KjHoRffvJ+M1ip01f/cg+1/nYwQzy29AMDMQnJGsCkGWR3zp52NhFf/upyfSHan
z9utqXnRVIJIddW9l8PE5oWpLoDyi+FfXa+1byPTYR622/rXX8FEIDd9CfxTUje38ZTX5rOGYVjR
Pf+AKGmzwLCdXQ1zHC8kvXXIwXjzNZJV2dy9YVby/h5QQXSgAksJ0U2URMAyuX8mYwzjB/h5rnnk
VfI8AqR0a0YMAmman/QUtnqyWGsmbdH0GaLAScGxc8rxOEL1J5riDeOfgPH57VDCAk05neOCP9f5
Dy3atJpU7sNO6njEWpAvmujgywk02/vaRTuzK2KKa7XEDh65r2WIn/c1zIQhSO934eVUWGE9+aSi
pLJEh8ARyXm3s8ZbQziBFaMbpXBqHwj4wE2KQHYSqpQnSLCsBmAH7HjAuq66jLpQESN40qvRji1l
SEnEuwvxV8BOZG3vB40Dj8tPs8pglpqwdF0mDa1gdDVfEBVCCyC3tkYElvdMWOZVDtcEIcCQM4kV
kZz03kBrF6GKZPn+0doKWDJV47M1B45WsZbEQussFOaQV/VNdTJ2ZODAnFG6ffQLtOKjtib6tA2u
+sgHTyV0ZfKVJjMqz9m1hkeA7hvTXwvW9NXHLy4xxucSvH0Dp+fnM9GLjVaImCy3LPlCNaIGXRTP
K7jdMjQ9yrqqW0cicpNyieiSqJ1wjkF5h8SYpT3yECbMoUyBIU6MkF7FrKS5G/TYvPTuG+TZMRx8
2djRoQo9CrSVjmAQCPfnBzPmkdBSk4LMu3OTKLIu7buJmaGiLCy04vBMHhSr2urQXhINqPS5JIvg
z+MYo3ZU7DQeVPSq2se6x3RHd93/SATfYyKT/O//MW6luMchb/gq0x8krGlAhH7tY4FEOjS18dDO
Uyz4Wv4D4CQtvFtINGjB2ZsmrlWsr9HnpGsIsYE7B4eTPw4TbwLVwlFHa2ipCH1tQhaPDpN+Kbh3
o+pbuzSkSpcTsAFefuCVTr6nS6wBXldTCobVTP0d8FT+sjWrMbssdFeawD8Rn4KJfdI2Uq5WQLmt
1Jq9s7XioF8twr3S0GzY/5RbZ/NoKff2QXhJ+hnIxt/7Yc6fHWAUe3c4bIzOADTPnJ0XantS9QaN
mJQN+VG9KCntGDYjdUq7Gjd6It0yBkhAYbxwDhT9Un30RaXYXRhdppPbSWv3Stihxly19yI4YJmB
TqAuUViy5p2fJPDyE8D2tI6QB548+Hrq2iEoMN8jONfLtcaBDwP+viIDcyCpj8QuwdXyKrBnrI/s
Hs8f1XN4g83E3PAsukfB5nB8+qeG8iSVsEl/jngH4Az3ZEkIRI+8qvDZjTWgS9fNVA3j7IJA+ek2
DPYTC/n+wzx+5UE+C4+CWCL4XSMOT0EZBzswMpB7XiONzyzGucM5xNZ6QG8PvWoparKFNkEVnGmG
ClAxo7oCT8GWrKZJ1a9SZf0F4UjVzxowak2x/l5KVJGQwlauCyMTHKi2o4MtUpJ4Jh3AuFlpq1uB
EmPLyA6WgVCy1CZWgny4qT5aTFZxLQG1LKaEvbpaYM++hw3g0F22KxYLWSoRw/gGmDCVcSLiHIqw
RFNklzoM8p7G/LqjKsNcy2/FgEYSXXSLhChawknnlJWWn8s8NMW9ye3nzY31Bt1BAvlPjGyMsmnl
arTT/XykzC8sli8TaKNZ8BR3gRXlAmBly+f4cEB6+FhWS71J6r1BOAg6qO9O9zUUaROIw7peCnOj
7goI1+7UmUy4sGmWQA2vjjkZ6580azRF02u1BP/LyD6E8LiHfsJ9CwPwsP+q0B72z+rws6b+TFQC
qTttXcKYHFxkjdkja6zHEsMe5XXRHp7gFb1r1YtvSGiT9iWCLixYFlQ1zpdPBldcy5+lXCjRaxUy
c73TuykEpplYb9J+UUfUWL+AxwKEY0agK3/THY4AXsZ6QElfsgt5TowPVqlZi3eS7l2162D2LGvw
LOnWGd5vSWdiQfSRErWzjCKFxU3JISDkmX3EWGSTg+HOXKYw0dlRhqKjXah0/Dur81+U1Aupzyj2
tKn1zDqe2G7hRcFOhbdXADR5WN9wGGQ3tfMknXX31xRrgg7VbpluH5szpkaVCvF4p6f9RnPSefSw
G8Tf8F+ErWAXBsiGG+RsxhmyzPmktzKlbgQ3i4N9+ciK0O7lrSTTha/wD8cMBPe2zDT0Jco+Sza5
4coahUHYPLmjYoNjBZ+Ee1Pi3IqXD1Waim3spJ31HL8IZZCTAhBu+50pM3iHfPj7Y3JAoI4ZQjop
h0fnixs7UPHR/9X6wHPe+htO3cKC/ee1J13uj1GaPsYpQG+551DgUZyoABATUa+BWsBA3ySbKVDN
C6AJVDSvjY6RFjTIkBIpYmWGO/hZLzm2sT88UGxRXGjTjlxF57i4JL7TIkGMxYD1XsAlWL1ZnGDY
RMyyVJD59n/q3hHdNwYFQipbvpoLye00gOYvz/fE2C6duTELldoIiC/jM7FcDgnrMUgKe6Bhk2fo
FnDsx9CqcjsBU2bfWQsKdNPCAjkBXSYiZR4GJKs6SfgWNoJ7WkJQ66Ji66WtDAkXpi+7OtNERTj1
LS9+U0v1fcOWQivXJIbaPFT5OS/sO2wZRJRUYFmkLB+ihV5clBGB7ThY2Mp+6WpTeyq1ZfIhicGL
ToKCFF+ZynEeEJIyq/m4LypDK4uNfNURI6Dx2fpdiaA9oULjjCcBOlERmH0SiQBcbsUfyxy2hyu+
RgeVbAZtkQW8x3BHV50UPn2ooCZVkdIZcHcHjdlqHKZOVIRO+pkeN7E7dVt9C197QqoyYATiO0vr
VWHF6zd8CGH8NQndsnanbKLiMcgoYrAsJVzxZMi6Y4B5iMq/P6jEQcV+SOwpSAy37tZIZLbvV1UP
QgAop27zVqZejkXSh2LJFszHeRbzli2UgJEIpaQNoXzTA6IWej5sM36g6KrftrreE5mXMREhY4ZB
TH8ev6Rjp0Ms2/j+qU0jOaeMB8Q6DR5HKKbQGZs1ZeFUYI7cFz5Il1tD0yOTamwMgLOM+EjlkuLF
5Ipz06kmtUPhuEbOvy0leodI5MxczXWQ53LjYUiC4nH19gTObesb8LK9ozzcPcLjzARfGbdpbOCA
DgcGwkatpT9BE7Dn7D9y0iPGTROiRygfxQhlketibbmpHSMM9dhJJLyK7tVa3RTpOO6P/5Km4RFM
i1AbKDfCNM8QlsB9wXB8ahnnOvtoygQBvq2ijomwje+xzJnkA9PVvEeLrFRnUOyZ5Q55UIL+hp2U
YD2PelAyiQqO4YHZS1FYw9O90Ts1IW3D3ghNRs0bcZwIziKAkBsQmMApEb08oAMqsAnikw1Mu6FK
kVzMkUipf7nE8bmytI3Ro1Ce8k3vvaUr1xNu+3gryGZ0pb1QHHFq+BxqvTB6eNfxG0ckax/gzztz
9VBsZALXyMPiwuF/Z5aQl3Vh5BRf+BlwSjIgAQY4AhoUz1ykieJMttHbsXZ+CCgILGxNg2INljo0
KcC2GPqbkpDgTa5toG6Mkvsnc93U+x1l0FJB5Lxt8Z0SIHQkAmnxmGjkJkJBTBp7HNar1kvhpI8Y
GpneePnM+893c/tVU1f7r2sLhYRQx4onbN0cij+qA07oNeASyHDnlSdjUH7ewpwTvKlFJdW6OUvl
iTzFHttrJMXgoekSqoNGJR15iRKBu8H2SrJ0hve5iBjgnjv0t5V/2mXqPJ4PjNrXaXgL1zWbwyyl
q3MaX7X50xekyxyJ/Ssjb9DGddKRBtwM+PU+UyF85S7i6u3s6hvaruBzhUkgfPB+47M+TChykvtW
R2zj2McRRqrzHaVARRt6Jkh1n404Uxtfzafl6FoZFbM8lN+5J8EwT5IVnGqlrEexnpS/PfMlF15l
Zyt2XSZHmTHcUXtIe5d1Qpnr2sdVFKPdQPlqtTcXVBdlDtTOzpjL8tAvKcvGaLufAwt8EkspIc7q
aEpSbJJdLgm+AkTzKRt54Sfpm8bLfwTdVBwvXX17+lTKnMkY4k1uycWNZy7gzbLBS9DhlyaV7Srs
Bvgg62j0sdmplYEItEwJHK8sClmNP2KGgNnj+F3PnynHw1K1EarSATiKoh5s6e5VMy4Bxv39JI7P
SPiYFw2XgXMr9PMVWUb+jlFigAZHonk6SY1U+Hxoa3/aFANMlTwibDwRwi4yL9F2Iy/3gy82quCO
gvPW0FQz5DxHuv24nBvGqabY5ZfRZApWOt3nYvKazpfp9Un70NEndpGtnKGXjDILOr4PmxaS4qHf
99kdneWokD7pyxdARLObcL0vltcNLA2y7ID1YG07+IRCeeT3UPAwOgGGxGQgykXwzIVkZ8Fqc2NZ
YRmPtf5eZH1ckRGQzUSSNEsCKapCk2HUgKwrHXMa6T7hExettRDAqYOavNhqu056HsHmht3Q/7FA
1xLCkMheyPnXPO2JDxHzHjZ5GGJMkl2zIQPqVTqMO9lEQZY1sqxVBhFtx3zVpuaTLvvYb9nNnadO
Oc3kTYz7s5h1w7cOzSHOkKmQPaiWF9/Pl7Uv6KrCmhR5em8cSnrH5CRFiclQ1+4ToaExjkB9FgTC
LleOaP9lch3DVcptSzbnUNFN6xtnSyjuB5QeW6qerh1LwUtRLeMMDrCpLjM4bALiuk8KsJDanVAj
WDZFVT50l4lbAsvHuUo3ja3gNMmW3qBRROvf0DbgpbGlNJshmJV7/n9xhB23QtYP9s21ZGRrY2Rg
r2JLoVnZOpT1eEp1XqqfTfZcVDy03j4m5AsidkucUgCmhiataThQ2I7MNUh/GBni7bpPWGZoi49z
RcVGdNUZ6pZfaYBrRq1y77Yxxv8MQXozBm0w2YNqrDYiFIj+fJXYoP8OV49jtaUDukwNxcg+Afog
1OfmIrbFo3n+RWN6xhbP9dt12R9usvYqWfYopbrNdF+OZ1BPh023ZGBgNTdibYGtJG7iipGsk50t
CcoxrSYjkjUbugoP91bfIC6tis4ryjYMRnP5ZUO97mwLDCGI0BwGAbXHr1pA17S8aZz03cfAaZ2L
XeCOXKMm7U+uF+opHs58vueE59toeGSuhvUYSYeoTY4FlfUpISmbsDlvreZzS1g/DfliTWgZej2Z
VM3ghPuCSNDjJGxkctbIToZduWr8GKFkgijI/zMN7Zoda8Qj/QNevbIbg5ZgPqZ4/ybFIsZgUsGL
0s7j3jIJ68p82HHkOmVux7aRbCGvVvMfHovGRszBF0CGtrdmgwA10ErpP2qPKsdDK4YgJTxz8Tyg
LseTol83y5NU5VuYLuurk8crlDTCZaf5RoLCQRpuQT9sUaxDBX5bVCs4uzs8GPxXTPbJX0eGMLMc
d0SggvTSiaW6JuiDOUCzpH8gH80+E/6XBM2yctgAlJSeS+Bk/SeUHLD0NWc+bWjPZZ6RmHfvJiSH
AUDA5O7Bwrjc6qy2OAWJq8YOUXYE8DNM32UXEWJ6mZth1YLPpk372bFIu2Tf7ZPz0bi/TYN1E6YO
RDUCXFLgWXSBos/gvTjfrCFqAAkpvtfUTtsu3FKxJT83CbHu+CyrNMsD5+y5z/76N3S3FaQ2lotC
4vEg6ghcfHHnGM2O3nDWDA1o9SEJhwloxexBewxxxx/p6BJPitMTCKg30TswnaGO7t+EbytIlS/P
+MINmv9XgdIE1P+vWr7VnOoASH56jg3zimq6DR5ZPF4roOjsqtvYGUzS23iToW0zeUavt8Ki1bxt
UXh31MOm7QCEvZnDkycfGzMY3aMVasPXqz8GgfpdPX+9CvMWBT9HF845vMtpO4bd8u1m0R3Ew2Nw
YlXfBniJjZfQG2A97Qt9XlxlZQ0vjU4qhdUGLfxpk4cEBNk9nu07lHU51sSLSO0YNp74XT9fIfna
bMIoGlkXhKQInbSPnyKASO3xhMazM4Md4/B9Ty5KU4jP0DQgF81qsOXKeOBYGWq2ARAVme3simsb
U9SJ/ztQANHc0R5Dnx1srtE2JNDfFWkoSu+2MmN7W72/Zv4VcYLIcFlR02HuqKp/N4Cc6ZnNlnZq
YocGSwhUDEWfessqq5bpkQD6ovE52bonGrrfbczqfsry55Lg2gt4RkP8mEKfI7KFYi8ulO7WMsi8
JjBqfA3hS36w9SFwx/BqOCUTT7KF6A53b9Z8GihjD4FnsO34LeKCY7FJV3ojVNyIaOteL+rAhE0M
Z7HgBT3/WEa2fattOohnucC4/ffg0LJ+lwGLwepVml0mt9QybqpN2w/4mjm7r0B43unFHRjzvUR/
EcZCweyohIJ0Xy3qNr2qrKj/ud2ciGQ5I43OyRWJ7kMyS2IvBU0dW3s381ZjMck3ysm3ibsySHV/
kCXAzIOa+T+4I4Cp1xsR/3J9HmBlDUWUGpvuNX1gK8DEEvpkf/zJHto4SMUbkYZ/JnT8pN6s50h4
28w6XKjCRchNhEFmN/l2lqOufYYuxz5e+GIA3TSd4OdhzqT+D08HEXzCryJk2AerZiyHcxUhWbmj
iyX4nyo4oeyf7BeasTOFU6cs367jgle1GUidZU0jHEPgpURgRtDaKxEh8rLri/xqEm00c4NuHbHL
Q9w8VA6O8q9JD77K4poA0bXR81EiVywa/CsKPanCbwv+6Wm97lIQXdJmkMw+CKAOS2xQdLupYRzm
/E9XtbICo13sJlafrJEL+DeJdVQLapX5pl0fWP7M8XHDGh3bM/6dwTzkyGp+n/zFiEMuSk4W55mk
NE7tbPK54/wAOYKadHuscfuqiYTCXCP9DwHnxVoAKTNoEX+aO5I9jBp9/T/LgX09XR0LOHgp8MsA
Jnrins3KD+1Exb+NBaB155z6wECP9IkQrCIint4+jBRL0sEtbKc/YsrccW1g58TblUzSZjMoQwXy
kq3jN9z+GZ6xaKstnLP4exMJHnN3rLqiMMrfLKIlyDZcKbg/UeGbQJZHvqcVScbInfEnFcL/Hozt
/UKLrxqZpwgEIc5yRZSbjtRY91Nvi9cRWOdTUghgUcKM5+GxBkHGwskDvH+o6N9t/o5yQ+xvxJt0
fi3AZ7M+MvT18KQIowHqIeC2CS4TmnXnTEnSnx63aFwi0Tp8+k+A2nkZkLw+/TJA7wQeLWwDodEB
HPCBkwGGuZOJhKCWiQGmyoZ4jOvWxkacmjYTFM5kAveVPamhF8eHnhpWxPLsVjYsN9ZkJb20nRNR
BiY+mxDNvlEPxg3PQqXADIYGaXKCsU05QGYvRMKV0jqciVEV717SH7og+coyAO/hU1Lj23THu4+m
x6ik7c4FXlGGXQOOJvV7ZhaAjOIE4bkutu0Ndad3sh/PmfDqi15Czby3vXnLHP3dbWakPqrxB/M1
8N7oZ4ypqV9wNOqxqYx40PP6h8KoJI0Gr8r/datMXq6Fc0B3le7gR+TVo25rXzNmN8+8eUgFVG23
1KHhV+fI7u69NhP3/9pRtA3ZDHgUedw/3ht9BclJQUOx2efR5Jq5aSqJdlJiv2Kn8J+n7i/vxWL9
POoHrmpp38YhpEdZLyePPCsx4AL9els/NFXxwKeDT703U8UdoQK/hvZ4fFMkp+6psu7ffQGMM0nz
CDpCDlcBS7xD5MrMCFBkG7Tauess3eFHr0JF8069maCaFshcpnuBKDiGggSoEvHzegO1+muh1+xq
sMK8g2Dwkjx5iR9UaETCaNbj1tpYZBie4qXwO7499jXmu7NlNfNBO0TKueZvTOX2NvrJpYw/8Uk5
YRdedzjfOAYqVcw4DgBy9x0U+uFNcLr0FbWWbc2geSkOWopCMOMgSg+u6rBCBwy7nMg1Dgz5oWqj
iwN2dfwNh5/684xwXRxGB6IZdk9BhIkDCpeudBFRiJQePALWC7cevflijgs3DybXVNtSMuBfCXPo
Ld6cM7SGjNXGLoomQoyF70edSVKfEo/JAFXsLRv17v9yeluzMlfP1gRvvVhjGf9a0qevGIBWE8Nz
+nUiyCmJuu9vIHxq6RjqrhnChAKwaPS6t2IaqES71EKe91YdRhhIGCHI/UcOdL4VASDDXlLc3voX
xIHFN7RSXFfnSVL3eGXGbepsf+7GS2kByaUePVIGqe3KC7YATNbWnGIHqbb5ChcwzBM9GTjM2u/o
+kajPgPSk8OelM4JfSWgbwVTvi1uM7G5zjD4FamuQWZNP3O0eRMGBfT6SU1etlrvyc34XfZ0kSLJ
zED0t0yFT1RAJFRui4nd5AKSBdJ3yOqBg9aKA2QLoFz7J10gC4gL0VHyD0A5QVOxix9XklKBdmnl
zR0gi0vMHk/QqY27dG39a3IXTpZAcd4yPHSOXNAzaq1TZGxrZJgsN2Dyb7qwWwWEvQohp6fOCndE
SXiWxs9q1rCurZmOhUGva00xNZ95E/xOy7upNGyn2n7SVZiQyr22mSLRAMt0KFi6BYleLHnf5Q3l
+CKbQUJt1MRBMvAY05sChSPkEA+q1UQyqyGcQCclPD0ZcPBswM3mAf45Uwef/6JQt6bdgE8CTTrG
lgNCCZlors3gE6pveCjU156pkqRxBpS2ilolJ5+iR/BQxqDudIItlaZkioIahbXvgS/nZJbrCBxm
cW3mTu7TESDzXvXgG2pvAo48+0mS79dF+UkjO5/HBSOEfMkCj3Y+G3eXv3d5Gk2FO6+8x0cnaJJp
esbTtqeowunqseMOKFDT9H9RXPGaIeI1OtOVjgVoFGZfcixHS0xXReXDzOf+FCls2Pp1VlBJ2KcM
rA2+Afg3WmKDLHZwKOlKT1B6vYfH8Pn0DHvtFOcy2EjCWqwGM/+ef0+5U/j40pZrEqB7Znox2zQ1
2Sa3b58embmxVSz0NC0Mbmwh+PkvFNptLIVVkqzQTF5nweVBAc+WWBg3sm3MEdBwhZpiEf/4vDtX
csb/s9l8cWcjyCkmdWj+5j26+LUFcGa6Y0rY8vmYu2WrP5grQvAfJKSHAC+H4rdTBY85p2QLQqNu
XSw1zX+LjRSNIWwD5oBatnMYOOTIOC04XEZfT9zzRzz4Gt+XJejc0AqwU/c3mysw0EOQT2YTQPVx
KuImh+y961KEA9VYG2aD7s1oamm694hWJDxOcppd8DcQVOrkA4PC30hY+jZ2UfFG5jDboOGwN+8H
cmTFz/up/sfonoNlS211NC3XEAnCZY1yhM+Jr+LcPXUm65m+rGqVfNFz0uXUI7plKKu/UVhhgVJ2
trnFj/6GnHrcBzKV6CKlTKEjOUfLdM5IRg4a7M0axJ4w9WN6ek7wi88KnpLPw5wf4pXBI4nj6AA6
t/n+eixk6mPJD52Z88Rrzp16WdD9auaXFG59qxTKFpMGlbpnj4Lwr+SnxcW8KHKgBoxiC721U0rZ
szzoEgoXD7Wd97LdIgjnv8gJVRHEsvKQtAspOy0CdPbJKtHSFgw6HAsxN6H//dGK+sOUABLQBZQH
6FOypaXg1FZd5jXzX3WBPPG+yd+HqzA4fXZURPKC85rI51cgUIJPuuA29TkYuQRFne9BG1NCXA69
9N7PzlLJo1+Q2Jv0h26ZJV15CpbLJbGfbNStDdi4tkFXGR51KY7Xd2MqhYnkhfoTfOWK1S9+qcJ3
59ODqgWkfaMAMEP7DbLBDrL25AxSwcqs6VyJZvUiEFj8vIY9WoG7ZUWWFXX9mI1QE9thLWgSBXF8
fL3RCC3pTcHY8z7rR1ynMZEV2U53NinDblIWub3rcGsYk0qoAw2RxygYDQ0qZKie3mJNISqWnz/i
C9dXN9xoO0GJ8A+MfCPUGowIyH4igQ1AEahyd/dMe+gN/xNc/RRYw948MG6UGZXjLHu63hNXv4Gz
pd9h7fchF15/bkWny7n9usyGSXMEIDJ6iDG73Jjb1qv1kUkUSd7i+G73PHvS17qKO1+g+0gwwHhA
e/xw2rpBhX1n+nN0XpEZS65tEcVCJDqlhGvmQQD4/HHtVPGLTo82tuWJcTJ+xr4E3hbrXwBT6SSQ
r4OpUvbxv7keLiZMJnxpyK4rpytWpcYlsIC8OyXGCiG+3UIzAaWLELIg1ZNYquy6tCF4kjlmTFIT
FWjQHNOmtBWV5/0j2UQdaB9AEDQQoX+CTM0WE/vMt+BrEHT49sXpEqfNM2dsG9T8m+2AXs/wiuvA
uDv3WplAAIisYEtnmIrKVSzVp4kXK+6jfQYjatZiknqE8ubdDcEwYUCqh8cjBeuzp2E0L6xF1H4x
EuqwuSDHBEhlhirZnJXYH05kSVWXHdT7BnFGjPO3yqY3BzVplm4aT+vgPyhCOuDnH/GjeEHqouIc
BhkTYyJwo8ZkrI9NUnosrW4r0MwVN8A522wzilrr+VXl6MvbeqEqoEbE7E9lpNb3PRx7rzvd7GPX
kMW+coVDM2avsxc9amtE7fN+I7Xq4PCAO8Pk1nuVBZ6SrI8kGc9v0y2m/WaGhc12zEEx17DPC9Rs
tpPtenP6P2bPiWzMCU4cFv8HOYyEZK9aQThFu66FPs76kJSWA7gmtkGFFKhBtzaw14OJZtN+iJ5N
iqZ1qmwZEwjM79F0YgqZygy9d/qIaR2/DzX12KBfLWWm0O42eyjT6AFe4ATFlSlaC9x9mTIAktNm
hOoeeldrJNs1RgLGnMfRQ5YHn29xOrDK9nCXsA24TJvXGTHUez7eMYmg8Ozb/l5IY0Ny/ncHKfAj
HvuDHUeIxBczun1V3HTASdp07wSJyf1vaMH1j1aQuYK9gWGdZ00oZqVlgQ4I+qUNkvnTmbSSlltY
fVBtaVPbhFQW1Y/TY/ZiXSz3KNMDiVZT7MC1HxD2NEMJhlvudmfQKU1wlW9qAiQ5bAK7L1a059Bj
S8SEZ1Ms7vDF3QHVZ1KssUJXFgiq8SHWGAwurl9HJOqooT2Iq7INBk9rhgKIsh+Vdj1gvrMBCVht
HTE4rKthBver0MFi0sVqFjRr7/LcHfoKPZWBC8GBcRa1DRlJZpnZA6ayvjOX6OqgoJ5DDlngMONa
S7hgMkz9vwGiSCmywKtS6bYdVaHBsEgmNwE4FopD9sOEcF5/R8zbCQwpmuYzruhSRu1BX8sAFmFj
xldudJGwCwBmsHQgWcJCmVJtp94IPOFRkyFn4FovPW2Ojf+d6PjL/sg0ehEdvL0okfk3altvqYYr
9QngbDO8E1+RUP9x/a/Rt4JnOZzunN8M81WB3kBCiaeDTlovhYjNlQP1LlO+RFwHuqKJPbYpQhb2
1FZtw8DQe5Kw+fA/DrMCZYcI5Sl37Xc6tKg9Ud8U8iq+gia6oYEpBhfyDWEGDtVMeWcTRzlpdusB
Q2Grcg6lVL803JNHHZnBxXXmy/Ka/SBIwsnnxqaoOUd47ny0qy5F9fVo1yzHD/XbWrtgI/+W6+yq
FPVY/+Z7/7AqFvqey7INPuP06fMZLz7cQqmu2MMWApPUGF2B3if1xEme/yijkHlIptLQeWiED6JK
yYlJE3alEJQWBWOeE6dtE8BmUWNHeGLN1GgNsFmFp9MdxJyG74QA3k2XNubnJelPTxBJFoHD36u4
q2k8+AoifDMBR+Du4iSHeKx0rbHuvGVtkS39yl4agRDZy+fWVfZ2ZJrW6fdxfzqSD307ra1IL9rR
e6LoFWog1EYIeNu6MzY/PzFWI37f5QcAcaU3Wyuz2PeoWAfJKlmibIdaboOL9TmoWks/KK4JQm3M
L1qJNfP96nXx9yQLfl7KJ7oMvO2ayKtGRI9kpNqzBJ6X1suWShlwqc/o+s1kTVDDXbcio4RqPCiA
6Dcc97hcqtCoWm1DjGtANbOZUW6cfsl9GOrpPoqcdjo5tQUKQU/iLcEKPM5YXoDwO43j36BFl75M
DcMCP+PImqoyMRZMJuchAqmnNuSYRKOanRU4Dui4B8M5a7DzwDBQ2byqtj1UbPz3L7wTgjfAbPQN
5gAGxQmO1WXBmJ7P1srb8iMRphGzGMdOWKL/jd7GAMtwrN5+hH676cHagoFmkSxew/DRBiPQFLnH
WpJ2UB+134s/nz8wi5mruioOhuswhCcroO+iF76OXHofK4e30MllhQrZ+LzU0CrjYlMG+2+o1Op3
lIUsF4f9QEvK/W7ELVn0BRsS0hUOhME9dHxfLYkUvAHEeaVMfJg58QIjh5AurJZSGQEWMF05pE+S
xW+yz1MmPbAsvbGpqhZV9Axd68nFgu9k2wt43uv8Rh65F+8WGextpayYXr3hxc2Y7sUhMi8h+FvQ
qVcURmoMd1VpgOklJoviPh8VISeQHGD/jCeUHM5feEe9sVqqTbDM+bgVRn9t8Q9h3ra/jWDS/ns9
9yIGGZWwTooE42ADUIyKucZnQ3FZHbHH8J/F8ug3qnjBJe4pkPN65HkzVtUwpfNOwjL9bS+/phX3
irpywDjjA5U9XxMElYxNbuiGgWydzAyrZSloPIFKBcZWZiKNrrbp9k7CHU4F5IRVxy6TeIlRzDoZ
mYoa5TQcisFaW9MRxhTlwWiueBCHOv4joqVZHV6dzP0NNbi+FrC8OVKl4pXHf0kYMg5PaoelKrLF
Zp8FDy2JG2Jx+zWOU/i/MPOVGAELLpEKWkt30s7S4JuF3wW0B2a8K/sj6z4i0X3cczOs/t3jj1Nm
KQyTMnck6Uid0INIiRAl91IBQs7fjxQ17/u1Z7duelJ7tVTB9X2r95lw2/UcRjiOQBguW3R5dTBf
y/aI7iP5quvfb0FLdSyDABvIFwv/DnVKQiFAH7MHaybQrqaSF9TaAm6GhsHb5ExIr1IxGVVzauKj
Ev9F/r19Wkt7p2SDpJpFULue2GM+sqJTSGFUpGmO7FaMwezm5EDV+HobEmLSGnR3JLgxjzhrhu0U
EKicWlHUT/T/ocWpJM4hoi9VVOrC9dAu/bq+kdS0Scdl1UxwXvzbk18iVEG0y8F0zecOlssLMPQs
tG6AvDkxAZlUeprYLkydX6M6+UYkHGwEr90rVbZd/FLen+FO0DH+jBKpLpc6bMS965EVAjjKPnoi
kWfNsJpqDmqWu3mJaAFXnN9xhXaJrPVITzqMzAmRb7/FSaxgXSFhnWXpS0JaRcwhg75wOrLmISb3
DEWQ0vhfTkCd8CMweuXVmZCYVkB3o5rOk8bNYLd+lMEVGLf1opUyR1E7efbZeDVx59CJ8iFsxxSB
FhKsq2A869gZspCY0XQh+ZxRXpQ3Ok3WZkxZTujan4oopIrMmZzXAhp5pvIMOyH+ZEbFZNE9FpPm
u3zgsLadbdiKI1y1J+tiilCgcWKHm4bQ6Cbbm7M708j9Tb/KGb8nbGmdN6Y4y7zOO+ikfWTDeHJ7
xVGsMNh4D34AHqh/OMmINskbhK0xcG1X6nL4jUkqQbUB0Aox92CryUznF/wR0oT2/ywlNW+artSJ
W/Jk1w73l4yTYJ9dPDsqGhCZ1+QujE2gUmg/stw0zWBtlWRM33/DE0gjCtehLenNBo1WgwxYXjV9
l25bD8w3Xm8wo8YcXcLBbkdmL6cnbARiL81cL51qUj7RXlcxyGFD37brH0zWmbduqqo6ZrUmiW4k
9eCBXoNUtakQGz8UbOPUsjASoZPrRCCku8TLqKQO9wemCeIA9DfIkyMLWwZhYe5uWRkP95KWgsxp
jn7rsuk22IWKK2WPzwd379ByfjGLyhYgTBwqJAIP1aqnsVj8IRpQ/cdwWEiIPEu3ZX1XUc/Nd6Lb
lmjwwU0qBRgDivvaMLlaijX/yC/0984XxpP+vVZo/sw3oXby8uiOdbi7VfIEplMa8Gz7lKYqTt8Z
bhsJgFrJV79nBEhO5tfgrH+1LESHySVj8l6lcEJiFHjLmjUSQv6WH5JuZOQAbhiWELrXyIaHMmUL
UtWlW/IFmFMbVv8sh+qEBczdhvyyAOczoOi5FP78A+OLllJxA0TRNlCAShp/1VC/lbFFLLdSFwyT
PftpsnrX9w1SsXkYqJBbFFVh+k2057tLOBuNP3kPCvXF/R/UpLdbzvMCa5AOREhIGMOUiaE88OkW
Z9sRuGiNbD/zHs4PwyM+Y0oW6ogPCtb2hd7WdyUGcgvSW2qNe+mXz6DsPSQSpjy8xgEcSCEtU0Od
nkY2/W4CuHKEevMevhbYxOs17AVsezWIKshHSdVVKISFB0mJarS/Bm/jdqigipdyYjcHDVW4oTwV
FehNIs5HSIu4hTrijajiHOmYQAfzyBUg0YMwSPo7j8hpQwMvOk//BYEOK9DY/XcardXaeo2CbQnR
6eShKy891NAiN0A23AlLBBMZU/nGh6ubFDGE5N2gP4U3bdDi2cUuwWDVLIzgNhhn8/IDxOTGQBVD
raqVu4vwDTCuOWOX1f8VRqZaTxroiaTMGQ0KE2HsaF99npOjk0WeCZpS6tkBw2SzhdMWrSh+pTGL
V2UstWFN44ZW72ubYU0hhAfdK3Pb/4QXoa0IVL+bXjW1j/oKAGeBqTaHQ3iIbaYfd1B0NnTMn/Jn
O0+vjjk6rFMkaHrjo0aXZd+2PO7lTQThrkI03aprw2xTXuZ8G+YBWHjwrQKALOF+ZSOfP10PXsa4
1ByDUMaSOJlz8OlRQppScvqoBnO/b8RexaZoXqAHeVdXHN08GUJLmVw+8RQURXQHenE1TkFSh4Pu
vHjCSvjguYbAd6QUABsBOAv0vQCNTKZPTZTMTdKxeDZw19WRLI6I6qIC8xnZOTAGlfztRB3zqJ6r
pDvneXpLrzwiNK+2ZowTdfus2i4yzxAW81kZiFsHiVIU7L/mq7BgUy1Dw7z7O+nkDbyUVOfkeBhZ
I62PYNBRmtFlfqHUMni3eTmQ2S8K90KmvyVQhWVFXzY+lVnVRa0HjelewokQrCs9j+l44FU9Fvli
lWd2bav4bhfvMO0y0WfJN5ULYvmvmbvBgc0TFtxxUIjCx6Bi1vOZs18svXoIcghd9Udinov0UnmR
P8Caqzis7zdUxp5esXVIeGDjdU7wGpJgdnq4f+/mdGiLGhM+c61mtIhwRVLSZJk3XnkE66JXYEUA
/7P1UvfWvxYyjtcQbIT8mIihmX9sma6Gj4kGy+9br9rX+bwa/8j9DNuUYy6hUrMq0xnmC7IDuQeO
9cBmRi1TnSlymXlRrGbwT48iv/cEuT07Q5Y8VUULJJdGeNTxPp2/IYsi8UIqO2+zpbKEuQsArHvA
EaNpyXxflHDzoS05a0e5wDz/IGOc53YQjHtr6VScMtHN0SEgqi6xVHxTaWM49LWJPy1v61Q6ACaH
ZEfXMPwLVooWi3LeN+4l0GNeucB0nP41TH/ncEMQcGzW5K0RvhyY74O0qJ0FrsfYbyoGwaxGM+EA
wg4/tmpMfD72w5ifMukoOzpIy+XdUm43T7Unpbyp3GPMeLhrHgBXTtKwK5F4Z56OmTE4oBWNy74q
/Fjp1Tykaa1sYqtXlfsxdO+6rDTlI9kJLWZPAgdZvj/Rid0UjMTewTiCdfvnlnncUrfAYW/nm3mx
UYe6P54Aj5y9fmF3prt1eaG+54YPcRiIYHIK5Yb3vVw1qH1uOG4lWeg0UOW63x3jFnwUpml+OhCT
dBpq9QjM77ypTXM8pGBHzcbRBEhy8Tr9fCrje8+Tm/LeNBenqxFAF0/C1MRvBs5OfwiO9QJEFniZ
wjS9sHyAANMCo/GDe1a3gnW02vw6//HQFy7poHEY0/P89UkxjKWpvZSgocIn9tK8KPi752WoLM7s
v5rvPtGtAREcbIxAaif9Oq0MoXxuUX5osWKbwf7GRRN29MryK20WszVUag3qcEJmwg6XT8IxxSKq
AfZz7oVYngi8L88Y01xI+ppI8oWmqmXlcMjOI7lJYc3KvQdkhjua7D5M6VPiLuAmFx4jXLibiOxT
eYQU6OGWD/B133CU5oAo3xZGgE4O3KS+RpeGhOBNiQxAD6iycO1alMYOZhf8cUBIv6FWAxnRPDrn
2nm2cMkLWm5lKStmigpT2AL8hqwEMy4D9gGc3Z0Y4rbZmu/aoRj9QjAq6ZPYS8Euwv6/8bIhnkly
hwCGg8rZXNukrsyUaltZqpGY55TnxQGpurTSdaTUQrg6a0QweoTOZa5dzVRLKyS/Qz8W5yuCnaFP
+xZ/+GsR18XSfGMGaflybetkpyiqY6jzJx66vBMj7zMhmon9VPuxLV/mKYRuagkOgcAYfmRAqecJ
X4H5EjsD4+ogulCGHVZ4CZiSJUO1IiiBrPDwmeTBK6fYPItEVeYOStO9F+QG4viAKSU7Yl2ETyMo
SGARMbLI3XmVj9xCCx/inoeuZmrW8lpKQhg3ZzbI2XGD+7QAnf7nrRes0w8caGRIIbasnSz3mrIT
AHyqcxpYqO/PlJQJ0IUyHx3tV3uZPl0/J+njn97JSflx+7pWfbAz8OuLf7IbN4IuL3jTxHCcrG9C
b/vKngEVhQXCvv0BWS1FHqTCqBSXybZ66G4yggQMt9fd4i5vH+WASkCLZhflLFl5+lMICUw6ke2X
5fvT8CIv7ljUTjrWk0TxuYzLNU2XZS8K0puVCMj6UmISJZOx4zwgLdigmt8kktFTk5R0UwleYlqB
Z/GxWVCtKXzLUDLZoTajGuYx6fAXDBtIZ3Wo1q+fpf5gtqxJifUEP5CjrEk7t0odUSXJrSLikksz
8cwcKNLhRFAgeExXpIeSlDlH1G1Sm8Jua+AnQq/XsDrv12icHluQOHdOeHLHGUnrdt+NH9v61vFm
MXt6iPFFU3vX2Cu7FeSrPJoo8A9bLaHAfQuWTDePYdQaYDHlymVxRtIgJHCaaxUJF1VWgx/mzTYQ
rTYXt+pRvo3iQo0RmbBUZ5HhIeCa6ZSGigytyrMn3Ul69cRDDErDypLxSwPK69YvhUeFyFRHrDKi
eY7BJRgAlZ84ptm8OqEVPNHixgfXbCLV27d3RntcEY6c+jP5gSUhYABwLlmI1LhALcg5BeS+GimR
ImhSfTmYYc97y/vP+Qjs9jP41gpqY/ST/vvggD+fgl9OS2HFfUlp/gSjw3Zpbsw/OBbQcIw/fVoI
R8UerFXoeAqAQEsKYufP3Ukz55qBeNJX50HeXfEwAjt2Jtk4jO3EsudX8I9O5SswGsWkpTV9JqOC
cCcAYD/titW4JSbhPCtLIcD6Z4ndhSMGaf7MqNn8Hhzw9n8bZgAV2c6qstVNFhlC3E/zT8DzrkJ3
gcpenQaP74mYF7F3NDbTRJib+Rk6T3YanH0mUcdMyuoienA7Qqh0STxrNUdoeglxnw0VtOj3dXxh
TfLqMsoNgLY5USBU+S/LS+ks/+BcvIxUtVfguxzebk8ViWCnCvRRJ0nFhrZpuvCr+VPfWJosnm74
p0pJt7KCtlWqIXZ5FgV4JhH47ljQPKUGIsRK1Gfca5GsKrt9FOCaaBrbfUXIC2owm+/TrQ0KIkDN
TaTXoVX4C3M7r4YFZCWq6SDZqeq3PmJIR+j/bMngn1SLUX4QJ2c3CIZJYOFS4aAbuF3iyRS4jqNi
a1BWTE90AWCmtWrak7vx6CEatsdy7GKUqIafKkC49kBZ7bhhN3XsWONXkXRijyVGC/wLi3beapPx
XswmZmJtNlemVGwP1i+3IY/B16zwPPci0bhGXQNZz0gELe2ba2Qzq5/peIhfuLLWKOFN1TXUhm1+
NIdYYvv+imcqI4/Vry1ysF6JQ9QZqhqFPI9Y/q5Y+iD8VrCSD/5YR6ic3/nQbSw9GGxckrXf9e+I
xcM39H20kwjm1pZNLj+DiLhAaLeGiXKr9rlxhrJXmg7jf2y3nGNB0uq+6xZllJhkMlIs3ljZcL0H
N6uOVcX02VOsuWB8aNo0HgIquiJMgTHVzTNlTTcWUZw1aeGHtVscjBlTftnjSAP/WyJUIgo7R2AC
fujOAfjhQxhS6EJHLFcy/kCXpeHhm58AzQrHYqhWRYSWkZBiY7qVr0pm6iAR/XORyfELyz2gN2NH
oTOzcaa2yI+RsmZvwn/g/WOgJJtoJyl+CHrqrMiPXRZHnRXE8i9YUlW0xSP4gCqy54B64XZrdy6e
u+aBG+IFOWlziZHeoIc9COe8/ppO908AqMRjIDCoOYfbNaFUY/xha5VwcddDgHS0qd0EQNFslwZJ
gfilu+nB7uKL9A+qntcKa6sNXO1+LrrnRZeozsQzFnFoqZfQ6RZjxsLA0j+fBpaJp68iZSMkxS4+
A08xQNY53rkVZ7qw9jkkFH695+6pQeWcU+USo/TWajsN781liKzNbUWv5+UZHPcpnIRcOaojd4gz
sdCNwCdSjDvAGTx3Rpkv9R7hTsgprn56s+VGOHVrt1ngnIG4fRsvtN9ggbl100EpcEMR4hmZJwjv
ngIioECGooZymoZk9TIV6CawCeNLEcSVvJlb0bkLNXa6nUsq3lJiMlPgBYcbHdkAaJFqN96RQS6h
ds4CEcKyip5yWEYyU3vqaP0ICNkU5ZgZm26QTMdUDFzzb+dgxqEQH6UhFt9mzry1itEtRZOJPyqw
Uo38EGlP//Yc6RXYgydr9ol+CywkmMSRJOMfKCuTCSa5aSnpsElx+TJkelVz4rDVmkTE8BOYqjDl
BmYbCWJ+/Dyr7M2LGsdGt/36bH1m5J0JRi+xoGSDZJYwKpWBcMe017hFjOh/VjVmP6+8MPA7RuqH
T5Q1MNOLeypK2vqWNW7v43X+p0Xo6AfVj/wFRC5r52GXJ0SYSY4GRxJ8BRqdVTD/CXy4oinMDtH5
3Tk2xDUU+zKwLpFh5zLJkzNs5xx4raEgSwzgB37/ud2sFRHbtOmFLD/5G6QsgeqszchzpU50i7+Q
FAUhFe4MJyuf2DYVZsFGXETxxWIcibbzAA6YDS/vL7FmZndGLqm22K8UwhiN/2IF5+v5YVY5aYoc
1Tq/dn/fql8hnipcUVR1+W6pLOVFsUN/UhByZOgfprvulrF6a+wo1vbbsdGGlHAtUDS/nfJDFD4G
HRIDslmKpjkpGgbVJB8q6FIdt8E+v1eg4DjElaf+ysttrepv7xt9w5PBWp+ACmUX/UeQYr8YN2Jx
6exJI8Qnx0IYxo8tHxOgq3RgDzebdbFBgWxzu1BKrY6ubEZLOLwsl31leIQfj6WXH+y5rR4r6lPw
4w+MBvRrKyTotDgyRwi+g1purNpYPZwzhRAgmvDp8cpcDlRLsW00h0Q9N1Xrvc/RvRDTSPIRqdI7
A24R5Z7VewywgYs0/ispdCwiiKGZkF8BF817ysVb2oKqzzzNbFPUtTOZH0M+q0xnEYb0tk2hIhXw
KfXbMuRrhcXECYT0yHMKd/isWNBezUy4l0pxztHbwPrsT8PijKVdlMywr0LV2qVY1Xm454di/hvs
ebWutaebj/69zhzRDOgP1rpmhByGFErCV8+8OpiqBFlRsvDVKpdFWZ/6JQU2LfyZNBTB1XbilPY4
AKjngXD5pGlzbpQidAOzeMfTMGhxko3HJ6iRpEG45w1YOsw254+yPeQ8sy/cnh/WgVJ2TavqL56k
0Ms9RleHFPTANUiEVK+6u0SdXuwk+zXFcogB6xxRV3E++Omhs02XZQDQEWAVnuUlJk+FEf2OLMbW
3s6OIj6FAtCWQbeLD9Z/Hm6+zY6PuxbJgdbMBmLWzp+FWCxQx2c0WZbJVSE14XtdBKiVBttidNbS
TJ3QEu5wUAISIS4o/y0q4dDgjwanD4xiTHNOrQot9Z2r7cQg4pHNUsOtnCp0YoOz6HWWqN1jkcJt
97uItWLUFqHnl0h75I7ChKf/cKp2WgRtM6HkesHv3q1T68guKqI/KNXWLaeaIxeoSdIptIvYT8g1
2olcSJDKj8m5yLKHjVO+U51+Opl3qyaRXQ/ML6rYzUBbpJI0XuEcvFGYg8qLBQyQ7kh3EYduNVl8
vvbBt0vWwNqaT6qFGUPo6cqUfraESg2nEO0P8lZABfYWKsY1IJiV0qbBYsP6KHNJbyf3p2cpoG1e
fh8udz/rsbTq3lGkUZPq/Yo/9I0e65SD/MaVvgwQ9KJolIGAO1ARrXP0uJWXPSt05TBZ8eb1VWvM
10uaLJhwGRk1CnV7Nj12eFWhOx6gFr+yumbAi/5+2WVcX3l+uW+3KZYog+N47fyFm68+YoFDLjlJ
+qdCdeW5WOtfrnqyyRrkplNkn16azecLlX6DzHjaAW9q24L11Qrduo6Rg0HDd2jNMOcML0UYngH+
/5itnRf6PUtb/QJJ1ES5zka1H7HEWt0d/sTDjsg0QEjZrTSows/wZJCXxOqGuuhJiYYBMmd2Vle2
AonV33PlzmBcurl2pNSoy8DdTIZ0lWjY8aKnxatEmrBR1NENy4JbVkuFQhDxwHY6RIN74kJ1UL2u
3oIeatj2CzGfTMVSsd0z1MvT4gha3+X30oKVv1qz4jCkb61YSkcIUpYWSf0ijKmSU5ON13SIyt/X
1Y6/r3ckn/S5Def8EuMBjqXL/PCPcFjjD0E3tb0JH9eYyKgV3uaE2a9p3TV/UvHC9OtuTB5FuE3l
GAbkZJFUltx9Sd383SW9kxbSLval83wpUfs6PpWtBVhnBYj9d3iRMzRJqfdj7Nq3/8CiLHYgIb6G
chZJyacBmS9oEEKoveYuug78EKHDFucWpeVQJsykwWmeSUi0GjDARUdKdS8GpV+0OStUk9woJnjn
FGZ3GEIofscePwpWfzJz03DU9NrUWazADGCYQoaxffQd4WVBz9BVc5fTi2B1BgNbC91okmgS+4ZH
UJKnLrxCZBsixEIdgnutlqhRZFeNnMixeAIoMECiZ7Kv0N9KPgRFlKP6ZDvTImP4WYRqg1Ym7SfT
or0f/zO5r0cPdQ+gWY22ys4zl9MDvfiXXGypYwv01/bQbbPvCkGhQ5SlUrvw8XAUFqNXscKkmyuj
x6jCPd5WOhfJKptghtMNhCpQ/b56dVY78St55mUQ1N65ZV1RFPevB6LyWLFJVwe0kAs8KP5sf68k
00CWAuFN5/LWT9BteMAT+r2jmVYiWGwimFwxrbXTO9GTxl2baF8kL9pIGChqqkd8e7oT+qbgQoCU
hwk2Fcz6jc81QwqYfoRVNn2kmscKGZzI+DQocjy6Tl1fN9YXQzmYzFxX4h4fszY8G6sVPG/flmoW
uyqV8gJpiIa1w6szXNxmi0TtUmIC/lFE7C5GNvZZNzvagV1sacBTNaKZNkIynBI8J1o8gfm4Mir9
v95HTRGf9sQqF40HbsaNpal8D1/HWwPnb8lkhrFq5Uhx1E+oM+xoVCziBctddak03v1ouIwSjajR
JfqIAqc2RO5Img1Uk3eG9AYdIjZ2qetpGKQIWLlnW126MfzEzncy8Btid7yb3QgffbFT/UCSoE/G
j4Dw9myV9uq8sFRg0BRYSIKhZPq9Ux3OBhQ5T+1QQZSwqXCsMfhLHbE9gdAWVLeeEnAnuy/ABX8i
wLbD7LoWJnzZmRZTcwUUeZJjvGw9pAz92Kn4XAzMI7TaBVvHx9qf4p5oEZV2enrcQLjt3rUse030
O3YvkkWkONu8Jj0KffM8gfUX7/rxDWXD12kakDc66xLvRLd17e59k0F1AjejowN0ZPGcLQHHduP/
INJJQWjC6/S9vsjrKCIjhYttrXP8mHNH3/YrbQznKJk4pVWm6doyIy84xZrmuUcf1mJ02nHdlH9B
vWT1vkDzUgTIbEZl7rMEd4VdzY3VXV7xbGrm3++pIj7dyqjzEjlJ0Tbt6bYUoIC75XJ0BCiOe76J
wsR9ldvEWq0bYcwd0DXB/fV9cfJ/72a6Ob1xTfWtepbl+yRUulqnwMxdG66ZLI0zNnKWGqRhW5wg
misqBk1iKYaOw/rZTulXcNQh7Qdl0Y8h7pFp6lsqN4dyB6M//n1ZdA9W1qQdyAockfZkTqhC/KpQ
6lcEbs/YHBte5UDU0sh8bgsPFFmkVSGVSXnkD/MTIRRfxPtMyaz2v/F6hg1gNhXiU3r9756GKtov
Bn4SYtUhRys6IyEprKfvugUeBWTGUdaREgVWIHI3NUImXXubEX0kM1z9wz163WT5PIVEGwdSNl5y
zwmiPiqaHO7t8cbAniIw8L2ZLQqVqqaxiOlLpaBGGKgJswl6jdNB1uR7GeGoNSXDr+AHjHPta+l/
A4RrhLZ9Agq6d1HuQ/8ikHWB5uTaj03BeF2ibMAOp0uCw9ASuYfXJpAaP0EA8k6mXuEPBs4ftdbX
hQYICx4L3FoCPS5vzFWkVrehaCYk6xmF0jxnKibzH0vutlHJ+8Npd6e+Lk+oEN4V4afGygFksCl/
eAaV2q/M82sdZI8ibDyEPoYyDvjXDKn4B7iyu+m1iWXKpMFErDrDL/xB6E7sIH6JvcdAj4vzvprA
hyGX5bTnciCn25UqSE1lJbqHX6KBwQWSyGwUdVJJa0XQwGnDvFmor/pTQpxREFXW4bh0Am1Ic51O
DELLEKUXQTyQHxBlIQNcktwamAz0F4sSkmetTKh1ypRzfeqftMx9gTZwan2eMhPWgishuAQueG7S
Wyhocl6ZVJO8K3CPcEnTsyDHS7kVyHQpR5xheZ4PdnBmLMVwito9+gHry3beSJ7JG63uvdl1N4Al
VzqCacQwmu08yJ5bcK883yYiqkNFkk9Ycg3acKQP2PC1XJ9NV21Yd3FI3SDUWZhKYT9oUGv8ewiF
ZpCeBxBP/uoA6mw06i+6BwHV3Bjf6yRP639Lz9n3U2nVqHG5Bbb3Bxf3rddIRd8jYGoJ8x9PP9fb
C7cHANfSI2l0t9JSr6iqsOLFBmbdXFRewDtz/7aA4gd4AWiQFJC43LmNiU4Ql3gi6McPKVFlU8YT
IqV8qYyc3ZO7yKDdzM0suvA/3bQt7LQ65rQe7E4jIETLgcggjnw+yUy9wTkCAwvSbHyrThIFKW8S
nceVldiCwVIdMupKM9uIyweWdFZSBzi1S2PPgWygFQpBhKWCSV0UeOa77G5IZm97PuX4AgETP5MN
syn3RftFnKqWyjJspcdC3XXQHr5xiXxLR/FP1+Br/PAcCU3JWWJJRfCt8N1Ac3S3Fzpm0eX6c99s
T+UvfdB7POgbtrxn+G919M408Ufwy2H+bGaGCYk2s0zmhRws2oK28N3RFYzrNXz1nGdrnuAkMjMj
nzzj799GWHBhADegnpxGERdPr+WHSuJ6nZ8hjBVj0WLXK8fEs8dYqcj/uTA9W1Ty+RlR9vf3mkfX
eYsy/tnx4oOeCkKH9zV7LV4mPYaqARxuAEX9wsCYcSCkx0az17vjRlHGGpv1RprlAPSukJ4Cuz0u
eUJkiSWXMAz/foHOY0rYz6Ld+0x680yuxc1eC/i0el7Bqv61+kkAsqrMRNUIJzsuLZRa1gpy0bXp
e0gEFdUeT/eIcEapmMDykZo0T4ATz/wCcK/wUXUqEcli0lKT43iOZ9qw3ZjMYH1UO+nkMTCiMjRw
5Uh3RWBDk1TCST4IScrFuq+VliC1ZlkjSVcqUT1oPMm127yNPPNoSYuvSUejC1RTix2wq0AgmmuG
Lgu4lWWSD6ZdM1Fb0Lhg6ZGbsLZDssNgDgxpdKKBQtoxqZcmK5zjSIOGeGj31JckgGEiibMFvyiG
BoXhg2V5uzyN1fcb8pqXbhJEz83zbiRpK2KPdoiwciDYe1E5L8MuMW51lSAvdV4VLnN1IJpBNI3P
kYzJ5zz7mU1jIQe9qUFPht+LcrrdQ0VdNggcTiWs0UL13EkTLc/Rd2rQUV97w3ME8geeGFe5dzbt
cKO/IuU6FnjpN4SwLDnuGj1LSkcN576ouGE0SGLncjdq9ENZ7dq/PQ+0x7ZNeoUqAx3HdqHtubQe
CyLDIfbla25FXHHavJXH/9qK0+uc3fNi6fyuLgHg8R//YAemv8FpHKlbJCQ2sLQ8ixdKDionOoY/
3r3u4RbyTn6Oc7c8UmYn9yzWa855x6jH2Cj6eaxph0B0PRS+YBLUevGqfjCfa2Pon9hydpcTTsF5
ssgHBKIUphAcsCb8sZ699WSfzk6NUOxRw0o1TuCho/mq/dvKEvpF1jkYjFWFBH3GJlWk/P3+G+Xa
XoCaRROBYSYYPWI3PYG7gHto/7fCvvtSIFG2MIYFy8Q4mzo35HzfrFXly1TywL9nnrq+vekYc+Jc
G575v+R5ZfBurjK3otSQRcOuuO8SOHCVkPY442Bm35rKXJIant/9Vyayf48gbtiRrXmk8gIGybIK
ccDK5XsmsIlehA17311OsGcdtEMvWEw+CNuR/aLoGPb0L7ys34/aYYvkHAzXVLIGpcvpfw02fUkS
5RGsesSLZF+4L2AymPIhx3oVMZ0nVEUbsf5C0ukXsdgV4so9JuW0mPXmGW+49jh4IhXsX6u9dpSL
P+9vJ0ivQNjohdO/gWTSECtqMI3N+++HXVSKbKnUgTN/TBSlX6w91H5IyB+9Mk8uZg14xmCyG9pe
ifN3NC9HBbenuCg8zObPJ111C2U083GsqApQw8NFe6giGaFCzqnSh3Md2goUky3yto1nHJ34CgIh
6CxzHF+etXjx8kAgspfYqW/7k+nzU/u5EOw9iEnOKCirZiFZvGNf0lWYv42fm8yDeb+3w9SFfVWs
rrddnMgvOKXq+ycdc3OMq3hUyhO2x7lx5HCpEQAjUBEy1CDI4+ZLYStUBUXJF5HJumZWsO1ps4OC
TgzTibRZdRQCVfdEHbybU0VXpaSkX1owtdvnHtwlQwZhokdHcHYSuCMlflUL5Uj5cMstZp9nadlS
aNuLgEvm/NrmkRxMHqSd2oBbMRJwCuApeBslyFZDu9GtiB9IXh9MpFf9L7ZGqSoS1aY90+lzk30s
iSZRQaRjrIv+a6heDq57STjtlaHwbNzBGN03DoZjGSjseDD4NAxfxoQ0fbczYXhF3KM+CHMEZNAf
nrFECNgsmqv50s5fiP/MOy9SfvmvbpnTwZg6KLCkSyPi8Mxi41b2jYVkJe2BqpUZQ5p2ytFBUq0u
il34mEg/hkZherHWISsNXtyIEm5JK8GHTMB1Bkh76+A5K5ozG8bBhk1fYsgYivmzs3hvn1HLVxUA
BHvS1TmyaT8meG8XV6tFJrrfCsp2AncrRMmHkkVGMMkyzt/LCQ/XwTCXzTzbB/LoqP5x7zmjhJgW
YSSDNBKwxmJwmocFlwtSWK+LDiOvBP/U/4C+NyrI5Dd5FMiN/qm7UPI+ieqVoXepZUw464/98A+4
lMrBNFyI8tgupqyWhfA1E3+aLzjRymCfk5VSzJGRawQZuK4ujoHO5vT1WsR/VH4EzK8O8/+FLlmX
36G6vkSLTO1w/fNDDIuNLK+M18a6zkl7yMmkzYGOGYUXP7j8mcrVBz8Ye2q+gkgghkF3ORI+Uqx/
V1+u6VgTsU1EircoXG8VUIi8yqrPDObXxzPeK/rv6oGFerQXCJKRPp1ThPL+sjqzZ5Jqdl8QjlV2
QFgDZ5emSDnBuGw2GtpQa0G48mectX1LXh1Ed3O/W48Iw4LLC+kBByUG+J4bzHEDbHieB0tfFQUZ
GNzhMstqXuxInV2H1fiKT8Y5S9JXjpeWUoa2M0HkwZ1l3txsB/On/RgNIJn3hET3lgsoT8ZriVub
zSMGbmU3VtkOeTwycmtiY3QL9+/+PTJlZOsZ6NDa2OwHeCLDFdp6bU3zuMvedQFANPwYOy7DzeVG
jzhknrVW+cANZ224n748dQRgtelSDz6OxSEGUxBSRsclOzqp40gf8jtrXaIiNQfAObfesxR9YOgj
ctphuxDdB8NaIE/wyYxLCgopchNOJr0YZjRLQOkL8Ulbf9meGRi49NDiYrr5QAC+KbAVDD9MdRQC
JdfK10ERXQCvq5zW+7q03OO4dkYbY09cBs4kvTqqHNxrM165/Ib55VDKS1kET5MSv/FQfE0yPtiv
kjkCd4m3tGHhArkeXUPRaaO7b66JPVWE9E/4gk/jDpkBoso/Y1TGmbHK8BjixMH+5H/k1uIESMMI
EesQM9xS67WPpPq4neW/FIAgUp//43HF83BugiXxiXQYVlVFflWf5ZfvJBATmdFIAfW1K/8koilX
WqbVTl88tQ1Z0sMLao4y6WrieBPKHc9RGdWfm1pheKAgG8rsAtUNudzgtRbMx95ivInRnDw8OdVr
YjFgQke8ZxqB9EllRX+nguZH9dWLg4hpZKhUT3+FIgy5FdpjkyulXJFQLvGpKbeHBCJKq4j/SSHS
BJ5jw4cx3HYNi18mruGVoPwKP6n2BwCIAujtwJokSwO7pRvviCTRTzn5PmIGVf0VuN8NrGYwKe22
QiripGXPu646DmJwboQ7MiQ3HPSYhL8/n5ZfavXHcvCxeZ1+LyhwnjROzl1qD/XcxG25tWD5lOLh
E3onDMCWibhnQp6T+2Zq2QVvj7X7dsvmu1wBq30zjvhmrzjQTgslr0mvVkK47q8rFAKqFZib5ta0
v938GajeLCzLlczu9jLHgzhYnJKlW4q+jWSapvxos1im+DvkSXE20S34e+IzMUXvidM/6Ue+IHq/
svh1geF89CMrFgJhUVeIPvf5krVld1Hm+LqdwFs8HaiF3eTpK8bBLaMp1ZBnZvanqmUSCE+btl0Y
oQlDHjBbjQBfw0GNejs7cVYqOyefqbOXCTSnOV2IddqzcM9Puu9EYYabb/JKPy71jO9sGOCTMzXW
4is12EofUqQWua5AzAYia/4kn4vztW6lw0j63M7bBRhciZnNVUSAv7UyjG58zO777PKHfYnptVCv
YV3e69wLt19XHWrB9i265auFoeCt6dMsAXHbFpfm4rhK+Ece5cX3QH6kfw27MOkGG8lYQxrJNQna
GlZjyh2MzXrm8DP5xYnQyIejcJLbYSvR1HqD4NOpQs0SAVtmILT4z2LOAyEsq5cCzM03YKG/VHp3
zyh5kphucj9o8XXogFZxBlrn4tZTUShdCzAFqPuGktBlyNobqUo48kbXjGGyjMdTLAr/jwFjANXI
xQjjrMQrSDSIrwsQ3NGRropF20Jb8WorBPxrNbygVvLk2WMiK4rjxangrICH6bXMqe2ib3tFaQ1G
R58HWmY3VTMgZE/hlbTtA8OubX19BBMKSb/x6EJqhZT03orUVWxtANpPv5qsGMX/MiIgC0SOsxnc
AxppG+rTCim3Anl00oAjPHZdMMbNE5EMjIdPY6JOcJdPfBCZS8VyY2GYc5OJboPTDvblUvvyDKc4
RFGntPrDs4lYF/fLT2HoPv+vqb1XZWZSRfG8JvO2Vqjb0CwNc+EWJ8zG5tGlzSyX0Iu7HrgRWvyh
omWuyKw1t5wL+vhAE0Wx7+xYC7tuR8Lt3yAlUCF2NxLbOylETkOp6xoAdUZs0wDqxGzPvPL5qZ8D
Onazq3xwqJRo501J4xrkgWlB+rs5F/goHUs4zxKGpLBh3z7bfGTYd92mU5cD0w4Iy8hi7QWx1uVV
ZYHPQNLupbVd4TrVzNxP/VBm+F3mV4BAzhGFQHqaJMM1EjcLTkzEuXcH9wcDABpfJB+JNOyZParH
bZ2xgcZKpjVPnra5U3PwLKv29zvl/cdsjOnaZ50pv8cqEUSTKIsC/V+bK76Lu0EI5W6Y8ZhA0nf7
amYMJIFGGT+wRoQa5bkFgJJECv4NvyXOH95nXejYeWXJu7JjTOvKQMdUDCe4j+w/JC3cjuzr4x0j
B+hWb2qQmmXu4c+C5JTUzuNgpk5alFpBR3hzMJCHfp9xoxvmMe+HNOs0hp6qDhoJ1ClmzzTrTwAO
ZFIqfOJT40f2KKaWc6crV2PHjIkdTLnWYAsE59S88Y6D/nxgcf6eIrwGeHazGqSmdWr4ZXSxG4FT
SFVsHDZ/hj31JpS9KxjUuBPY1sC6ZvPJt0hVY28i8EqWTUbhhG18s13z2aCt9ZAEjFbcUMIhWPfm
9hZDaPv2Gfd8oh48fAA4ke7qCTpNI81NRqBaZnJIMjB/89qgK29cYCVgHfmiNiDeE2lphDfy3Qdk
XhbeQTOqMRiMmPwAUoxnZqQc72V4/GueNYop8XAhd9Qz3jfqLhp+yieu72lOOfahWiIzlRuXG4G3
FejgqiWJk26cV50nUfQjS+fvIJWjTATwy85Nf1rB9K4SyFf31XI+FBx4/bFk9K2xh8E/1bcfgugV
ZbGuAPBDXfncTBp7t+HN6ujH14Pb9JNJ6QR7Qs/lMImvuewZ+YgnUa7GpFPOeh5PSRfD/ci8otDu
V5uKHH2f8ZZWGDkQlas1jOqAlkTv5YxbO+qqqQSArybQ6a114xVMUJkiXaK/8T9JCd5X3SHZyyc+
WxEv/qNg6SbSUq9T1lDPfk9HBDgn9AfpgkPvp4PibI6EUp2qxHspzk+d1wPpzZqhwlBqS0TcMgjF
q2TOYe/V3z5YPwvXZ0W4mX+T/y4M+REQb+pj/eMcxqP0sXXFDug/MgvPNT1Vor++9FVjudF1hs7D
BlJqSUr8vuflleRTJvAquSR/mPsmOy+/xPamGeuE1V0UnVHwIse6HDQfLIwy/Hjq8/VRCLPKVQWF
8gfEOjmwH0OSskO7WiMnZo6bwLIMXvEl0sT5QB5pY5srrnZvelC3BubWHj2M0znvsD/d1qTJGemf
w2+oSP01Jrk/o8i/ALI+AeFlrIhUEasdR8yWnVNjsuOgTujbKJ84DM8SkNcIfkjSPlewVz25iQS4
72i+sVmeyEIDutIodgYCliBfy0Quxlcs9Z1AORj+sk60lI0k0IkXVm/zo5bDlepXsSx0IfM+jIjj
SDwmfjtbhKHYFRkTWzxqCJ+6h53TP8HJiQM3/aBA2XehuybeisL6JMECLaLJoNLDeheCjiKKdjMd
AaW1AB4rDHQ/Kk+SZEmTyD8uhfKIx8VQO0bHVPyUNZJcWRIE1tSgqbXArRLwGRAgX7HvloXZyoOE
CkD0jceO5KW90Lkt7XTlq6ugapjpAV3uO0q41NjSGa95ead90eIQRQyRUFa84xpHutSvm/FL3Mzs
F0/Bv492zB30dI/p8GF5jj0aIl6fx3F7tlseLbWeud9Kja+P8ajo71/3VW3S7XhUYVvBpzhgxEyt
Mx03lvms8iQnXBjc5sivaLxFTun6exS0nT9Kw2F3cW/6WnECBpPyxyriAIHPCAC5uQBib3nBFWyT
Kz8p/3l10lcppWhbOCfP+M5FSK0UvIE9sM5v9M/B98o+oyhM26RLMubGEE+c7etwuv+jJx5wb36f
Q69sAFyRy+8n/RLyfMfMdyq5GiMFMcYLrvIT3mk6vCQ+wVMOB8IHEuovr5Nj912NacZHWsTxABd/
1XVcl32X1OqIynilHXxn0stNTk/JSNgDdKO3Ew/a/3nPOY/3yxeUrx6sH2ZylcNEXx/gd72BsM6b
q6d70prb5LUosU5ZCANXuLWMzi1831S9yzf2H+b0vB87eaLbZ/IKpwpcNDrjNgvz1/00m3zQxy2a
9WfEWvyHrrG/c/OiKpz9UwtX/xBnmVhtRuxzf5r3Sj+pfZfpwJ5Lkr6Spgfqjm7cFcxqFpyuEBy5
pALj54JE17ZmTOZpo/EV8h99cS3tstmlK2kFYtCD28BZ/RvyOwSv7ZwiNkDAOan4ILkNjaFO4nNE
+c1H7rs1aD8y+KNcIo3Q7+fiaYFXAG880JA9+Kb+GzOBoB+xgKU/01EFpqRAeloNJrmfpXxysCog
0DUIQkVf3JZ52TdRy9m2sQDuv3i11oH5bazCCyScOIOECnayEL5tHk4vhfwnm9mZv0SZyZ/tssZy
gF5D89dthPL8S12fVGwpCPLNkNX9kj4y8rSFlCvfjkIZ6+6+8qlFkXnztc+S253BOKV4Pu7Tu63E
yKxrMpnuWCdqj2XmzQP6kKU0MuLsWgqUHUQAgRNYMzmhFXwy9SBFTZaOqzf5sOTzVyGC3/J5F0US
pOGX9wfkQmLPj/g0wx+lu17j8rYHzj5aLCzujIaugm6Vc/0PMCBjEqfQf21RTlrrYlfJCb0PuT/A
YrPkRV2+8CmEcn4KRx33cC6TzfWIG0nxJ2NVnz4Ssm8IqkVtFM1z1WW7S/N0apNQd3TdPsUaqxn1
8lBefdGO9Z4nNjc8IvHAb/TwQkQwKws4xKqaaGWiOdV7Uog7pidbQNynn5FQP6VXmcztlyBbX6tv
D+RLcCpogq9SUVjS+YWAP39AaLsQ/oOYIGxvrWJIF0fjRwhGGBdltnwhYo9NDkV0Gk6GkPFIv2OX
gpYqpMk6FDtPHHzifWS+1K33h9RJvhDSplL11QJl9WDTeAnD1QgpKq1ORhs/69BGK/PktISd5oK8
TgR6v7iOd9o5jB2aQca3Mf2m+wrtw55mrS/T03rNExnuVzRseslxFpulNGVWBdXz4WtWbOXvLaqC
BWCivu3j2fz4+dEdIiSAuQlXv1nVOSEHwb//zHfl/0QLsG+naauOnURD2DEe+jBFXmJlP4hklT5A
7xI1DiCA8Z4LBZEO9sbzNUvLj547bQrcNP0RCRIqGR4NrJdVJ/ha4Cb/H1yEgL+POQGE1UW36rJz
w1cQQj3kyJszCirzJZ61bEc5AnBrrxdQQlVmEhFaVAqIl6huaOzGjBbNDhfVJYt8hDKwvcFQTOEA
uT3MhsQG9U44PU5FhTQGXYwLceu8rL3Oz/QxidlrpZDL4Q0RLllt/bu65GpKED1sKj5YdS5O7VT/
Jb287JXpo3V3Z9N4DhSoDJqbuRUwjw6ClGj5hXqrX2lNCbSg+2ij8yRPc02yYfGRemAez1OwidvK
RyjcQfFNn6kaFIn/lssVfRJqpltJVxy7VObuLrWYOB6ithzMdNTkqqVhMhkfTYMk/1Y/Y7IY4KeJ
LLhRHcq11XvMX0m+2V82lO1SgzjSzVGo7rX6VAFSr7ZV/O73HMvOz5zLkhnsy48+c/2YnXeiWhZX
d1y3GjvSQrv1deus78wvDfryNb0W77wqpF3rHof4oSHQLSIVPZwrJ7rS1cW9ChrqBNWDB+3kDUTh
vCQeURRoDh77/pothfb6G+QKcrQojxpbigqSy1haHx1JrtzkY7Ym2uSN0Rul2FVYaisbat34Rs2L
dL/hE7xWviJwybnB4JG0gIlQ0dTDgwS5NF7NFjX7Sy5Oni614vKb35Viy6hXR31gOB1QeWOrKcuQ
2e5iWnIddNw1qef/O9Ab8qMZiDG4YxoX+hi+AUYO8NTxsZ1gYg4vhyRELXlfK1cIRMNx/bknK/st
B8WnoHGhRNPLi1piVy28t6apwXd3JuvxZ+eQ0YNwlQnfgj8oKJIvtC7faZvurlGueF02C0gQzPDY
isKBZS7LY9Q16Oo5z/ipwDGViFfiCevZIG0ap6X3U09OosO5TA8S/hpTUA35r5qmY9Rr9rNFIuMq
6siLCwcKJ68fvv46FWup1bOEeGSkqeHEzmzic5iQlSYWmsKUzins9ckdAkuKlXdddQ4PpgBtGfsO
zBOe1U7c4w4gHn9xnnceSpR+VEQKklX7obmmWKm9BvSiZ1zrrm3TAZ/SRhMAVSFdlJnLdg6CjHxe
BL95KfCQ+owjKmapKriWKFCRHuH9LbPFSLQWhd1/g2BoryOPTFebVfiGflM2ANw1+qYlzrPIiKSC
1KSMttKbKh36pppdluTibIGlsgJ1JpHHUB/BGbCzn6hM6oFmutpty3w7+SG6OnBKGGqNVovXrCTb
AeqPEOru9FTvOh7lhLH5pOKPq99PIFK4auiFKpeLRLU8tWp5DqiGf1kCViwjRW87bK+MNSTOOWlb
xGBa0FGUPYzGF/qlxaObK9HifaiipEIrk1uBblCGd1bFPSaUKnRfmvZwFez57SME9Hf88sGAJr2y
kdRNS1bDSBCGIVzvBxX36rq6UluMK02//QZj31FiFgJtQYC/zysTTRYaRjbw03Mq0bFsBT8jHqat
dKCo57RKlvBT1Awxj3b3mZ1QhxvCbbfv7LDvVLLRUJkZdmJWUmgmkg3DLdMRC6YUJ9W1qLowgavG
pZNd1uvINZ++VnnUAnB/nvuR41bemRVu78mFdo7XwOBy14fVFfFXHzjq/TblFehtqwVkI2XYKdzg
lvpSJu0DJl/pg7pwUmiKet/yRNe4rvnEnYINx1VP/YXom2KCe6gYlNOexeuZBcaQ1O7qY5o6QQCE
kNKqqnzfttKVC1ey1DFKvo0AuQ7/tmyNPLImNqzzivtrhVZCkgGVmdybI3qhMNrhmMB8eGIb9TDt
aeovsP78sEFIN8ObuOO5e0LV21FxBagwbWGZI76TRYc2yDrLuvr1F+4jR0PaRy7aDQJkuw57nYW+
w7CKRhrVkKx07wGcTfxNSC5A7dVNAEs0XrB//L3n+XIM/vTV51e+Hcdr/RRbwam9Iwq6i7atxvWd
skY+QAxqQXXnoIcpfWcKAagxdg18ibNDqcJXDf05QFXrKsuW0wz8Hiq/9eYB2jiactIchnNdmrq/
MfuO7GJ9U5LJQUctOUVW3Okh1fbi1Y7OclqXSrj0Se1Zf6QuGmAq98CF9oVUfgYeCCiV09kRxco1
NfpFve562jkmEwrjs39koEjDDVoH+zasqk2MhiG29nG2Tyio2TVN+8FUMm361sCTVRRp0V67V0r6
cV2C1Hbx4l6EuCTE5i8YStGSadvT+9qckj65OXiX86AzLUdEdBdBKFCLrqzZzG/P6UuDoFJsGUG3
kIOyfHRYN0sLZfJzdgL+KrLwWK+mZz7vOvEJZ4H4PQtUUxta68nRA3tG/eMMyS1GlikHzIOOxcWd
Td3G75STyIaV0kGaYzOvwRnLQEq3co0Os+erjC+bki1jsmBVHcYifjRY44d40o4ecO5daZ9iZgqE
9AEfctGPvcYu0bcQAMMAv9y6mJnTfA5gwvw7ZuCWzcUx8YDM5brNBbHR2pgJZ2zICF3PsXNY4J5O
B6uiVdxj+ZLTk1BMNPJR6KBICvtPWWt85GYb61VkItv+axYLAmYezco3YYzML9N0twewFf9XDf7c
WOK+8zIxuGZySFhPMGSV9dl4ajZCb+UU5pWZOwq/54LkjJhWlz8KgQqRWeEj4XsWUx1HcjS0g7B1
R+GDIFpZRgIzjfS/KaUtCUvepsRPdp84Se/MGRE+fP4cpo1u6EoNRyaDU7gMvzZtlXX/w0oIXaF2
534FZKXYjlgxOZYzSiU58Ml7hyXdzhw1f3j5EZJnFpQ8f/qupLPNZRb8WrlW0nB2ifsxVLDREzF9
+SzH1jwK29tpD+0r8l42G/SxvAOJGuYWp5+OAV0ShWiza4GPbMJbmZ93sWG0frWRw48VOfwtj11d
RW2YLxJwaVKtda97ITPkgIoN9iYyz7iudeV8/y9YNUkrKnT4soJXKkHLm805RkxwaiNdIMfkHUVq
24s0H6RwwE9Pllmur3L95RNLxea3ZmtQ7uRywBkeur/oE/beRAhfmTB1OANe88cJ4Pg34H8T04Pv
x2j7rD4vsbkxmS9NKcJLZvomIDVQ692AFNNn/USuu1HJVMmf7sUnaUr7siExaJiCRVs+2rnlrR6I
K9GMolLcA9C4ZdKVBsnk7Im3+xLYdYeWUeafu/5eX6q4ugun87TkyjzrezcNNO11oT5HYKOu41Jr
rU53KcVe4nD3LEt6hHgCuC48WYFuArcAs4oklMXN8ilx5lCseqAQLtTOqtTKTbOTSpAZZNeM7+TL
TuM9F/XS//L1jXAkttX1XuVo6OrrFxZCkxIb3prP7IjdsDsD3OY30SY15D8JE7Zx4WpZDKr9MEJf
rnZUKWXPcfd+t7YrJ0WQl1L3DCqMn51YaueYEfKUUfSNp0y/I3hD43aqaJAwjMTTaJQWe7XCS7nX
8DZLXGwjgXwhZCVMIjSlqOUYk5ATloR8f7FL26TrT56pwizy6wp6jD4zA3FuOcgE9Z2i18NNwKqt
ci9XuVwUr/5VEvoKCWfkapzoj2191MhSN4+qm2T1GMGQYpLbIkfIA+bV3Z6DZmYyXRLF6q6vZ11R
f9gdRzulXQvXbp79FQVv6/QT6inPDK0i8KN5E73f5AnUxW8z/0e9BlK8oqaMYDRv2bBEM6zMVBDy
9OFNukMq2GE6ng7kMxJN5Vi+moQWIRnvT257PlwWUZng27jzfBNJcCo6MMjSIAintWBNHoFxPbey
jLEdUxSU0KMe9jSh+LeELSsBj9blSKejAHJYMSHUXaCrryIqHTM1t20o6/Ny/lta6ITkZZ1GiPqv
UoDStQphZvBJ1Vqigo8UYt5uVMtK1qEHhUecRo3OK/mgOeJ+Fy8t8ArEkLmJK8Hm++oekMcUgaGJ
D+X+nNrKz7C15DvCb8nXsJDA1EE37oHuRiRj/vWUUO/L0jcJg7HnnuZpPT86Yse1RNb6iEL4n4He
5LmHxFFmOmj2uaFXAOSMXsuK8AaeptvN8K2MZSpKvmfWB0ZRCTjY+zW36wiKt02IVFz2rzrL2bP9
Su8vjuHcVX/KY/kPasSl0q7rt5/p1BBR5iG1GshuepHZ03Hbe5ah4MguenbEIEWqC7HShmEZvyLj
IHMZ9tJetNep53xOVkyUaT2vSZbx9S7jaaORzWserAeqBm2IipVufkukty+o7DsZabp2HHIZId1X
UiDXYuaoorR5cXuxvbniVd0J31P/Uy+GrZsvot4F62oTR3/6F4bZR4IU4I+Mi/AKzAGcUDjj46qa
jgVXJfywm88OQlUsqVfvasUejbBEpr0WCvT3OBv/V1qKJrXFpO918yqw1JpQBpFn/MymMMp4BbkV
bYYBAJHde1NolzYxpS+GstIyX5rrgHlx+OHyz6MWGQAUPj5cf8YtxWepz4nMwQl1k0x5Ymwp1nJ/
IsGCvUGUgF9CEOamBa0EbClrwnTnwSN13Tey1hpSGhRAk+2Y8TyFnfvh1lASiCH8MzuK7dKkBext
MRkwv+Df3HRAIe/Es3B8YVSvqxengSEjQxXFETpga/fWTjLHNKBk3Z6JJM6ghKfKu2Z7krd/deWr
pwRAJSuBPrvKWMmfWPZbcNMLuFlgzEKs1P0p3LFLhppUt+MXdroPJJNRo/c+s1SAmZXT2Av/B39c
E2pkwM7axPydH5S6qS2E8+THmZBx06j8zKSOJdWbjRYEuhmUPKWkNF5+YIf/fcOJJIO9aZs8i5c/
xEjuelBOJi6dF0PXxShmXMdYFThhbCpmEPoEF7XkQEysNgOmeJ9Gtw7UUzm2kFWr+73D8RIS5jkd
0UbukUr7MXJ8DGRWgMluDix7Fj5OOv92HFjiA4Ofe5AZhXRwQHJFdbtXhhVPFb/oxVrSoYl1Fr5w
UXSmx63ohCeZVwhLMUmcnBVEKLaP4F6RuWJKorRHU4aSqe51ANkXheVF2DkG0WhBYqDuDQ1vNUuJ
xSirg4+2k16mqlwhDzE/pCAmkRIuRfak7Pifoc9tr1xtpRziroCYmMPzTLPYGVz2qz3hBir9rbTO
+LEpZuXH4rw/mX2J/CaAQHbpKBdMuDCKKtuU1DcQCQnro+fVNiq9Z0QB3WzVBZJQv2OdrNFEED7V
1MXABrHyTjzn0ppg+J8l9W4Syzz1WkJv1KPwN/OAFo3oKI7kcAyTFtvXqdg4yGZh9Jx0vilgH1YZ
ajup98JsxFEyg7Qt6Frlv2GFaty9Wzj28FE2D+tC3E9FQw7Dbl6Wo4DpUfE4hVRgYwtGfEbQm1p/
WEljE5Vvj5ppZ54Y5xDsgFYLESvBNgqGHmmlExeMOMXhLEzrHMsSLlBaqm5dOQbUUrwJYy4Jdu/c
VXSfiJoWvLzprnv5RTkboWobdSoDykc0hOP2gx8BOadxluLb0a6JBo9KH/NShQe9B+GC7iGwTevW
A7G6Ja1QV4G5BLR1KZtpYQsp68S9IE1rOuCbUwfpMJL321KglqnbceMYiVbV54N81JN79CIiGGU+
yfzA9vGOY4uRq0gMqnn03fbkBcXBNw/aGFpQDfXvpux40xmKUB9vj+rVOKO9OYrX5GBIEsS5Q99Y
3nsuwnkIbTAxbgLjVW5NMTgz99aPE2FG42N35tOn6XLGPld2+3zTrwX46vq2hCDgPXIkYwmrVVti
Q3DUsKIBUSIZXey8ncwiWZNQfZUFewfNQsMKTxY775OUFK7boVcK6FO31Qn19VykF+vhPEQezfOA
CIoYszyA5Ih+g/NggRCZxws3y162XV9PG1eJnemIOgI8Angwj1/CfG6xBQ60dxz/vXBYln1gLSFK
giwnF56skRKuIVED/yH2NnSug9qt/v+K02b1ULgnUIaSWXhd+vVC2lw2eq5V5VkuWHmNPC/abEjG
h85xyQh5cZa4l+QpHPhzHvlOJnWap0/6xe39c2KV9uk3C0ivaXMOh7CJo+bJfjJMYylPgMpwSWlv
FUmg8MXKwKs0v/O493cBVuO5P6l5soeCo2nRPeHd8JX9gsaDFyByK/fGUjq3WnvmipN7Nylax0Pv
6o0p6p78Gtaomvf3vCYGeBCcHzzOhTctBO9Rt6dNtEqmDuJuZ9XZbHq245rRDB0PLcg15nro4nDd
qVLFFpDbskAo7plZ6SjBTp0+Asds+gEzrndsKd/+eiL8GpHy0llIrk1tmQ7WybfKD+p/v7hkF0LH
5vg25GWPmqWZgTbmC67BfTV7++ylpm6icJK9Y5g9qq+vp6yf5QM9YpTRDxpmw1pNrvP1/qcSjFXw
mIRR0SsWYF1ta3qzJ6rNNXbNW+Ug6SZCfrzZO2pfB+djhUfJRNoT2mrdS+JzSN/gDjhY14obX3XK
8eMVNRAnVS/BbazjiVu2X5y/VhP9btuSDpheqRs01avBBt/g0x3eXJnkYA0Ohh7gPkmd6IlB7s1C
s+TUEGJuMAYb0o5zPXLFIovHUzA9Bfo/rvvR3+o14m7+FEhOZKRqJOFXuB8wksuVtI8hxovWseyu
bZ7lKESEqScibA/f5UHpy9jBqbTEociRxQNdI6PldMPsM1ZOQFHGW1HnCfeJjOdVvsWFkOSgRLrz
QLA5x2SNJ5VBBAfEYv8CFWlBu5+a9ZDj7COYfKi9d066beKoyxD57j5EUwqLb9Rg8icXQRCQpzrL
toflpBr1URMYRrsNAG8GnHP8pq9TF4mwQNvy2p+rjX5a1PEDWrh6guWhXM5NHy8JKNCP1ppb/zGh
hEITywhaXdVVYGq0dIs4AxcBx4fqPYl8Q9sKT+evRQ0r8W+9++1wYaXp6lId1pM1VSJLCjWRzsoZ
wUCjtn4C4kPQQjM5oNb5xnjLubTohQSAMX/EsAv/gM6Zldr/S4k9wBO9dUTjIq/P0WjXapHvNiDJ
5uvN4WK8viW49JDVgJCk6TX2r8YzB3tXi+tNc9oVTUDCQ9ZpJNdm/JMMj5ACjnSpunxXs/0a0GgG
dct3NAytmKWSYj2WE8CMaZh1v2YiX36zDn0sdHGW1XJ/yqYBSTPFVg8f3jeqd/Y39JAeg++2E1Lt
dfLzCoCK9z19nCY8f92HSdX37WczUYG0R+rFdJy8mu++RfmLzHrvm9+lNAmdSto1Phs0iKdE2nJV
I5DFv5zLl+VG9CMNdMCl0LUynd7tYwtM7cfg0X6mV5PXcjdepB0/eqITZ8mJvZZqGBMQWHa2HWUM
kZ/4bNB+uPn/t7Bl0dIXKCpKXF+qlM+7gn54yt68B1DoUQMM59REO6tpvMUPjgn6/0C9vVk057to
jxNoPqwvoo2HlUE8Tmjnvn3IYSR1agB1uSeCtvrz0j83c06xXTXrN+ixnc4J7zpgmwtIs9rumGHg
mtWdYV1k7U+tzM6M9c46022K4xwb7qPLEtcoPxo4ydeaeaSd+N/oUiGlQ8n2yvQhAxnTHR+Apigf
WjG6YJSQPyHAYV01TL/TmrMsYlJJTQg8UfYU20parpYKKU0wm3s0+Dhv01d3d+NcPyOscX1/G+bD
QmGecV5HDuACYqjvDKsWiERkkf7Fj60mCuWjVni6AwsjX57xJs3frL6Y+W2Ec6WeEbJ4SxiVPpP0
xDDrOJm/Ld2ysIaV7XUybt76XoclBvx120zhmFYUWCpg62QjDEDTetl7HsrrHm0qFse1d3K9jzTb
gWxmCmER4Gya1l/oSY1v8CgbWxIWstNrdOxMY18QzZA95KABzHTjzDsXdk0YNntiFYTNxAbtxQiX
7gFJ9LsTzRmIAtnqtrkxgOKTOFI++1tIVkX284zNFQurb//f1tNxEjbjK8iqyCNUefwVNFI6wskO
UJaoELPwCR5/OIzz2A6fR+pGOSQFA0V6hMmikzhMr0pRM/9ZXzTcZ6IgGHAPoucFEfhMoTQAgZes
R6/247JnkEjiOUtH//ehIgrb5QTaVQpGl7ZfmIbqvcUXoo4XeZqa0a99sc2H3ILki+Flnt5kY7hG
nBorPuAfq3+pxa7etP2ic+q+GouVdMRhfQ5E6EGU7vGU6+ItGF+OimLWSGya5xDWQjh/FWawdASG
Em7Px7ccEZKfI/xgzf5qo+qV8LZ5tR1XEVkhXLWjyOJz0HKESHruCA3E8NSe6HF/G5hZ8wfWJrUm
5qMAF0ZJgUu1bjZJ0hkPVDfDBf8fprC2+6QZBVZHtzZxOlitOEfLlpKZf1TqSa9ON+cz747e3enP
/0UsaadmKydXvZ48oxFinPvYKap+qZ/eGxB2aQmptvBiz/W6K9T856shooLHu2ENFS2CFbO2n+1w
IMv/4HdthfbUseEubGAELg6WABMBID0Z05KM8X7KzuL3dKkfe2xgO2jinOKbjB+Ti+QsyyP+Rc1f
DrWxYmG273WF1M1cDAdIs7IXpYFqiTncB5ebmfrl2sAJf5SUhcwj+ObCossXCCGtI0Mbf2863Jai
D3/GlbIerFtX8anRNDW5xgKIzkZV+hlm4rDASSGBeeiu/9CtxIkKdAWIGDdG0w9LPFWMofUaswLl
S5ZTMYAW+GYPVPHdnMjP0bgJq5c406IHx+cINdVz7iiDzEhdfY/WNjGuqmUKhBg+HOs+soA6dhqU
yajZc9mu5wbr0/9uJ1z6b+oR5cgI8/cz3f09a3XoaWMPwN72VB3YysNizjG5ZTEMUY70lI1M820D
FA2+/0Vybmhl5/xZJAn19+s58Pgtmlcj4GSTPrRzVMJqqU2VgtzhELiTvUlWO/rX3NBjeKOGsk7P
i+tOKx2wc6ALkPvxTgbZ5ldtOTjj2x+rlXaryLzTLousULKrW/l2SnLl0Oh2VJk+kLqiFotzD6wc
pM3vABZ0Ja5NliC20DDF/Ev9k4MyPsyM61lPDCmc3MhCqsgtsk6Xba9DZaSnFeqJ0N6UReObPVdJ
bJQKMZSwoGVem0MZnqjnxHRU3+V/v5LUZbuycVFlWPJAeN0NUlSff9314cgkS/rz49J4tzyxjqBv
CTbiywfFd+vAbPw5G1DtSNhpxFXsfFPcU2B7Kpf6Zkz67mpUNSUhpO0Etv4GjRk47HXvKH8f6VnX
j+1mwNPW/RVg3nG6UqLeeOAIKXQyetRfzeoMa3k3XuurGh78SJjGEDK3NjsHOm0LNAtbhS+BsGAa
/gUsdq76Ehc/s+wJdlXYRo+EchwuyEGFFzD9gvlfqYa9XkqvQpnG7mwhqsd+zpfnWuuousjpG7hx
08R3wXJPjvYJ6AyKWPOVb9Y7+ZCLSa7agF2xai1qSRLQGySKWlSp5H+6qiL67/s/oEiZI6bjuqSS
1DVm7MP/yxd062BdOe+Szb0kvFCaNlaU3c00S4GiNwH7Uo6FbSuejJOdRudbIdWTMHQU110biwD6
FNMfu7JRJ0QX9egEY0jMHbOp1uaG6AYXmTpq1f09ytCuwXZ/ygq9oQeFoeyIehHJ3c25OaxLzAqF
AKFpoYsSLxk2tFBbQxNxq2GAOwSMti4CCfwy/pmLIWHa77CiVH7oUQLTBFxrMRS+fDwBKqcv19Ka
WcwoTW1Nez6WcQhTpL++I4iPSLg1NLI07Abe5a1Uu/03xQvC429tE1hEdK0aYjGMs/3F6cYXOO2y
f89cdOHK+2g0qCtvNRbC8WPRIUF/oBrF4nrC/dsFceGslhWfK4mmW32WbIoxu6QZ+kOlnwfooded
SytmP1ej5OttxxNgtpYm2gwBxXuUQwhDSdzN5X0qIH/AG9MkF9B8MkPRczZZHgZ9LmOhZRXtoT7j
xYxpIsEPoofr5pZrWZJonvT/d2wCb2g57iDzMyVfn8FkyDsuTrWKkgqhBCr2LK0prVEDM/GSRWy1
pO6we77fbnBupmhtL1NNh6iF9fKHuo/ecNaoF8asCk7ZWoAX1b+mwFSyt4rgIwKur5CkKpLTaUbo
BHqQngX8GTmUWNms3KUtgjges6NZgwG8+W6ni09rU0owtbn7iujhE8Wnyjp88s9op1Mr78v45NVa
tOveLFFdiKnHPBnkGfhx54MLc8FT1VREqykwgopXlz43/sqoS9fdtRebRckKLh2R/bh8iOaaManf
HkHijjchtzgPYcBSJ7ND0BhLqm+368Fgs1Oemh+P1y+5xWNIqyk+lSKP7I8xHXBCI8Lx2QXTvemw
iZBnHa8CyNhxphjwYU2qf/MTqWw55PaEaK88KPAv17YfOA2yL6y4azc33OXQLTWCHoH0VanganBm
BtX2Bcw+nn/eE6C7b5aXR7yuanvfBZ/Y+HxcjHEHssNfj/uO2K1AvTvdWneHzih8bozvxW++XyYv
UNVlb1V1FfBKywJ7nKCyTlHT9N1TJpAL+mYo1+N6ILPawi6Mx5UwYVoVUAWo1xU16IK0fHxRSTfj
gAJ5cMk17OAkfWA4p+6sfgmPy3OaZck3G6MB6Zj6pHwjU7+CqP6jfPcIvvNR7qU0iE0H4Tj8hDM4
KQL7uRG/y0/mGI5vnt8IKjPzYDgQhZTHisqEr+4HN22l9chV8jUZ09Ky2MVBk20GuVI38AIV+PS1
SIDvEA4IAi2NsUZZpNjpPbMnTTGvi457r5y2xOSrFdTK1UFFXjMmA0sY55R2hF+h9/9Afe8PLDsE
iOTdWRAg83QMsSrD4zQUky3K7kHG8+2BQ9iCfyh3nX9fvch7YIBvwOZroycbwI8foksM9Tv2nFMN
8fzAQuhQPL3a37/Ks4nbQFgrwXMQEPPRCUMh/4cE3aEks18or9L4+YMkoWgbThRl1qauqUqZyC9s
BxbOzY+gtTNo/uB09JVfypp3UDadlH5+v+URjzs+HejegY9E3+aliMIR6+GWZ/RYxuvA+Cp5PSrm
C+suhef/ci/TftSes6TF/LPlhEzt8cW1diuoucLwZCP6wxHSQkj60jBY8l/JOCUcNp8eJ+/jcQfd
d6PJC7PDvO/AbOa9Z/qRiWWcEbyNLZbs+iIF+v7pSzeeUk21TI+mr+ZSrUUnF2ufM1dyTgjksOic
JaQ6LHC26EEi4sOZvCvX3K5AwPRKtfEFGMqPMy4OceFAtYO1TgmHMjY3/Mb0hl73S2HAfqqrLDQX
NXylhy0bY8kK5SVfH+hfxj3VZIw1qmOQN/XWJTJAumr92u3/YSAWb1vcD1Em3zb/ft1runDR1CXw
yWm8nv0/h600rdbAgIQJtS2AYaNBpIYcwPp8DehsgcCi5hbJ1pOvz3hZStfC/RW9q7naTFOsxzhQ
50KVKUuHG1b14zPrdHgN+lRL7hG2lnvqZgr0hDAmMZh4d6csMqVyUO+VAFU/ltRROSU0HqmQzsk0
/0ZAP9EPvwzG8yG+UiDdvOngCeV7cVbrmwb3tHfayu9bC/JPVsg211WUODvGN7vl+c0AnO05f2dF
r8jcNWaVcELLif/W5UF+7gRNluITVu4M8fKbZvR3TthQzEMKizAxSJVefVsVlXTvFUIuBWxGj8CR
4gsB8fAaG7MMGE7fy5xOKRdzQ6XQ61JAUrLIpqDe3+Rls33WgsPaUqCRqnps/KDpV6cfX+xZZiAP
blgD5GXmCA6VftmRm73UQO3mqevMWwok6saAUdPMwTlH1MlYtWyoAL7KbEHE+aawj4TDUhlruPcc
RQwoft5YvuwB7IRAF2sOVS9jQ8XSUuMpk3wkuEMBhloGOuTRTPbdGSueB5Q4ukBLCNfphof7QyS3
2MlxbJ/INMXyeAaxOh/JF4/XpVMBdWkKd/B6DxS7fIxm3iWC7ElgntjGbBAUpO30Rn/6Jo6jlfQO
RwWxGFX8jxm6knODAu1iERkCY144YuF3yCumiyyWpCt7t+cgkxgMiEB9+WRNficx6qP3z/+6LQql
4vM1AlEk+yLd/nfYOzI2HOXtQwOl6b3ck73h0K39RfRdZwvZ3/SeGFNnB9T6jAoz99HFMeiFPn6v
sl+WT7VuU1P7L62wc6dQS4C65BSdPXSjFJQ2hJXHKaeztAldViqcYqGXphfJrgqGEHVVuVn8nnzC
cV/+j9k1waR80TT+nlKH9I0Cf/WN23yIP9xleUoRujmL1T8vMGZ7QAvLqZzr9C9ZdThUzjeFOgcE
2B+JFz7gXpz1cvIttXQWeM+4JltFB4vk4GNevTt6SwO+SmR/xs0Pf5oN9l1BH7/wtAjzoIhaatpT
igWFF96sXbBv//Eiqe7uunFHKPl1MKzo11GM2qceV/L3QdCxcAViaw8EoPZZyTzL8YFxuyKgwwtD
yDmDv3HE4JjAXADZXBdQa2qf0dA1XDpwuPTt7iTWIjYuHZ1n64sOH/MHSsTCeW405xV1Qq9WkF+u
1FIwvOSvUhMH6iVIUOBou4ec/EgoAYUlRKUayv1C6UiLJuTPNSmoCvuhBE/WGcjb/yIALT/6FIMk
g3EyPuhvHwpuPH0uVR/zXNPBDhVO8d9w23NjVVbaIupeTUhW9om4LZdpruYiW657MOMo5IId2/y3
T+SBaXVWbBIQu9c2nyR/MWGHUKvVwaPulcSY3GzHX6DkRI4nl5AvAo2nuUZ0ieasvQQUeK4poXBn
lL8NVj19KiLBEv4eOX37D1eB6JV2Vb2dj3HUZK3F470A97O9xQQ4iW/IBKwiDNlYMDE+d2i3M3fN
w/iCIxxZx6idH/A3jBd1WZl0C3FzKVtzt9vBa8Np1LUvRUdAn0S0pmylPuElCNWzgRsLzgcy1YY9
Q6CFsvhFM8CuU4HVMg6QSNDICyZp14EzBQHsQkkJnTwQwrxR3KIAx5hMTCJCsfRfEIOLQx+3CCTe
rit903fE67Fzd2/9BtydXP4hPHa/9Rh8riT8oeF3sXweonVMUrLn+sjTrm6PKchfkHIQu6AJ4h1m
MJohIjfrskFML/xgZpjqUPa+wkF1TPR+7MJFeqix5XuQl95X1NAkZBnyvSdt1wxSKkoan2TGvfv6
+XO7HC+4AXvVWjMs0sBu1pP68p+VfqQw1jWcm49Hdq38xeIUobBYB223QT2MiLGoKpUi8CjxRX4b
b7l4kOtALxOwOuwi4Ua4ejOoFYA96ymlNYu5xcK4HMB9ZXln3n2Z226sudB11eESKOyejaS8VRef
CC11vvTP2DZTfPmQEIt7L0E262WI3jkQX1cG/CcCZY9jiXY531LahvG94GGywLJNyq51puWXGruM
4mMRIBN0TXbf637kYc7c1oVGU3YDUwCNGadPKSgRVy998ONdoscUbAHpsP/CKV3xpbgD9W0W/Bqo
9QOk692fwUumJCSVutoGCqKxXVwlUgc+r14wX816AshH0o/RvRLf5IuPSBIQuknljJkYA4WL0QfO
asmdENTO6D0q/4nutYyXUdhCx03ggx65rRkYrQfin+BDQsFBJtk8S7Y1bSVAsF3HN77OP7FDyV6u
XD6/quSY5KJ/laVHUzf8cUGNHCzurLeYGwmn8QlGrm5rWcYEi/Z3bNBfQZFEKIsSKj+HYNH4LAgg
gLPQMElBZ2LbWFkBnFo8DUQ4cuGLXgJ8n1wqc3LWxIk1xN636PNh5Eusp4ycov3nj816wV1TNh91
Hr6+0aqI+NHGRUJdNDzNKsoziZ1pQCZqICnWXkmLCOzTv59Ey6jZPJDe7D6GBN1ncSl8yz+bOmfz
8uk13LKL0o9iBmpZ5H3B/wHiOLLnk/vjarSf/OotFMjkeFblyuiGf46cL1WcBWpYWKs59x5FNZ9l
+E2CElG8hhRmlixnCoMxI4FHB4zCB2KwByxyZGEykPvTeETIjQoepduKtsK9LtapXpgW8g/cwq+N
dy3jOnQEK4ml9i6EhCH9A2+Ows8BOZzCN3OEgxJsQ435G915dwlUNlrKaR70nOGhR5+/C2MyDd3s
nRq0ksoAyZhiFy8qgB5xvpCfAa9Q21rQlk55f+uhoivYO5XEcMNgmDrVr2vw9W/kY8flvKiv7OIM
AF7VPigfdC7yjP+0xZmcXgdkNfhORlqp1BfclehqKlYO7ZSyERfYb5knHS3zAT9QD94NWTI1gJxT
4ydTKszCH+9nmaluW16BflYzO5l2OgVyxZJ6YMFI5YUD04e9iyXFF/1UKCrtV1lnyPN5TKUlowDM
ITNRM59jzf5fM+jYElaeQ0b5zu1QQXL4u0Q9EqrkqWzEMx3UbQOStfAOjFdBS54yjzTEJasf55hF
6qZnQeMibbV/WzGeIUT7JwFY1VaF6resfjN01g4/hUALmTmYPuMNaJnTwRYfDUMkYNjX8JzZJ/QI
XdrPpVdQPEfxokwlAacBLTAoKbHgqpHKFYIiTU5aAgYYpcz9WGKvlW63vbolrb3Yx5HClnreupsn
abhHuXdJ1H8dKnTSCjhXkgeOm+rDFrw7LJ5quU5BFtqYI1PvQRmwIPnFsa1k9sWl/nbaWUG8JSrF
tbRQNYSgxexiKf2M1ZjuJCZQ0TzrvMcmjKbTDhm4sFBKiE9WN7Yk+/JRQBOEZfwCrTshUNn7X8Zy
Akr4JswB9GggptvXhLtGgUKTHtmpBRJs7FGH11F7Y2pFsInxdQsiye9KdXv8ohFNAnvF57WSZDG/
W/lnd+wrKQwTuVtjmLHhkWqDVtRVEfYRzpKjvYR5nFRxGJLIIX0bOdCYlwhGYAsJFoq0czqSizD3
Cpto/W5JREb5xw497Vn4WZ2C4CAKeavSZp0mXbKz/ps7WsmVnXk1UkWrGit9vpKOopEp3hMwVCiU
QThzMqR29l75CtUSMMDpvElb0KPCPaST9QPbhfe7bsu5yKeNo+H47l4E/DUAErjWLtBIsAJYl242
57l0HA/a9BbkPJNTuxA0BjgoJlaH/tJgWCxgzq9wAkitALxZfXU+31w3nEJNUyFc5ocsqIgUdzJV
gHbLynIqCzZT9wOBgR7LxI5dDgByEXaDHPajPtlx6P/Zex9Y3tcPkntNcnHiWP04Hqv7sGO6rnLS
SvO/KYsKcAYV56Ug4674AS9ilfIpNfJMxr3fvFO0LsIxr4FmEuU37aqmOvzL6JSlQLn1pXXoVnok
CpRUwFbR3XHRjH3ulc6y+7eckH91but0f3WvnQGzWXvXFVEji4f7QpqEXInSbfS3+wE3efhc/qhR
GVXdBz3gsSKy+rgg0giXdhIvVQvHgfH5m+EXDvGlu6NJEWYjOm3Hm8xUGNYInSscEYWxVd50eO7I
l1OQSdfZy0PxGVDOhFCHJgz1faB9nwergcmHFvIbluJYaEMof+LSTg/Dy6jWXIa9RchUGI1c/OWM
wa191H5GJNBYfWHaBp9YWzZ+utPUjj5crN5jtQKjk+aWZojUlnxaekSIWhmhCEgkK8E3kvZotX56
E/OjKXdsU97LSoTifhllD1G+Xs9pq+U/EM0IcGUpatBBzDKDy/gYb6cCggr0pdkhiR4zjzIX4Bt8
v2eDjHu9IUvHPmI3c0jEOA1oSIJR2RNWOajfuZ8lqhnk3Ggd/aDlbONGBmDNpXGonQ6Ko43y6g2C
EY0s7i7ZhLHffdpHbGd1Apdh8EmABoPCKttEwexBdk2Gv2ImbPk79UW+ycWbqsgwspprhE3EYM9S
K/+RyqloBZGhP9ikzV5FpHq0Povj6ru5TKBO1iCaSZEzgp0HzUBJZ7DNaLYaTD2MOAwNcFbLH/k5
Mjdq4izABiDLpXM+TtQkVqyBrBR1xEjh1nqnn+VHM+c73V2DsTJOD5oqD9lxH9GnmsE8D63vHhO5
fjXe1p93nfowYc6OwL1P1crC4xICWYZoPRH34lg5abmECOMUcyKCN9MYdxPrW/S7hdkoV3WYzK+t
ODkcWGsXZUTl24LfJ6esY7cx1p0MP0JLrKXgB8Vt7iaU5ymkQUZsMB4AD0AcATcEvXvN6H14+CZ3
n/h/RCuP1KcRgpSuXqVIrSkAJHDjexme3Yh9NfwmdKHEwUJhqr+P0Pl2xFb7hwQZs2rpwI1zvixc
m0rImTLDwr80kghOwgqvi7hf4Fe6HGYA4nmfww3570gbX8u81Wl2LOEMxrrd0J8CBOCo4gtrf41e
XSyv1+MolKuRDQ/PBF9rKwNom7NXqJmZXzuuEz6DxJ/+KSAIN907Xt+Czl6tfNFjomUNjvNiHilQ
dNr3PPY2D8iZWx6xNY4QTazyfifMqNDFknu55p0p7D0jtjupPQ7czLT7r6BWn0H5YE7MvmC8JBRV
urXXvH75o9+qZ9vzeR/AfZaOvJu7v7BhlpxlIT8/R2IOJjPK9W+tnGNWGuhTAjw/shgl+GONBZGa
zj/G7oCzS55PswZH56DemMQcpME7Ih3AXrPb0XEA5RERvnGT08paoJiZAZ8sDdweKBpeA9F6v9TB
aILmdTfN7PU8Cczxft5VjQY+L+tSRAMJR8Vpcr/I6492zGWmrhpKcMzWPS48p/3yVpjyV+LX68u2
rNJTBjQXbJAAGsjihfvJv+sn7NrHGx8LPS842WIpgEYrg+/LmyzDyCDKUh5UCU44eTNLRqGx/3a+
hI0eipQ4tH9ft16HBdX/VufrwZvaa+v+bj/+rc0nytaQ7enkXXmR7Rs1GV+O1ApJo5GB2CvtoD77
hpR2iVX7vjkLrIO5t7fzYX+tfrVmBTCmDQKsqmt0HcLOe4sC8KtyL1xOmQ/YcJR6Xux7Vd6ma9K0
fKOKtkyglKsw+JytlIxzg6XDG7kcLmZDxJElU7Uj1+/aLCWDHXw1wU/u53U9k3yeIUwGkOQMGKY9
uEBpO0uMoNYb2zZZxrRgtfhYuYcXhCTqvT78aGh4IEgUexrrSXGnJ6wuwBs3MaeWWhZPN09dRGpH
TtAwP+me5PKSppuPS+zIm2aTe9iIGxe66j29milz1Tp0J7AtzTAlBuQXckZWSyC1a5itKXWWzBFe
iqefjK00K2+vUlCoJ2UladEZ+arIzRTSnpz/8tKEI/npGM9Bbv0P3hMvrt7CWhgVcw/4HCKXSy0v
n5zg65HSI22+ZoHvNWcazpolwil9nD6XS1en3IyTGFlD5+b79KIJ3s/a0TWefpIH/ucLRGOj9Ky9
FsOOekKKm9Kerw4FMUyZYhhA4yxBrjHZy5ofeP2vU6DPm+i+JGWdpjTxNEfefjqMSfnMSid4jskD
lelrZt5EDVuz3AH4lfmWmszwv2KT74xQiPQsQRIreGYS3MisiYDlGMYDqK7Bg9BHjprbJZkMNp+8
EqNWJQjciJ1vuhstkkTa6+lnj4QSekFqDSTa9UBuhMvQoUoCsQ6XAjdRexzPQcsIpIFGcRiFoTgu
0u2Smbwa2Za/P1j8C7OWnYamdjqqRvtPriurKJc2/rGiyoKWwknDKi/nahmHgW/ogAoVjYk6NH95
YfXEb7CQ42V7TctGsn2z3co1LLdhUWRXSPFbDRZ1fXsDSxdaszIF3v74ZvXvsVxK9nCg5JxaCb1h
8EcLIAHQNbWLTK3hY9k5ZJXgiqctDMFvKkQiwm0BgjSDdR5DpjJeneptxtvFAIKmOdTZVlkNT5Eo
B2jxKiKRq/ZFzfzXDK51x1GzL3/78TBfSQtb1VR7lOczvIyKbdbkd0gIbqP7oJOQafbnvcV4a4Ik
cApygilzkWAZ8M4J3KD+fNdn6sLX1jBhwmYIwZdzqqtFFSS9WIUmjGhngBlT/sOd5OFzLhq8qlHY
EGZ1XfKJ3iQ+xlsb7T8w3jYODbPynjLN6/GuTCRqsuquXRVijTIsU/wVqwS7yMNNcLElv06CykOc
rTqk4o5d2Iv2cMN2G4+PcpfSIRH4yL+0q5uLmB8Ox5zuhAHnzldsS9oIZCmlwcqc2lxVbjpCuizb
usKo1Vaxz0JBXtYnTQ1NkCoMoLFsyMnZHzjdURUbl+MTfsU6WmwxjcnzypU+BnI3ic8oKk68s8VI
o8k7f+YS4rXVLSSHTCM5Z6F6Lb3cdU+Fv68URZNsBAI2aYfkvaD9SBU9mgw4gRy5yOAqMNtbaSyv
5IZqd5s6+nfKcV+uMQm8f5gLcVZEYyfyPNcP2jw0ddJSDKpaVTr6W7Q5QVoNybKMhZ4ml1BKpuEX
E8vv7dUFM9ZJ25vVWwMvIkfweciGzU01PWVYEEEplqO2eWRtM15qLo4BgCqMBccVHxfFrVe0oSUs
GYXIl9VTxNeLTEK2p5XtvgZTEDXo6u5O6sXvQe5v/5CSKYPHzHUkdlOvpj9WbuDB+w20yhiYtskC
teD7+GTyivZ6ihX9fLpl3FYVmPdhh4XR95oaB+dP13fz78RJYiJRU/nPBMQJ5d/H0nxLPjfSOgy+
s9EdfBpepFA0/7fBPwgKBVcPeInK/b+F9VXSEuttz+syK3m2H24WnKJrHYsoBsStzAgGvy2+yF4G
lyADQ6XPZt1CvdxnxFjXJXUusnXqBSZLL63DIAg0DJKMEvdax/9KKff4i3My4MlKp3YKAC4wZwXs
pcXIGgZJcl68qAAw7IU9uye4LD0XFRbabgM+gfkvR6d01czZERHcQXh2/yyAimudtH+pujM2g9Et
5FE3MRDv9Jom1Qutw2qODh0iyFr/30nV5jOxhI/bYOCO+3UBdLt4ZXMjuyaV+nOURoelekSewBLW
DWUvhpDiag1GaljE2O53J2/OSRjl0rT3Bq9WiBIwguwUqEcCtRg8RXblIPf5Aw6uO3J84SFUzCKo
hxDRRNwrgzJiVIPyoYE3C1Y6nerVAxYjdyZMDqnh6VyOUZblf7gp2h+ttzmsU8ZG1Zf5f2vR8iO4
yu58EB5/LqpQ8R5dtn+XI/8TwXq1FaF/K0s3wg86OtEy+T3F5HxAFwcAA4rm/GMLpNtXWvrOxqUX
6thhvb8yQcAYe+mcipBLytI4lUkCDRJcB0OsuqUjK51F3+N3BtAs3hQ62emhnS6nWySDTH5Q1KYr
l7LxMxDbvJ6IQgrot60gWYQdxgPoCX3Rs2fSqgAbOYJgIa965PU6ARwVESlutPq24aXJ+ZVI+GxJ
Y3v8riIIx/14JhNHNBbIODgMgLPNHd9nSP5D8rENfiLZ/0ONzZ2LIrVu26XO/9a8Ya3OaLdyoQmM
O/AScFG3n++UOX7uaGQhHj6ORaYow/Y6WS6PnT2CRQuL5ZfDm5A/o5Ej5T/1j3gF1fmTv1SsJkMe
s1n0UslPaK8SJr+fHsgQxtX0Ter7RdjKy92x7PdzfZiTMmOkodgZJfEcUQCw1/r+8hnX62TbOOrJ
aFxfUgufoKOIVFvZbx+w+Azy9bLTSn+2hDq+OvnfMc6qF01cxJfB94DbkbUEtB5VIgLS6SuZ09Lu
LRgbZQnOLCH9sNf0ez8PWmFmPyB/lAQVy8b5duB4nK9z5DuZkeYV6lWgKIWGzQqpKMv6xvJqiq3e
Bx5S8mlJ2w2sjQynv53k/5qjosrgLIr/CI0n5nwP2wk0KV3HScZv5ryMIQNbH+z+07S2bRCEUsxm
B5mCEdgoAn0NObOTF4aMk9i86MHsRpfimSWDV/NEOlhNtn+HJODjzJpOaFKml2Yy7SkDP2BMDCzl
5WVm5WHBYiDRzQrXrCvRBHWl0HuPavOnLdlFbg9w9IrJ9r1kEnLseB5P+m7AMg5msp73IxlxNdnJ
G1AFSvyGJ4Oq11qbJ31Iy2RW3R9Vx32RZFkkdW+QWVp0XQ7gPTu537X+OdaOA8R9YHnzhGgo0ArF
t8iP+gPtRMrHYwDBfc8XoTus4OQUm3DZmrVjd9r0WveRSKdfehFeJtr5WhhR4ioIL5nseiidM0Hg
4ViOWozVNfMwA1eeojAHoY2Xvcfzmz/F4OC0Un2Ng3Is+Yv7Uo/WCkGBh16QADC8n2WX1vIGcWG3
sBPFAJfkHapmkV1dXiLsTlWZCTvoe3Ce5kNZ4beSyrujywd6V8YazF7bfiyJIISpkJsiC3skgzuP
WmvyvLsv9+vr/YEmSJGjBj+WtVkk0KK9qmmpZfz5MqxKw8F5//X0WApNXu83Y8vn23eotuy1SAIB
st8uvz7mQEnfL3wkgJ04ygf8keJfgouj03D9ulh+lfH5ZPdj6MUeEmC/ClH+uNR1WMW6Nb5/6Ji2
hjUUAgQItsINWrZKyeyt3n1r09RN4WJTt8EnGQB+iO+abGSsv6iadJ2gy5DpZ/5Mh4iKMWB1AmtC
ARjY/G1sjuga1YABHOJ0eIq1xtQdtUkrZJ+RlYQusvkFFKK6E5Q54CQ9RkBR4XbjgsGweJAzgdtZ
rp8nWDIYxoOCUQYcDcCzobYqYogMC+/+x7X4C158QFLmdBNLjzcWcBopEWPXbfLK84lUqxIrIBNf
G8o6MGDIjttPpnk0MelSK+3wB7LRPQBTAoH6i3TGZK5zq/mTSXXJ3S14CwxHqejeYMkltnqB3CTD
ZtCu0aL+4PwS55Gz+ZTxfANSo6525mnFjCQVLFbfTRUCi+JTzec2OZfsl1c5WQ6eZLl5hqrHVtZ7
KS0Rbm+BaFTNr25XzsY3snSpzR0SvXYgfmeOoNyU2UmFLpfMlNWMq2zo5Om/3tYswQXsqMVfgfts
v1nJg/XDE4ngL7GB5Lqe8LgfzP5jydnEVFfX6ya6hj6mSVDwm95pz6HnnqrlgMiPqKJ/0ihvtZhn
EznUyA2kHA1aGvLF7AqzcIKkAIYHG/6NILPeiD2iSN4HZ+d2fciuUS04csXSjKomfLPHnlWqbGp8
g7UOssmrKOW1hnL4XUNexk/wP4Ic7fE0KxvwpCViKVb0j0RybMVlYoeee9BZhT8CneRKWTDkEbdh
jUAR9ZUMTNBDbp1606PLq9sy6Sf9DewDwgWNkTi/PYUCjyCevdbFZpKvNJWsIEH7/I5bZyFLOeAt
YV5yadDHg4J44rt5MJsXxEAlQ6A/TbDbdcO8/E5+8wlSCuMKKqaQ0gec1a8PCpcsrUIZYSaKgGBc
n91gDzYvNBDJxnuMGIImXfSdsxzOlWSiNYloBPKq2JUlpem6PdN7Pb5GZwPuLzebiCTVxrmbwknR
sTTz6v1O5Cp91+yBBMHOpoFy1YkRFvdM85JB0a5z+LnGkTKq4+yvQYFRNg9LRHwDmhHaGFB9tGe5
jjDbpd1XIWKNJgiMLLiZLlhQWgQ8GDYjsa7xSC24Dk8prOGrcrK6HiMtHyRHdfbU8ApkRQDdJJud
kQiO7ERVRhmCMyfdyiVAsXwd2fKGTyPiNQeDfhiKEVlfR0tNQeLSZALBxmZ6JRUDKbS74Q3bnUFk
npVhWAMH0jUgfW+X4quQ8zNOA1JEyeOnqwE4AcSpNFMfJyxvkooZBPfMMRgAKaJh2xs2+D0jZJvf
oGOGTKeOrJqYBOYOh2/01l9rCrc7pPvJOdanWJQHtbblPYgW+JsPJYd7zeOxB7O3X0MI/7ufIZ1r
Ea4cNEd07YWKkoz53Vur38Y6RO0FcKy6dqWxsbG43H+UivQM6EI7nas5DSoyFED5/hL+b63EYfe5
47rHBVcwbrJT7oUByOjgl7fSPLhKCvxBWds211iF9OAo5/soze1PmZA9s3HiichbUXIcNpc50gcW
vPOgW6LqGJBVRemb2WoNG4eD+4355CHKs0yvwOBHEkPKOyuPm+CqV9/CjNyqRE9e81ua7KcjBcb2
jv36M9Ck4v8EvhZGCa0l1LYe2CbdIkMuxvqiiNpo4LhIqlk0rr071bafHYjIaIMsroDkWIaY5OSs
Fx9IJCnlTDEk7oJV2YSczGwN6L+CSSavlQ0y2rAmt+cHLjTyKy+ZYqsZDXQtImO3zxP0PTgE3tLs
s18tUrmxfA4ggNdnAxKUoToEmXQNFwCU7qbvjVqAcChZIHq6k8BbAEKUYgYyR1kMDu5pPGHtg6FR
WD8sc8+D7nsvqEiqhsP9MRDExf8+uJU1cJ9Eb12wcU+9Ml30omx6sI3k5/lCb/TGxWsowOQWHa4B
WIstZIeVJD44B3HROxyJ+PfpHPTRvVVPof4QMMNFHzOIwJITBh8Ud8+zUOrnbtJwxvbDWcwoLoEA
nkP0gieWrXIsavO1AY3c4QplfweY5FvGawKUFS1k3rh23BOTAi9Jw/7eRYQp9op2WogLUOdclJbK
UfVnNOkR6++ruf8GRbyuf0yOau+GCiXIwH02cjAWFUP3UPRaV12H2rSaPh2Vf6fkF8mynNYLXsFf
Agz7htUprBX46e2qheeg9ZfapYyQ6YER41dZPWGhUtRoi260bJGZ0YTmoQDXCHamDpDpLtOJrz1+
01Q/S99DGnqa1q/V2Glqt4T2bElAI6ZHo4QFjmECHG/T64ZTjr1wtcGG0MDI/Oa68LJMVCubiLGO
nkY76xYPIHnOANL3q2+VNr4OnQwMg4UaKhYELziEDdL4HnDbEfvdvoa/+94N7u7OWPUOR8M4wQjt
nncd00hG2gdTdaM3kckDQYmIhjeeoXMZQk5/aEAma5S0K00gBDWMlLh4tRG9piPiLNCbcGGJ+9Jz
4++8p95e/+QPB8TADXUVwFQovFwpN8k8wNr60R6qx6DNusBWP/xt1GKShnWN1PI/YfrFcG2KG8Xi
z1mndKzn8ntU0fnHKA8Iu8hoNB7jR1NMfHve9wSFVrAuRFe1cD1avEGQ3o8iiAGUw0Q1BPUM94uj
QKmBEW3m/Zj8UbLmSK0mY+zt8OLuNtRkrmkyuAFttRLCeJwGXDOYislgKktdR5YDQFOqmNE/AJJY
DzJxgBgNLGRNtcncmiwiDUj9ZyYmhvLcVqQBQdGDkkbSHdhHcoQbBMbh8C/bTY9rizXhnzxb4BBE
DgfuPDE2jB6t4Ya1zvty52/PYrXdvR/DDr07kkF2h/oIPpiF7onG70x50HLUFAVCCsC83tBNCM/p
V6mt11NWDdDZfZvrSASKdHRAKkN+Qjun1d8qVnHu2dYskG6J9AG27TzbjPkD75GeHWkBfCv2dI6u
uO585J6MHwqDkF2YV6Foyn0b7ch8DhVJbdGsmgyt8qWCzVeHtz50hs+/39LlZaKTIWNb+XTIN4vs
NUiW5HVPVQ281/ZPkJFmW6OT8JgYebpDMUcRNASmgkg7udGbea1THPa/ZPQ7A78Y5pSwKq5ibN0t
ez4zWj5XTMNR0ufVAJpOT8dKdNIupyCloCMi1orP2xoEgvA4pYeD7DaS/35i9hR9qYNBAI74qMOx
MqWAu5T+4gZzBk6Sxpsh0kJTDZwHQNAd4pO709J6EmvAmfB09fBc6ML0Xsmqq2/pk/KsE26brZtB
U1wQFXYofxmvsbuBhtD6FSNeB9iWT8UHL9aOfpbKDGW+bq/4FBBNeRfAaHLTTazuO2JWbT8W2knD
LuwnavAN9XPKeHM0ZeAHbMNQ9u+ICIftyQXlDuh1UhbBMR2k6LD2d0Wv6JvMcmEa6ToIfMhJikiR
BkTaeDZbdrd4RjDNaHw1bS38z1OtkNINqYR5U8FvFGOYLZM63He3WbFHPq3P/o5NbNUBWy5G+xP8
BuGyK/0UGAqNMGRMHqTtfAtNMBQbJZSnQwi0j71J74aIVCRG585lFI0CNJ3qpG+SXSyJTOw6Rd6e
zjqg3J5m8HbHlI0nrSIzjP75jM6Pqbscf4P9eFnJvcnmRWyTRzqEW7IOamU16zwTE5WwTH4Squuc
VmepNMNNev0/RR9vYeHIM8AOUHdQUS9QoMYJnBfQYKXNoAZI7kay0CWNYWZIELj7yDF3eNerrAks
+pE3WWFRTGN0ma0ToZaCy8i8EF3aGWQ7Tf/nh9HX+PlUa7vMUdxZ+97PJnoHcsoswZz0OyXX1dpn
FnsmDWVNgsF/zUrnyqZbzl3sGgpTEhVcwht8v0d1OxuOCVZAdDnWCaJwyMVYTWtk9xMjn6RJ+3X9
7DaZom8uC0MJXxC5rscjV9TihiKLKV0B/C7SOobCggficiIO8sEf0myKJJyGBQzfLPzIiEJrHbxb
+x8mCWnW6nDEZWYUY6et5O1GCZY1yKZ47ddcBwReXbtq/coxJtBFarnkAMYIFURl++zkhTa5arWk
jr9iUyVAWx7hMCjnN9Fc9ULaqxB4d9iQih6Qn24hS+EnASNluBmdHh7+0bZp7020leTiLP6X7508
3mRjwwXzuJzavfo1sSinsWS738/Lioh7MCi88+NTmBuLv49gKq66TXFCeY545RQdKlFuJVjPcVlw
iuAevRskrnfrGW6n5hdtyfwIHchP2bGwmNW6QR/uT7VlhbbTZuxSkmQtzAuSciOlY8iavZitSy4R
hjsIA2fya6Gsws06iJDEcdSeXlLy0YmWgixnYvgTcV6xqIfjN9oTPV1c2bRdQi0qYLhQu76xE9SH
TgYpXMzcaxiJcATJcLAMN+/4K0Vc916nWWT31CUZwVlWOLG0JwCAnX75VtsEI/Ya96uL9wlgXm7h
8yfqcyFQYoJYlfwJe0VvnUfXFEW4GFHY+qjKBgRn8jVvouseu6uK2Cfq06X/na+DI0BpOXU16Tok
R/CLlf9uaEPDw8n+hwJvoFhQYps8bwPi/WHdU3xxQLdsuv14X+h7ShNNf2H9R48KXskzwEeRTjUW
OhJtTAKvVYJrl6uKEqGQtKtehGSOnWK+wV42ay80NU+BMsuko3l+Npj510Bgz5ZcWa+JPXo4ywVT
PG+hIpN/1gjJAJAAFVBcyDBJPUf78njuibw1B87E74d2EMs6Cg9tsrMSrpSQhFHG3Bh5MX0qm9HV
caHOrffmh4Hc6IelgDC4mxmdcPrJQXbO0qZv+mr42lMj0bX2UzREmYaimj+hcRTxdunjJQbS60pW
wn8LfkILCUgL3iHcq24+4iLllylxhcNRkbkA+51ER1c2dSbNukNcyF5SHd0AUX9WoEFjokjXHT6W
DOHeHwj+oPhOMp8tLPikN+PUbj71gUa3L38zKYyKLJAVt5T+KYIFcdXhev9omHJritfBXrJ85klx
V3x+EV5lODv+QtIifpE/WTpjoDfDqqt6ikMzscTcxpfrWpf3zS+idrZQzj0hxPuyqu+ND7n4FLJ/
Hibqk+dVLoCikBfmxWmEYKaIZzGb5SLj2aIxw4b5p1FwuJ2L714h/3gpqToLzMc84tajy5KYrh22
1RrCfup1gM+WRG1LZBVj6+5eN5TCsZvOdWNYumL1SKVQU/UjjTVoUJgKHxbfCGSyMK2yQn5x8h/X
MgstpH1yjMqlY1sW1lprKvIxixIUGKe7Adbs2Bd6aRuwWqlPuBPOXU3FaHpApke5v0a2sq3/LUKS
iDsyqTXwFPHhjAFfQ+jCcfUcEK8iXlxRQLfEGQDRhpDb/LAP0sWjXE+6fZ3Y5d47lugi8yZ2ybsy
cnv4fqVNZ3B3fqgfvcKlV5gdWlnR/rRGW4NCs6Li+ES2pCRVPFLKnbbE9Yi3JJ7b8QNMRyztPdSO
9Ki1w22knlBB/olWcKhU7ZpYvful7fCM6sKbkG5B1kNzWe4QxCEilcz9N+fNCNN8kmEatcq2HxpR
MvxapIlwLpwDu0GyZZYSTnLIErXw4tNuiaR4aEZFV6X52sG/B5FqCHzst7s4YcOjrCY8tm0kHTnO
fQ/tbdUAQ4St1XjG39fkhLCZ4/tZ6t68jIEipxiieJJhbfyrD77azO7lbFvY0rIAF1ege69+qRSK
PAPIWwWt/oXOSIUgmGuTKIFMP55P94nvYxQEtHefoNsWC4Zx97jIFip5sitFs5sSEWb2+6b7gAbp
UjTChvoEylWBkKk7tzevQQB23IzNqFzUj74qc37fvIMNEGjx7t5KmSeY8lbQIJXNq9uq7BtLE7NJ
xYwBs+q1oZ60maxQk/AZq/uPS1vXMiN/03RKtdrJfhQtg/ThOQpzIY64kdnjGkwIVepm2OIwOkz2
Rmodygv01aEZ7E+zLDUTOgg0WerxbjQU5bTWA8VV7I5Ig6ddy7uB/okTx2u9sg3Wk0jUPUIHIppw
Q1QSsSlzeEfLhRb3fBEPEph1JJKZs4jhhN3xq/3OthSMclgrI/YSaUAdg4Ul2a/CK1MYQ0m8yDpX
ZrsLx+AQTnSK+naKu6/lSM+xNJ3IbOu1jTiXIYJ9WAU7tV+ndE/e4xQ1o5wlXEPAdcvRQppritWx
6wRymGJGydSMyNtSqdKf3aE26ioWLvklg0DkSEV73prEBKpL6pVKXoZ6aUoVfoG8Zb7CKNEmGl8z
CX1/KfgbXRj2bdI5rPepVEWZatUnNdKaCWf20CXSI+OzPmqaQ169qozfgsQiVJVZGIKo844UvDI3
2puUDf7oiwkNm9oWYg/bYvTbxcWN3GxOvt56i5xuOVjdO/ZlB0cE2+QTE5z6NXO89SPOGvUsNRp8
8y7M3Ubqq3eGWwA7EYy80sVo63Hs4ywtSToIfwYk5l9i/DX+iaGTrkatcrfBw1yHtPuReEwv3pjV
rFjvmxDCX6HtQHjNOISDluB+hkGqSYSh8hvdupgzzF85zMf7fXY1V6V11ApzupQIae8gDvxuuWVa
YeyzBczHnJUvtaFVDdaEJC04A8mKoXwQGTgrLgw9g2dO3N30XAHQqLrC0qMQt6biUTmu5eoxnbWp
Mr5fG3S7xX8Sj3ULZBsjeZdP0om5Lj9IYnO/vH2umsOjdZfgka9UTRwIzVWd+PmhyrskCIipiSDG
eNYhQr89R7XQxZzSX2s6OdtXktIuNjZwkXUS93v4abd3cv22yn209PhlS45corUP2fCeS9JzK/G0
R9vHKJ9YzO8AKG/Afpk+UnR9IvAZzMBOS5Ruo6ogtkvcXnIMCMO+Fw8GnK4NDrcrLsSNcbkeHSSr
blGlzwmy838EgKu9coeXmStNu4L8bdSydNteczZHM0gUzOYUb5nfzzgjh6BsmjrHPzish5qf1sOh
CzELfd82UoypWCzYgBqwFpKd3WvAnyvnMmtae3R/Tn36KDxXujEQyNs3qX8+WihMTaU6MLmfiwll
Wb/tBf9Oo2iIPvFyh4QN2oUhOnfw+twaIC03+O3xcLCK6ETPCI5Cr6gVlfXxjo4NwaqlLivsiwdN
OP/bH1kpagFFyx0Ie4aP/ztCSjO29NJwBbFgepYv8DSR/Q6SGu4JyIHUdhOO7xg3sIJP2BzKK2Sl
OUHFD9m2Mk/OnrSz41+RWdacjbEfqLhVMszlRzZb2cJuaKujlA2kKMVUpvtM9FksAvBK8UYx1A31
MFhghhQgNkk1Rpkzbv3dWo3lcVUBW5LozprqLtrOlJAjh8WSKNSC7o7LtPgehdHVyfuST0Wtt642
aVDHwx5allTG6z9HGw5Oc1dG+LTZFqReduJeq0oaRlVewqyBdqLhPR1lOsEKDIuEyIPoUG+RBlX/
BovQp88+B84a9wZibOhJTF1d8CYG5PuDM6oO17mUueYJxpVuPg8r9odvCVy6uUuDuW+JYRCjSd16
HJAVMd5EqLNfsmuqpIV93wqZMS37bogLo7KkIWqXR5fTMn27Krn2yjeRGf2ky7xRmu+LF5QZH1Cn
Z37BAbG9MKmIQaGh+pdmBNbK285OOEg2+Cc7y+Ifma1y5jMWVGLRE+xSQAaVXc8h2+wsDnqQOvB6
drBq9uw4sA+Q1bs2+hh1bWMvfAXnSetW7UJKPP3arsbHtnLEwrO2IP/jYB8oEQMyK7fEzKhP1GxC
TeeBd85hdJoa+6aOhXxz89ULl66F4W5DCEWh2wQI+c5glUG4HNOqVBzoDShRDIfQ6gwvHDNOakTo
sAfVvPZvF8BBMvRlDrvIEHFiIOtoH6mwJP4dp0f6I94KuxD/iVEFknWPjkaaYqMAhWmJ6RSQ1/sS
f/l0UcVKHtvmGuYOnIcOh3H/d6ljOiPcNf+68Fw8W7jhrhAP6m4Ts9nNGQLajjI5kib3O2YSf2k1
WfhEixc70UniQfTpqPWHUesUx8PLropHGzBt6Q4JzHsDOhRDgvnoKw4NOiGS1vlaRrfj1M/agRKL
nDPStJVHwaeuIfz/ytRBwSQt+KeJPcXTMxrX1FmsiyA6rlu//bdVwX650yBVW9ChZKXZc0qWBRmG
yPuT3CF8N7nyEYEqO0hhDD/7MWYIfD5bDiEztI27VJeFhcDvg0IHepZf/o9p4ZB5mKNRugQiXSxP
c66zGH90ihkkdRSgpI/q2ohoxXi+e+DrrZjNg6kureKzbA1IK1x6dUTN4aAgHGNtwlje8k8LyX/t
XRfNa7WwLbjn7Leuudeir/6G9xFQZ4aBtItYphW7PkupUoJUkBJ+zKKW6lIgPqrvUdboZ4GDcIJX
65sClPfmFAO4hB0A9zjC+AJfvpxCOCAjSYty64y3IEtbhqagqotztFUqOeEoddwZt82+WDYVbpI5
GGzjfh+Y2qADu9c45m0rKCCYRFnOqLMVRrndkDbA3BKDJVHawtZY3++be54VUeqKVRI+1GEi6rLX
O+pFk34AFJv1N0gDmbyjnec202ROGHkaX+fD3keSBRz54oHclYJHK0knL1Nefl3lAR7gn8Md2ihc
1IONJ5wEM4+vUgcL3q4LJfamziUqa+m+GAg0GeaidrzmMVv7yZRd38jP+Hj3TCsiyESpch8IAvoj
GgPoCQRIDOd2sU8ht4ihSupz7z8JGkcYL7Zv63skmSGgaOJHTMMZF03wOb56QqzBNaq12G9+GoH3
gGrk9lH7nFNTIDlrz19nIE2o6w2/BUYFba9iEJ7r3Mum0lvj7/xnw4ODKTlZpltYlictWp5cO8pl
Ejb/SsJLPNHJn9ys7czyAIJxx8lguhXAXHhoz7E59r9/+COE2Qbjsum7t4dbjhmNs8rWAMgkS4ot
7s4lMv8NgAcJCFIF82Hribh+98B3R3dDyURdXhLDUTb3KBgn2wxPIKPGQ8TCEDMcCH7C20O0LXia
an5+rLWKDUjQhEtbjb84UxkDMac7uRL2YklLNAqAuovY34IEbm54mz6AORsqq3I/oh5s981HNC4I
zjPxqVW0zDj+o2s7oPkxnEQYeChQEp01cPSNhRemBAtQfFQvDLSJyILBn3o52GFRttpBitGlf3Lq
E0oYlLMW3pFDz9T9YQ0AFaN0LzuJbhhIFMlx/u//eb4gB3MSnBrYlP8abk9UX6DcC/8XhJZH7Bih
nAwlNtQ4W6Md1YNVY5+gfrt4w6wzm9vJeQw1T0bpM52ZfRt6oCe7pf72hHO2zCSvEDKTuG693F9R
KyeoQY2nLTjmz9poF0Dtv9rO0Wt7rAmtrx8cWZOU2aR9RzxKlF9RqLyvonIdgC/CjXni/zzJJHs6
JkqrlFS3LSWXmzj1Onw0SEQ6r8MXk6O4IX+eXSquBCgL2y0gR45XY9Jr1DWJaiZV1DLbhIPVilpz
HrKucZ51SQ7ex2eJ6qfFLsrOaXkVyi5XpTr70oaJDPRNt0qOdL20/sgbGT/VXoYcJbO3gBJpnfjU
kCLWKCor3onDgIdb8eWOoenfICGi6OYf79lfDaEchztShxpzI6vl2/k7O9qMUjDl7c9MGnlgIwWL
lvDJwbjQ0YAUajRWKEKzVxpbgSZnOthrnIzYHlUblLtVUUfvPKo+tcB+VYfCOyWU8l2Em6JbXeVB
1vdf/TjHOXboC2oDtSwfkXHYQilZgp93EgZTbJ9ZH7PrbTPnBMeyZUejAwPf+zuhjP8HxCjWiSqA
ziXn9cbnIxSfOnSHJO37wzNDi7FkudBdcPnrJOqYSiy6tB/JFCieRhNp6dHdEv16N54JvA4QWL1W
lkPjBpmLDFl1hCOnF6cmGIZGkmuA+u9cQYN1hMTOcLsJCwXxcqehVSjDGe/3yEyQJavAi5ibCHkf
n2/EjIfISmyYR6fdLIEH21AyFV9gri6wiMjLnuBoE0jqJmftgl/zBPJNA97+E9GeyIlKDvRwhN4i
/LYMihcRHbB/1ZLd9YKXRldJ7FfmQJ88EM12tYMiSswecEwaQBHe4cd1aEQw1vp1jmZdOWUxRA/1
Taoaf0xcWFKiAR8huLlsbku6q4YQRg6Pljt1TDJ0Yry/b6Ccr1zIDaj7CM0niz1wEM/z3NL6eLaQ
4vKXRb35PxgkfR2YXc+ze/x1clz9alxQ/jK3CWprHNVTGCcaqnRJ13daqudhP0wLcF7f8QffHB0J
EcwXeKiNxpzwZw4PpKH6vg5wnrTm9zFZ0wjABsFuDNIw6Hzxp2er4fRqOXW15qCl7/AahWDhjaHC
xp8xIKPbZ5Vh/PYljdm/BgXzjWRsZYKRrHJxqnoN9kSloapag4uAm45oO070WAvpGy9wyWs0bqXZ
COdgbD4zRkCpCkzjbAoWk2rK75rYA/6e1gDEzibJhNDWysbUcYmuBAs7uRB5syxusDQhBpLe1X0Q
ti9stLuIjZo48zLdJprLTU/FumTCGZLiLcbIY/swskpOg4tyJdtHdbHpNcK3nJCmwEWvD5OqNRSP
9byEKkiEMyAmEaWNMWGN7bn4jED9zfogDR+4BtzX/YeA2cnNVx2PXyDKCFLquaWRopyKab6zZ//G
3cZMqCrGwTP9VbzP9pxI1maUi/4jlYCNb0BGAwIpsMlGYnnUFDcq9hIU/asiJTzcsVyIL8OhlbIy
vmXYCflYldyU5mQnRt2ZUr+xzhT8cJyFcTQBkQRbCyhE3JUH6fjxTPLv9SPcfszfpPxTllBvdl9H
epWfXASdLqGMKxya6o8jK+TBdyVhZHktfg0zF1tuGn6g8tQjTilX0qKXvyGa7LoelfEpXY/WiBwG
sTipFIwYd8sa3y8rARtOohXn1hrtvvxvHDnuXHbY6vQvOH6biRbvjafxcin6A3s0bHttxHCekowW
E1i+bAi28O5f1oN8Q/eyvT3pb9Z8RgKuWmY3pit5ivVSpeFPry8PK6FqN1W+2KLk5EjN16S1MFn+
7NXH6Sb5fU9QNfeLHugihgBtImIR/WMVHBoeYMadjPoBQ0FbCJIpSNYH6AKqJOK9PpIF2h9/1bQG
bvt3yGGgtqvaUxnXs+tHDPt+f5DiDYV4TrlBdb5in2+rrqnwW6cQciIDPEFBn9zjsa2QJL9t7/zU
Ns1b2jKVY6PKWNiba9yM899g2/W5bWxT+hw0mY4LZMBM90BvyhlLM0931LSXANVd/ZhjmbJdr5/a
wTwirmQt5l8/RMuW7FZ3OXZA8HBXA+6P1Oc6ESgFAbf4WVu0J+ovstZRKP5lJOMe1FFhpSEx042e
RkLI5PBuSOlelfSJz33GLnBCPgiO6LPTDfiJVtk2Q5EezQC7BfFPj81YPZWLWLpKnwZ6o0vgyj1n
1vfuCnTx6xAnz0B2Wf1WXeEn6/clqO7UMLJODqY2Z1hVT9Tn6HTaB1kjpfjC14mrHyP8m3NVJPgR
j0NEvUC2N3PbydVW7rOTO3bZzPaZfWfXaL4VeYZ5RMnsL4Pia8r1+bS+ew4oVrheTdMZc6QssV4D
vzaBoEKnXHeEV0BBnxPzDV8dAaVUoVtssO4+v2UPhDsHn3dicRkIUn+ZzFgi7b7Fjg6KxNJCD00z
9OjP4NCIABn+wo8ICh04SIUFUSNuMS+qSKE2sI34NH+WnJdlP8+IoKQ/XOjYdHfbN2ufHUIzRONg
ass78p2d5lnvjGsmCEnozUQ/FxTSqrzh6XTTLKUA2aU8tE474HYdQzncBY/QfzFmphgQzqa1NM2U
vKljPzrtm1vg3U2ayTP1m+DZJm4vkZ4nXwnsEGmyf6sBpg+thHm5GCFNYwWPRJHJyzHmIdNWD7Gi
W21+UaOO3Q/S+V9kNFPXGxvHZ7Iu2YOwagDkIpvgQ42yqXFp0ioKK2H58X8gZMgvWs/51mbq0ZAo
6TQXEqFKslq/2j9mzDu9va6oTVuUFeDhLPesLtrVOXVQXzQHlqePx+EawjgUM2Ke0odfI1xlgL+q
72DBXgxqyLZpXTaUjmDtI2oKVf7Epmb0agJhGfq/pvOKMHLTnEe+UMwhrDaniGOxGBf1NJi17g7u
8Dxekoi3DcPAlXPME8aGrnI2fNpik642aeXc841Yf60yEgK0ICwUK1opyII7rGr3WhG7p0CoZk8Q
uZ6xaOzD4AnhCp7MTu7GtPJWvXkIMhlDX7Q0/2J63I/y2tspZOy7YXYG1ddSvn0Nx4WP3ikHHjzX
VHBd6XKrlfm/E+t8uvC56/Z26MGc46lv7lX2DQwaJzB/V6sIbZFeK79tlN7Bag4/TxSwW4ab0BRc
oybFNU2+NaGG/EJ/r3pI33bEcQKf8IQTVo4KHm346TzBEGQ4S62VXYg05NuygLNyre4gqzPoYZHu
EjYCjmQ9Whv8TdqBYabGZ4z81vQxd8bi0jVEzb/CHXhKlfkJkZhuOR7pU/hY3OUVnuDdBQhCjcZw
ddOle6IijBtXd0iHZy2RSvOit8xeAEg+v1AOBrxEVTYlup1DESxC46NLjkZ5/AHLjyf06l9d7gQ1
TBHEpqxVQpONI0I7tZ0hQtVRgxgTYHlOm8wFPApQJP+LAXazv6v1c7Nd1Oug9Vis+awE4/8f+Q5R
obAyaCeggiMxjlPTm64Iadi0eSCL14VNHMLCDX3aAFXRSm/fTogGPujtK2sjW2acReVVh8tljXBw
8yFXnDP6iR6/AU117i+6/GwkARGFqdi+Zq8hOAd1v1x9Fb6vtIC9AJjFn3vCB8EFG5ILLjwPAqmj
h17Ya+2D45IwYyWmH7cqdWVmyVz7DIr8kBppCI3OnqNq9vW8IJW9A8bXnDZ3RmMNnuGV0/AjSUrp
FWpcfmmaOig4fzXWDse9PYvRPKXBeFj3iK2yV1Bb0TVpCPwXlvG3YSYwgCGdByKtcUpivCh4XKOS
aJwOyxpU3ZXmtp0B9A4y1KCkFsAw9YwSIsSUbq1WfcJ7qM9CdCAQMWyAu3YxG2LoxBjSZ21tFQK2
dibn1NyiKTxWBZg/QwX2JGqmXVvro2/GkHp0g+dlv4i3WFuBvY9rAwmuf+aJANnQICYow65CmDAw
QW7ZRusGtlh0XmFaFlUG7qI46xmVn7TqwZkQ0aoOetLqCOezkTT9ObeuMFPlZfGrhQE828EjZQyy
rO5wdD79Y8FKY/XZmT4l1qPg1RkE1G79XaGEySGRbofGtPHSRXDgyOel+ceTgpmy0W7r0I3XyKiB
O41NjdwXUmoTGMvlNyKdINfzam23yn86qmLPncZjfa7/JWAYByGf2B8lQ0fOPEEiD94+5R3vHbKt
VcqTQl7mLWW6lYZC3BMGhN2Nd62P0obHYr0Nm3m0+vAcu5qYvp0hCm8uPUH2NGSHPJadLMhMzJmH
ho3CkzxpschsUMvTKWDeuWboFcqeymPTPiz1Jjy7xnrBOVYSPf3oZuJbNrEyXberQ3fqvDW+X15z
qXW5FlHFo/i0c/1tdcRD83FbIKwj0XdlCNnnDUz4N3WMmmrxK9ixAmojk83n/ooKyaACUYIeq+kn
0OHfH0U0TFP5KOWqmS6rE0V4hgL4TxyEVJZ/2RXfCA5eTyoFD5H1q+ONmFVr5TT43X+rGHzVzyOA
1rk0eNYF2zD/hAutPLgFc1aZhSMb4EM+ZNreWAvknzDnNKnwY6OzuBS8YQRx+rjDRXDaqKwVfTVZ
bZB+NWCK8jU5bVQ7eMXHLHJlVdclF3A8d7plh11C3YenWoY6+aNGQiBOdM5tX/rB1IQBi8UfrkmR
OnTZFwhTDxCcFToGmljfhwg3rrZvAzAH4+7vNPWEHW+JqGAq7d2MXlybwL1fu1lrPmKT7FST7nrl
tn/anQOWaRbyGa7NtGABSzrt73b+S7c4EcWgeWzOUSj40yjrTurpwLrWkto9U4bPcDTUqnyzyyIX
YRP2g/ZUM/rfow3QUO22kDcnBNMxiSq60tUJL38dOCVLYmk2gnnuaBIkS5cDerst+kKp/yy0SuyL
YnfGeGLDJVMFvON0cyoqdQCTLzKZrpzBOMsXhJc68jgboc0/7w/xgLLQYSX72cyvtYXJwaNf1uCh
Vgz+Gwg8OEwW4eLi60524kzxyyzldbVuNXjVNy4590m5LvQSNYoALMxlFMki9CCAYuvU/W39WHdK
lfHsV4so1uIWgdk9IY7J7zyNV7cBRbRbF3qcPmE/RYPtfXf46A51WhUWF4il4JQ9VTiIevmSWAn2
5fvsIB8NZKgAunoCAGErbDlhwJtyb0EKgP8OAZc9SMBEM+Pl8QBhG7sa5xnazRQ7QJ6YhER8r77Z
ZudOv0Ts7exwBMjv7oXTSNOMa5ilQ8gUpY1NmLeDZNPOyWJwrlgx02Tm9OmA4zItgUMI9xHv2Y9F
NOtGBydpvY2tbhDi8QtCq9PEU+5YZDB+R3nijer1n6T+RHbclOkDqyGYt4ChGaNIB5Trv0EPAGER
BK48mamiR6UWt24qq8RxFDzfoa0XRzjmHZdfkLa98UdUNyevmtZ8Vbtzv7IzcvMpVlA9jTehuUjg
QWU5thZ9qgdTesba01u3mmMYqaHgyudUviexeyrXD9efIw3LmYCYrAJlBvFVOMF5fOlE/nflHhKa
8/sUzc1dZIF+mv/r8VsQhZy7V3/L1qIuidul4Mi0cGAoLn+ld3NNhSOne+F2QgUGZq/gASiMiPEM
aA/jzUZiZjmPL/Rnr20IX0Ib4+mOZeqPbT6FAylxuISROoUFkgMpwnihXN3PYUGoohARfBq9F4I6
Umg+aPksRkdf/QgpKD588DijKgIzHqnh5RKH53y2wMrqPv/x18LUd63wNBoOhIjxqMT+iu2hvf28
XknOHCq/AV53OyyDBB/TLi0I0zbHobMskJZGdgn3DT7HM6XiKF80PHre73J6JoW9aoEyDn2VtQK+
PoiSG/8BwhZ7mZ8njfMc5TAmdR/FyAu6D3KvUf6dpI5acsHzsjWQ3wkiFNouLiINt8Qkfc6qgBrt
r8X0yMNpauFO1by4+99rKEu7xGsfE0kAd80tAp+Qv57D21ISyVWRQU7qsFa8bwBRv9XtC/7F/52z
/HiFBW42QRVH/IjvltZt6FvqvzKZqwPPzXRBCMP3gNzwlTkzgNdv3yhuXWoTz5pNDED1qWanEeue
blyyBhDbGmM2j5TxFYWOpJ2MHQYt245b9vOFe60f9un8ZIsR1THhVDKhbYu4np4xjy+igeyBYms6
A2GGnIp8LTBhKOxt5XRoNJw0JVUlY1cA+VbBigXHs//WOFjByu8LiILehnUzhpXpm7k/eyGETZAW
ZGbwpbU+jX8nAkfTN6xCYjcgF9+FyAZns8FBvvDCRxiUiDb0HivLtnPfBUrEe+ZrKVUfovrFu4yX
WI02jrv8Hl/LoH0Wn5kyoqmaA1UX8tiwdjhP82huWc45ZB2zVSIHgDVoUbE4S3PGlK3OHqhXU0Au
uStL5haDhFEg3GDmGlR5xBeKDlMQj3vQuTH0448ciL3Pc8Xzk5+tNiFgMWcS6uHD5lIHu1n5/pLd
mp95zsoMneZpUnfSIceglBTlax2cdqxYk1FMCsdVN32P2Zkk7LwPi12BlIB1EmfZEDrRtuF1h3PG
fkW5DOqSr+VlN1n8EOCskTh5v4Gt09i8cYfb8+y5RNKOYdWpPf6MEuUkdLolqxKEeyfjzj7EzwHz
1T8HHDfrqFMeiTQA5i4CtEPxV77nZvUHnAqG13v94mYdaXinepFGwVgyrfThvLOaz47/eysv04O6
xFRw5jMVLg+gWcdduUD9FDxT21QqBWb0cfAt5ULBG6dEmmizUUZPodJG3+f1jJjB6l733sdE3+Y9
tMOlUqL4QqaMFi9+f3Pdsc7xCoShMJy/JhvGeNGUDZqD2WKqd0numjwI2mhgI4YWVfYVlk85KWUi
p53A8QHoijL6uh3aKnay2045ao5wCIJjhFeDdiu1m5Bo6fhmvxZlgwnaY4zBOT24rID1weB0iGfH
+ux10V+oKdcEyHRHQun/jbQ8Pz1+SY73AI8GJTg4Z+xGF+ja0JNqk7vr0BmfpqvoF/PLALYXX4qe
EDDM2Ffn1IB03MUFVDCItEREXRo8StvJ26guiyAl4ZE9jM8cMQZSH37Ws12KdWOU83fllQpqPZqP
SC8Hy4zFT51hSh6sTGF+jjEFO4ud7Fv4N2BXc+7NkFxNe0rZiWDAN5hYvwdFaveivDX0AKyYYYlT
ziOHx0nH9SYTRUOlzqtjOULd9R17TCZZQbZg8+e6iIGaVO7zPsaBOxszWeRPnHsnd0umEMAPmvbr
2uk28Q91egExhg7zB8STLccdICNkwIwVKt0S2YMUeFys1gMge3E/7l9/TgxRhyFpo056APInlomr
0RrmKTMVUuRWVIvLf9sH9PJvHUqGqG6hLKhKkR+nPQwhJf1h78WF4lEo/9aJ7RnHFY7f6ovNrMHO
bt5cWXHfZXN8g1fPAwYpBZWzgJxMhsE/SzgzSo9uz38bmuneoPTitBIsu2bqwQx2UbkaMVSYIKxh
TF92PhOR9PMIQX6DLzxio4XQh0LPx1ANCGEf1TM5hzeHCqsD3nm1JgEDUAy8gt0zdzRyGbpEM8a8
FwVVbzCe29z6+zWqRdauTq8jy1jHuCzuVYfEBunrq85PUaRkAqiUIbDztSnxZWcg5VZQL35/hieh
ZT2D68UsJBrnbjbpuTdWvETUSHN+liJ0XjJ8GGOXF1Iq/A1y8TgQLScD1uxvC7bo5bk52kKN/lAO
5dwIJR7Rvf3gJxnzDbVQjXDS18ZRm3zsMvONS+BxqRFpYpIniFuU/Y0SszNH60FvofN1FaQfaJPZ
S2CxMHjwPE/RnZCgnqnv+H/NiwYk+TGiakA2bEHMAz1YA2XMOhTS7+qyGEhhomttTzWTeXIsd3U7
wE1VRAvneEaSanAV1PXqAvNIexWBr0aAxLQKbx3olamFUG/F5rQn/oZioAxutZRMCdEQdvaZmWsi
MDypVCwDjSQRp1CQ2qJ8rPgooPPZeLOVvyMVm99Sqkf8mllBmJrQHZFdhGfoAePptjl/Tj/28dLu
lQtHIhsrKI9DTsaZY4lci5ILykjmBMxcBdggBKeoz4SnVOqX3JEtEu87tuvRNb5MGp/C7ely4jNU
MOVqj5zjhVyX6cR4Hp9HBsgJWjW6o+GzaF4H4Mmrpp+Rki6NgTKH2fh23Z5+zZqqjiADTrjYBatE
M8FOVyrvx4Zh6sVadZ5E4e9NUv1+1jUJbNlUjMhNN8lETdl9WxNiUmIbbtXafA+8+FTkhAWhdK8r
Pms8LpNkGIL7AzTPOSFYpb/EO2Y7P+FXtco8mgaqAH6ZqkVgu6K6sNqcTNu20vweJkMIiZnys3Yv
qKhmhJOCGl2QdhYFKUDwPpttDsmTsbGFlr2AC/u5BmEDiosIL0EMsuLJKe5yc1GwdREyqFDG2350
Sv/klredgacWg2azMVpiDeYh1zuuAPDHdRIqOY6Bt9n8RWZyw2uPrr5y6xYzqaayr9IgV/3gXei7
dLsh7zjEyNdrMnlCHF+hPq1av/8tXHEuqdAfGaGvu83KaJ2o2sqMdHpYrG22oCdkkNaRt+BkcmeT
6cbdqScp4ViDNLUYRW3yfgHaMC2o4NaWV9R/sYUlOrYj93RgptpG1wa+qvswzUbviQ9Epn5PnG0B
bh4lhHA3gDNqahinisCCd6f0lnaE/MQzaheq5S/9V24CcrvdAiAQ/S35GROKIgawNaK/xNt6P2kC
SjwzSxo1l07/DqTDRgM7AmFOtzW80HK5amDIcc4jOEo9UjKZntuPH3CgahNUIALIKlAg8HUudWma
EZ8xK28rCNcfMgPe/DW84b9XlYhTs5qkgf3j9oyN7WTuKvtbzklVEns91gCj3Mj8Y1wt54+o6c4b
PDfLVY2w5kol//mHGvmEcCjcRp0Ij131TVhkNk8e/Qix5TA4PJolt9l8x88nlZVaYZvWLLIXkoKt
AyuoRKlMMHnq64kCxQ4fNdVxDzIGMRgrHFnAdpJ78X+KMEC8ZFpja9qFGHfr6JfjxgiHIEI9h/WY
eJ/dB7tSQLvYg+1Zs11mmyh/+o3dQhz/yASb0cWr1AgDV3ksYqoJ3jN/7shUSJXtjnnpY4lCxNL/
xI1BdZFc9glWt2UPexXj+lzhPwAt0udYK52weFDhTSmsY85jMeBtbMA2Fe5S5yKA04oPnxQ1IfZC
0+XpRzHIW0pvF7L4k2B9bNf7kHVhwnoKjKpoCtRjCC13c57Ix3fm4knKuxuPtt5hb/ANrn/c0K3Q
iAlcy5VIgdCbasW+5Q+5yi3jP/ZHAToZQho6cS/XNgxzij/wB07R2It5uRml56ucMkndrYTIMXaR
iCyXLPvN7MEA9n2sfw96zAmdTeH6wQBaNnfZ4W2x1cYET2nV6sSdTn4fjj+b/Hc98MuxWuR5d8oM
j01bDbGwhM4CxzO+ylc4g7mYHuS8q3jK14u3gBB9a54QCU6YMzmuDZghEJcB8j+gut08xNcUVwM5
DhU2IOvxf1uXdu4VJIP0RG0OWy2OxEI0lPLnavNR4jP3tTlmgZIp3QF9SIGhoVAXiT7hbEP4t4c5
H6HeDzWCZED5C7DxVeVa5mnDPPpmBrCeaUXGbcTjeA9txCvfaEey7qtIEj1vYWWXFEfWHvD86sZm
Fvhl8Qe/cyuTp9aEwu2eaF8ck+GLp6y1Wxefo0NjO0R7z+QueAs3GDn74tmHmePl+LYoRSJhTYyb
E/YgB2BSrlaOXE68j3i8r7+ewwD2jI8yqRaFKsaPHKQxqeCyvUJE2yljeY2BYpcXwdpwLE5Bcq6P
mNddKTDB3UAcUvyuYP78ocVQ0GFieaPAsmOqdKv2HhIuOWUUJCUFW5SHqy8raGRJclIi4oguXBY2
QNfNaY/PjCMplbwsVcXDBucIWY1XU4xXTlogpQF6vG4mFto+EgXUHW4F0w2tfxBomhdmWzF4yuPZ
IIL/CYsxC5rinyjQgqYYKc1s5O/aV6/8Rkbdt9EjLV9DCnTDijJw38ppsXrLCOd5sZxvc50v8h21
f+23rhd7jA4NewL9sfLE4mwSaAl0I+7vS44+MnjqrPpGk3W0nwCyztHgdV12lPeEqgdTwp/Km8oP
mQycBTskowDjKAeTi0VgLlVFI82ZLQcW3B15otFoZy8qn57fpohGgl1XgFXxccVRQBnKN7CYNYA5
hu3fnwu2xuhw9710rae9esbumGlQIu5qaMN1HVlTb2rfAOAj/Keuwpfg7jnF/1bPzOkPbcY1Qqeh
yNU405tiIivHEEk3PbRs22kgAEpxXo4OYhX08pxA/0GK+l7sncrJDuM+eEgl1S/dVf+3mZsGAKvr
wh01q/L9Nvwb2JsQlPCDUTflJu34DAH0vD6tG6qWoeFVlQUmoix5p1ZpmfRcwAPVUf/qbaajlBM0
hLNugUn1MYJypjueQ86Lt/TaXwDrKHz2HJNUF4bHKlCMnptkUGZVrfaI/amrMFqwXtVqFRa8wvfz
JXluu8WKLSmBHvRh9HPDfqPFTbFs+d9mh/gDCKEJZlWCvTLrgsjIr9uaszBRu89UdkACEDKa3e1U
NjuU59yGlsJ7w63xTLvuejyXJU0ynvmrnLKfMND8OgdFveKg9S6acyCnyGUhO5SQnjp7TVMy2GZ+
pLv9fGbFOsSLDe59Wk7cKhEWrkV7oKb1I90AMtLAa0GmC1XCexx9KINPWuvxjnoVK20f21YySPoE
nlEKlp7RkF3NrM7QkIBB3bbuOGaBf3pJ5OmNi6eA8oe5KX+XQoLCzQPYWwpmKRLffflU7yIk9ofh
JR67GqzXhOg3sJkep6bSuZrVwgxz13UcKpougbhbYoPzOtCehzuyrcLfuUY9SNDglo21NyXQWMe2
ft4thCH6350oNL92bOD/ZvLWBWvbdzJbKxf/qPeQb345D4OlVN1b0jLOd5pmzPldgjfoG+s6BPQx
CeO4aYoAMGIl5tfyWOoeZ9GpYVR9b+0Z17irsaAJDSEWe8+KRnnVBaYAIEAMezOz1+NpLXtex83e
OEd4V9/bwtsIe2mmmYlY2MKFkPBytAY5SENKYIDT6Z9I4j0uyTGC6miH7ifQUBuM/MPPZC2i45+B
h3nAed31PLhLNI/Y3b34QOYgQ9A0as0zFw78R87Z/ER7oKv4KosT6LeQXoVQ0Zdr7clGN/gSbWRW
ExfJcbGQ5dJvywHMGgE9hKc353NV4ke4hhuyLmskapUEWZCx0uJnmo9umlB9aVOjWXrn+FFEi3L0
vRcNIb7HeYH2+uM74SkFjvQCWY/JiKvjCKIUPhyRFL5uTqsP6V5xewou7zwk/rQpNPg+fKNZni9j
JjlJm3KgRU+0UrGkM2s1vTqb8CsmbHEQEc9KxQQRZ6oYsvypXaQzIhbagAvON2EyYRJZfVFgEovn
4wM83dzz2kNQd5hDynKzZ94IXwW3c39W4bWesXuOewow8DMH5FClTnBtGReqK90GohTIkqzdnsrN
0g1GtfvogbMcjURgxeZ6oJatyfk6RzIZmqiousQ9I1K6PWfDRiFmJUZvbcaQmrvb+ALEPADXQRbP
EOSnKdfg/yAEm1N7mXWKGdnJfe6a7hTT2QmD9om+shivbqkVeSmS+DuHalAWQbNd2niHScHPGQRH
yfI/9kMkgx99dJsL9EWNL0dfBPg+5QwQi+gZy3VQzRUDdM/ehpvNhiXlN7nJqRcbV/hqzoIqSMz3
LJ3dmVeYLJX3IvqwmKrz02QPp4WEapusDUkRGGGSLBvsVyTnyaXOAlMFhdnAUPsfn/NE71A3i4jD
jqF/4BoBYY05Zl+raLktmZd/b1i+UAVHjHW9KRG7LtLS8BY6iQQxWU08bMoZEvokgKp8dSZuNk3N
K5u3ru0fbKcTweI1Z9NxAaHIurDwBAqNeWHGN01GEi6baNWspMuXYkQR67mbvZW3K3LS+MQOKOjY
dYDhhkaAg6GFMQ4jRBX3X9vCynY9XCVFQCVo8NblkDCbcJlfL2ZS9QN07qEupfo26ArKCX5XG8Ry
EFvC9EHlEDwUsM51CYc2Dkk5auuBhH1P7kKZff5/lHUXEMmOxA56/cnk7yN3ZV2QhOmz+Jmi6/Hy
Bu2iL8+GSzPmN96biOcjctNjYmkf/bZu5vaS7vQYwB8o/ssLi3LoVavqc6iorJxxbWYEvTyS76bC
TSinH1bi+IB/c6d961PqhmWEn08f5EAf9RsdDB9sY5qeyGI7Cx1QOrNMmzYSxCsrbuVOBrSpJRs7
tuohNw34LeVEDUVfpPHp8FjME/tBhbAOU/+FdOeKAN+xpqB4C+D/7ZZ7YsBl2/ILLcnoXyd2ic8d
FwKGAK0HIBXrRHfL+3qQSMPO3k8gJ21zI4lJGOU8tQ2d2o49tO1N/FCUnV8l7kXGQYV6UtJzAMuu
XcN3atOT41Vh5IMMsnwiwPwRhZadhQDjEElymnk6OKT+PIRs2TlDbH1SUETJHiGD18kEzwUiQsDP
BMcfAbDmcgP9ozr5nnLGwKLPE4kq6/chvxatuzByJzk1OYLbSM9hyLpmjnc3TkHunOX6YvdA+FK7
9vNDRWwJNC6Y3FQ0W+PjXZL4G6gGgI6I/3W/Q1ExwcLBD1OH6CX8uQEnhfSR0bvP9He7d13V9sko
m+TJsY/afA6lmK/VMZTwiBzo5NqBkeuDw//M9FEsauQJb03605bIbjWKncjdrHxIl2iwT4OfFAec
gF6Po77FQsN68xm5sVlvcAbOSNfTkXrMflAr/hhPX7yT5/v6t3sOGk6+gkZtbB6BEmLuPRjFd9RI
IYSSCmTIWCta5WzAHNib00px4Gk0PIQw9YqseEYCKuqzHAfbo2mLVYJYWqcZ1et5K1S2C/VLctXt
Q4AKKQywinTXQyNYOvf1IxvXo3TYcGbh8mT72VMxjBT0l9/FfeG/rTJdcxnAIPyU4C6b92xKyaCu
g67qDdeeVwgIIvXjIlpCGXIEyET5nFgedjm/+p1oZVm+l+XbYEcg+BiGK1vMWuozCEBJT3wKr4dH
b/C0ystsubjGOzWLapKz4uW9MqdigCdM0YdymYTaATJ+NGY5Biw8Xz1XDAkhOStnLIwUly4VYkEb
cd4pmgzDMe8NuCBnls17joMDvbrpJcEdoGYFGtTf99nMc+AY+3fxgSiPg219+j21DfmyhVE24Dlt
zJuhFm8pt9XPXhVgcrjRvO/kTOM1EnXQFlSdp+yFCCt0e4kmHEHcJ+JWpPcwllsx6dp/S/MxXjEg
h8FA8G3W5uK0WzoU3Va1R7aXmxspcz4aNdmBHF7EVSeEsfs9v5BkJwmBcepCUcy0LX3LdriHJN+a
j+UNvDKyRGhhaDBv4V1miopjL0sDN+8fTyMLzLPh9yHxEZ6Q3JuXUDedGwFSS7RlAkE7d/DfjEWI
dWEpschEqjUyC6kRrkLyeknhQx9rNAk0decLWvT9tuKWS5Opuo6YjUGI4/Bqv3X5kxqvLldEcBD3
QRin6zfcw9gV4U4A9M+2fFSUBHpDPix0MeSjnFHcbjUNwaKyyptBGz+gGKRVV7aW43Xh4Iaq/ZF9
hfJIU9ePxX0EQtGyyCJP4Kt4WkseVPBMCFDWBZkTrGM6KBdqoh4M3BqHyQ2bsrhzQRegGoQN+ln2
qNY+yOkiJHf7DyNncPpmnTkyaVJK8kghWozG3n4l76k4j6JbzzmcXr0+DuyHutXlGAhAh37lIXFJ
5OgNC+n6dXDG8pOIZv2cwAd/EPTJpgFoXnooOL9tWsqhOnt37LXb6iqlIJV1OC3yfT0ALnI6AB4I
Bel+S+N+XE2gpFLKUJ0YC8hwLHB0L1ADnmuBvtDKf/LQDj8FRQ7CPXwgY5m3EOioRl+TReFlIj4q
3FSktCQZ4ajIJ3l1Pi6kwdpI/FYI3YXsiuOtJCSEGzV5J92hhHca0anNr7hqUxIiT0Ilu8u/NWYE
q1i0QEPOXUh81sCU3182ItsC4dKDK8xB9rahKWkggMpjSCXV48Gki6XatT/0G4or/I5+9PnQroqK
hf5webkhCEZmZddly3RhAz5f3Rcn4R5y2SeQaoJt5e9BaMd6wQU3YHK+n2yxEUyC4np3VwC8jZ4d
9d/+XBW0htLjet7+r7f5ttnYpg6niQDp0MA0A9TUb9IoTi5BJDBTUr4oZgntUClgopy4bFwD63hc
pan2nSbmEqgWVqXtc8MjnynrdUoPN2tOQMS39Be1TIqaHK36qPWF+ngGw8wt/NpvZbqYscglEMSg
jVUmvWcBtxLMCBYXwNR7uyzKIwfDiyn/YC/iWMHrBwVlT36Mj2umqLtp4HtaP6fmnF8nbW+S54Cr
/bUHTaVVZSDmeG9q6dGJwglDDrwhkPsz7g6hWgshFI5bhr/LcHgBvi1ORZI//2nq9dIRw9IWepOH
t0746bKc/ST76EUS/jJWYVAXuAxy3cMe+o5tDmInSGkg33Vh9GQOyUsQmuQXBEX+bPuwjFBMzulv
QPeXtvedNhi6nJaYuBueVU+eokfbZTGTBhmOkfEum404O0yby3i4xWEjbEmauk1waYIso4r3MI0u
OCi8NikGuQVzeGHAH/yDzbelAXVRv5xI4PDCDIN7Aafqs725Mz3ykwAtZtdAGoCzT5JMJdVul323
nMXjLT9305q4aiu5rZUnuJLHqDUmJZQIMXr/y9DAkIsL5ie+kUjdtdk9Ld81WiFTC519C0gRGobi
BylIvy3rJ37XQRGWnDewkBwXqkRDqgmXncu6OTCgJBBgDkEciaeDzhjYoPHILm6FWvUwmIt8epUS
gBDQu1kyEFQ2lW4KDqzPIrJOI3S9K2AQyrXhDjA5JpCAVLgc/dPBQz3ZRHY4jfVKs6XqQ3coeYx3
a31R80ni+o5dzEhRnbAIdm3oO7F9jQTdtd7P41i6D9EfZ+BiVkeA1xupl56SYkjIal6b3t6ak8vK
/AkNSE/tTnfWto38rJ4THZKemVFXfIBZAvjRqOYd9Av0Ux9S8dgfukMcCuPNa6JO9Nnrc9DresjH
GUbcPLKYVVtP+IJb3ME2HacN+8y+nkiRmqTxXqCAuE7o+7dmnjsas9tawf3HEVuOtlQ9HRBXlg3F
HJY03aQZJKFQGJsNvD7uimOHLs/fgdgne65IiCmTvuk/Fr9n8I9gUvD1wqMpcEpZ01mqc9YqzZlC
OrHca3K4T3YVndFzMubujp/ku3zv5EsEszlDKq6BV4WPNVSSHit9iLz8Qxlv2PEVLuBA7431XryK
/4qYVuCoYujfzAvlMknIlR43gjrNRi+RwrpkpydvNvSWKAChWMtDxekJK4cfjkxnM1Egim7J8krX
YMSioLx648m20BfO7FM54CXVc1/T3ubE8nUfMlwvAUBuMjIN/FCQOsxr9s8Oo5jrh8GFOVRKskRe
GsaDGHb0L6r2x90mi+K8peCmvPLelPaV4WX2FPNpTn5VEBxU2mR5w5xUB0xChMfo/iJYKUE0bs5C
EbeJwT4EmhVawLOEyDYxV4dxa5hjq1kwAyXMkYZ0y1DruH2+jNG6ychbLhm7qDgBz+xn40zhvTXY
WHhXAsVSr3bzfS7VIRtUzH+FMj2YPFmeR14Pc7LynpkH9/XDoWlG62feOIKFIPtcfki3cZMuQHNI
4X/m7Y8a6hfduTPpeKAGBOSl7XwBnojd6bJ/vFJnCPn0YXycJcN/hjjuPgMywZDXAQTM6xKP8Hjd
1aCWdnEN9JOmImPfFfrmnXfL9wefprpCiSk4HiFFyyUOG0SNZ90Wz8kxLbeVLrtHojUz17ytOMJJ
eMRICgdeTCoUai7UAKa8mlxmdLAriNzAZSeR+P592gqrAWP6uo01UYm8bPkjybG3M+sOgo8QeHJT
dEkVz5HGwjOPk5VZkFJ/BYk+kcHR8KKK1lYYNPka+OBLx4we7Z74G8PF+yp7GYgKOW/Bezps+DrO
1XMYBiRAGYVSynDjsZcX83WeQ07iWswhuwwbHMiI7nA86WzVAsFeTyNJbAcGumAZVMK/Z4hGKC6K
7tfpj84L6LZg37+9DP6LmLz+tKrkuf7oWsrL8jGd4AkPZaRf8tBJOKRH9B7gSFzur0eF45VagZk0
+gAYhLL5IoN1xmh61+S6INQwOUkoxJ1/5CGjDiHLdKPt9T9Ecv/Ld0sWhLzddwM85VYDLKFBFB8S
Iq7EGbrYGBzCkH6Jj6tOL4bLNQOHX5tvnHfr+zt6x5xVEdQ5XaJC2qyAtgAPYUYwV/DCNQOnD7Yl
IesCNZ7hjo0u974Mz1sw1BdJeUjN1POozj0FLy6F/QcMJBsXr4EoNB3FLCyOnpSJveTE8Y6XpXS4
aFi1SgJWhUBsHVeFkwcPS2gxAnxgNU5jMDKYL91cCF9gwJuR8lVZPftyZ3IGZlcFs+W7WP+oWnCq
O/fMnI6iPRIJxLTVUUNVnX3u3tTSvSzIGuGb0t6UGHXEMHu9tKAGgpiIgGaOF6ERWJZIegecebVp
U6Zqi2BKDlkBrhCuR6m0kysDLsteWrfJ44TVnl5vKrHRDOOG8Y29veA7cYVZLOIFAPVSD4EWGgSw
0m46sE2zT5W6YZpKovKEmvK+cDOr8zfn35wbf68fqW63GlJv+SgymfVH6cRGFdderDrbLPbblNvk
2B93tBniHAy1i5ypWxA5Jc/c/qEMH7NN/iYi6bZEsr2jqHpRWIUaPDB9EdPUhpcgecLVVrEPikjq
MVQ8F0fN1bKR9foSehYC8sk+dPEEs3KpJhQ0eDD2Lhya+I/eA0Y+wxUF9OfuQfrJM7hdlkMHAQwG
chjniaL1AszRLUUDLxzqsSuqo6RwPVwp3N5x/H8eOFiEELrz1WeFeuo0VjgRRvZIk0T4Z4/2llQd
nUFh0/BXyx2DEmBO1uSewjhLoKEeNzbuUXfaImS5XKMuWIv3QCFF9U2d8DyirTbolizR0idlWiFY
Md42DxSJMHjJbvYYYYKiBWZ7jluE13Xuqjg/rDHAqcE+nR/LNFhfG9BTebBitviBKX7G1kdH2E99
vSAuPOPrBpdBCCu53g7BSSa7vJXxfPmLROKA9cQ6FgyNGuz+j40gkRQPTeZaISVtTPp5k2pqAQNF
5eWQ2JDVxSCHGMfyvhoqlylx4SXN2J1fX0FkF76NHJGD7Z2+kqKhzzA6/JsRBN5yS2p3TpZdIzCr
132Eo6oI30bqn7eCgnkdVyTgHbHyEXV6C5HpGOg/hx0xO4QZ9eyBYnKDlziwqoQpWWm55MGDNNKz
90yIyEtieL9ZbD4vyv5QPFnn6cPg66UIgWUursO6IueEc0lq9sq8o2ojeFYJ+egrE+IDQoewVPL+
VfcQYtHZnDPTP48iebpB//0V4rmrrwvVGh6+tAK1m5Ah8j9+3p0PLVIGVy2d8+5EFcHuEYyjnN6z
OUOibnkrfngSnxV7p+Rwmtx8qy1zo1PWV65cUdY7taGHATWF4MZqclL4WzJd/MXSZkRm9NtLA6o1
lqz/NbIJutZs1F6tzrqnyikU2TbnBOoZunYP2NtvDa99QbtKhKWA8991lUUZGFZcKATNPNGLvuD2
F7i2wVRafdggOxYmchs1wCsc2oB2hay++ll58VnKgal1Cht2HO/KZ4TtnZO1rEJQ4Z4ylE61MN7p
YHDYIK9xTeb4+mXGvynn0ChQFF0wsGDr1hOhrkPtOgM69IbdIH3T6XyYzhTGFjXjuKLA5d0e8Y1Z
ynuvRbtIUcNBd3X61biAiqY5VcZEglhqMVdoZ5wscSZNH5DEIGb61cERkBD/RK9C4rnJZSFs6XKv
dn0WUJBjg5xVW8/Mn8YqSTzIFH6uZ07jbtZwI8TBIg+n7q/HGHgWRjy32/WqyXPO6mp4bSICg+gR
o1PTrimZGOfOmqktPxo5WNEaAAa4+Li5jN6FJzCohyBCji98aXgkhOoaQ2v7iW77NNDj9qMI1YOp
HYw37xGwDWNB+eH8OlryA47hg/l9zg8kH2hW0ybMpTrxvzk8Q8j7MhqpERS1s2wv1Xj4XE7nAmIH
bDwUPbHBd+Tp+LXGjOgMvdpLW3HNPaRl/hzv1kEQlKcYyPPd2xHWxKNH0it3PTc3GXGtbQwZIpW2
Mqxce/XATIcU8s03P6/Fim4GfSc3jqXNUdaiNLnjJlMBYExLJbAUC8V/OXvZhgMJ09T0eKZeb/CC
ygj/doQm8BDPS6OJcR2KPw3MrghleDZbSNbgAJsJF1zAugZlnUrkwlTBw+N557sRcg97k+sGYlvA
AgNbXve6WK9Qe5yZ9av4Qv7Au4ZkWBBR+VyAvuALNMvdZg6fpjPuoG652gyLm6d/0SYhK2gXI4rv
NsXaFZV8DWWV3ZJCRhlGsUvu2ICa1rlc6bXJJd0PxusNkV879O6MFGkTdgMGZXkLKaFFg1dJqKuD
MnYEe3+fD9o5QFPI7nNYYpmcvIzmkGeVay+Jvw1+oBdLRSQpq0WSwGImfiJzyuRj+C/2iRz/m6Gp
jd7cFAnx3SNIoIZNM/gfVNWWUTGDdjHTCdQWEgnOGoFgXNxSoSo61OCla0tWOEgok3RfjQBKIhxE
L4IxCofHSayd2F+dgUbo/UU8+ZJsj/cJi/OM1LbC27udNtlezMmNLyHRP+tpDi7IrOFE0RpyZdX0
1qlGVSdC7hSfZY0ZmmBHxVay2pJAoHSDuNRv7Dtjiort9c/kyeCxg/y2n4Clu+txfp5IGYhgt2NT
rnYzgYAFn4kWNul1PO0eh7DcauEVbjC3ZVHEEU/YXVQ+HsUvon/6hM8zwTBcDnzLWLFpPwFQNs6h
CesPMSUm1Pjmdj+e+McFUGogx2jJeSQXcQELCOxpYgB90S+TiTECZ6xgji94w4I+dprpWbS8T61b
GYbHlN1bayW9zuJuMppI5sbO78Pcm70TYk5LgfqCD0+8+TibmOerTQASiuRIpurJpJHfVdvSnu0O
ci+4YBF/pzcqVNOOGU4tyKPzcoR9WwweHOfj69no8sfNwj5gTJ66KPUcHQxua0ICskTwXrBWE7fl
51Ig8gCvWMMvSXNolbrvpJUzNCiQ3ZJHUYMWxauo0chepHMVL6cnhZfUR11XuxXhRiVu8mdZYVOF
i7gMawxrAWOAuDndr01Nn+0OpsQ3ppJE7N0IxXnyiuFPo+rEFtCawK2XxGgdRRD1h9FUerBwO932
ietRBV3z5X6umhJgfZrfrBEufnod2uyVLEZ0G8KSsZDg9meGM6hiWHS+TxwkuPFYXra1rmmJ+dVe
4C/BqDhILFgyqq8WGM63GsB0bKG0UL97mzdYeFnMbw/k/Yze51jGEalYdAt+iYKtne3K4X097Zw0
Lpj7oOq3n5H8FSkpr9kxuN1OHhcGkSmizaoBV8qLbNG+8K6Pk1Rk3hC/7Z7tsEqC6KHkHN5MMeB+
xfFisEDOgPEaNltvlgie4x+BEtiWleRwPLa/Kd7Iv7NQ5AYEcOW8zr5AZJD7XwViKS31jO6uDSAh
Gyagj9yTxciEpPzCioTMfn7Hqdx79QSPCSY5rXYPELTKiXPJ7gbjiPL+H+XUfot87PevN8jbWham
XP0cO8Wlo24rD6yH6lRZx5/R3GhCJdnrKoQU/GkJ9LGBkMeTwabq5BM8aOhlUpNBS4W1Nynt06aH
Pw/nwexufV0ccH1bEPdyEKANJvA4CE2ZQW1iOrW0FUgjARowVMOEIrwGAdlmEsrpAwt5LCpsX1Qn
NFxZHykeZD7F6k6cKEu9TITRDNmek5DzCoziEdcNGQB6JZQww5Rkwpafj9Xct9UIDkKwZAsweuA7
wQyLDtLPWCM5Q+5OY34wkdjkrj1p5b6k09KWzpKEwwBXj7NNmS2uyCQ6a08tC2GPDIddz292JrtK
986il9P7i38hrHSCyMvatr4Eu75/G5UL9AmfBww3B8mKAO9Tw5gEdy/AYuKMN5U7xKkuscGpmmdn
NLxTv0odkrYwyBokCshz7f+sTJ6kbt/QbQnD9Yj9a5rh1dLCCsP6kAXNAPREJPuJob37K7BU+B//
mM2b5yQlnJw8ueGMdlqMiqfQJ6nXMBp4nymTDJfEJQuP1sUb5OEmVVQSlAnyvfAVl5nNDJ03u/YS
fObgYgPCTMhX8YbNTZZk9QOnZhP9ksiDJorCNEGjC5LG5HOAbPb2VMTY02lwK9BZZeCA0uiJfKTN
wMu9BpeK305sgGul+O2tyKG6F3siuljFhxE3lXme7JSJd1oPU04+f85qdR3INosgj6wGOsswZ7C1
oHCCcCY5Ksns/AL+hawU5uluxobl4oVEfbpIYeIT2yGTmkcReN5ZTNZaDOFQmmJqaMgvUMrXNrO7
YOSTvSQ4dTkF6ixmK3Fxrx4KiRiLf21+QmKdVolfju9WUbXt38gWO9bMZoV8j1xskoChiEw/l7mT
t5mx1QOifwrKI+ekAln3hEA/ET7liqCaw1Qc4YX3T//Z79wDCwsTck4LsM+vsDct3C6xWViifaMZ
W37hTmc8sSKaw4A0VoIY1s8yEJ8/vZmgwLUaJ+z86aHhuohvfi2558don7KTxL1tk50wI/BA0qEZ
krObfQQpnbOUfhmUYDrhnhjUAIVzqrThubbjm2FkQG5yudTtl55VGfwqjjdVA+jipIimDO8ZTilB
3CkLfoz39ke6EjSs1NB/Id2R/A+fx7Hl7sfXslrZnTx0sp7tQjxVL56CbUjlLaOmOr43aYDsuRLY
7xF8NElVji6gqe+Vp2cZSQULPKbKBD5cBDlAucbqv4sw2aa0RtjTRKXSSwZJgudQy2wJnH2yBD1R
A+Q+MFqkJ6r33BnKEgM2RSMk0okmzLN2MP6IB+H0LqzkngBVN0tjH9ZTXTu0KPBhl/c86XOCx9gT
17FeyEl+rDfwxN6qfo2YxAwO5q/kDVDjtPiDstW/BtcgtPhHzTATn9xV61MD580T5lZ0/G0Q6IuP
kvFPkbLkGuZ8eGHaUlQ6nsRLaZ/25BWQPv21u3O2+tLVzcsvGJ05M9O+v10InOtIxFJS/TCPMgo4
o6N4L4sUEnjGaVrgHvXJehdfAwABNTx2S+KehS8QxwTvI0/PyKpeezY94wdTFzgutZTPyWx6tK9k
IIyOJst2W5nwitwzwGcpoU0DuG7YslkDWd/gnGYhJi4M6AEgD3Xuaj2qL4M9SB7sEEf1lN4cnABk
/gh/yqa9p9T4QOJ9+pghaWWow5u5otY54auObo+iHCrz7siNzNz+lxBBmcW+0s6X8G9xSl150ABm
ioTSSaGy/uxvthUTBZVyksxuVWVqkxa7nVdimaocMrYNiefET1N00Ik4lIzldilMFghzsGixdy7R
3IiG0ibCbsVAvXqnwPpnKyoLpVQE1LQmPMOsaq8K10n1H96hOUL4Sb8ZptHrV3jb/TzoKZeQWRpK
QpG2FufVl1eEV4ALovXwjb4MrousqOJAdiKSsb8pH2ezeUqn2SkDh7YXuhqTUwEq8YKcUWkaSGbz
8s89WqdllcYySpq/nIDwnTkILBmrP2/z+woFZOk/TnjRDoRLJ/Waz7ARDEi48wpFnYQKl3rpwiCZ
KuY5wvgfwlNJpcJ6CB4IYjTbjpv/Ifc2wnAmtTS5hKERJGR508C0xlA6ly27AX9QTf0ut32pr39A
BmRhacwCIVgs6MThTdVqeVIHzaOkYMSaXFPoYSuzkQyKW6K7mqeFHr1937Rqc3RvE3TChEv0Zkjy
zCyk0gOzIbqrVQh2EMBB4lXZ++JHs8VNBzDVLc60msCgFViO1jC/V99VkwK42rX6xbWYQCWNASR+
G53iBys3MkqvsmlxrZOycJaK3k3J3ctodPdTkF+uBGyNy9qJgvkWhhDLPJ+CPOHdGNS9wjFVMgy9
QZmKpY51jHNyv1boiGEEKeFv1wuw9Eu9DTazUYrCOJcWAJqzg1FSqKiBLYPYUCVvxlUVUtyxM5x5
Mpp2zzc4L8Vc9GKkKp8RkwH0crqOM8qAh2RQVK8fLXjc5DIHA2yLR1nXEc4NvGVtlbPasEIMORWv
26lALOU+eZW53HttFN3fZVaxNRpaXfIfIwBWDfQzgtzLJKPMWFrEf5xDcLaHJwyZwLUKqoEXWWhr
xEBBEcPuSMLEUyJDUcetbt0zbamqwkuev8ux6+KQHKLQ6FnAEmx9gbquds+yus/MV0qkipW2x5Ft
yd55iyZaQK6cLHG6Lq2w70EwKcHFi3WP5KAt3vnwgyYGFrx6Oaocb6rTy+ZaDtoVjJjbvO+d9xjG
uuLdx6u87nKh51/xpzdHOtnVt7vuTMO165i/bFK0HGxy/MKN3Sl6N1ZWZg8CgzYzJWl7HgQBjDOH
59+D2+uNBiflfdc8F9Myl0GWaNfyQsQ9v1XaNDXdBIaGXDIO1RnyH3f7eS89/Yz2yEn+c2GKy285
YKgokpyXeSgdFHCxn5I8GKSQB5QRf0aljSYOhY4TwtnmqDQ5myl9d8PGUToySLTTM8EZ5FTgChcR
y0+vJq8ueGTgzLy4tA6HxPsVT6xajhNMXXZogLFmv8DCT9plaNmnrAviB/gKulk3bjIiyGbtI++4
UjoYf9Iy+KDdDWLaRF5YZafJBUqabyQfB0ijArSIYHK7GQFvsgBU7qCdZ7PAz7rIXMb48AgBM63O
kTjgEL41idckcPPX1ZZ2Hi24/KIQiO8BEJvNSUpUz62VUGjq/wPiE5wTQv6F9Hb0+94/dU2iqPhZ
7evTCDZ7I0xAn1obvd/TUj0dzFoY7uxSnaJ0f0S59nBLyWi96akC0vg27yJMCTOxfJxqP8HnBf/p
MfqLzNYaH7bEDXA/Y/kWcnjvPqVYEuFkGMFhJHurBfzpUrg6vP4TgTITE5Sdkoa3CVhjsCobxYJ9
x1M6O+9I74vUum1Atg0em8+ikpieEOJoFs2ajRQiVZYH7g/18v4erYckpWroaCOTQH6gQnaOqfVN
hFlyT8YqFYOchtLAmIVYj+Y29QHOA6dxiSFI4bJiKiK6kmAMXa/AbZjMuRoTBqGmcQ9eo0Avcfdz
mJlx+W8hlIXITb+XgkLyAKEja3Iv5mfhjRlAVt9D8lYNPgVb8qDnEsxWNLgiQdysIpVXgZuSEAJW
ubxFe4N161F4g/Gjuboy0ulErLF3O9yAtrYD6jfhwxSxwucar/fpZkBBRQDJVf3V6pFQsQi7lkpE
S/VX2bfC9chc9ro/95SQFgFgmD0rcX7bZWFK8auZ4VJiVi20gjuEg0H+4cjpN209zryHUOtBX1KJ
Tw77P087ig0xB3zMgrkVxUECEHVRBwmBvf/52mCWLA0l2JLnpsdhlNwMlfXNNECgXRvHWI2CAnNZ
268jf0NCuw8T2MRxMoDm5EgQG6Tzv2x8ob1IiD04NUScXxHQz/jkChZ1L40qs0xO6u9qP/t3ufBq
NrW15IIFSMTAqLi6km1doKOJoDSFbyKF2j5O+T1Q4lST1wSyfCVAubauKfCv5xaR+9lqlAxTlwCB
mKPqsFq4ur+sGXkEaUeyRI4pCX0ViCk+fzDUYxITCVPz4jxxdKQoSSgDlDwPZ0Vc2Ouy/NhhTFxg
Xtp9Mo+IdhukJtb1HFX/R8c1GnVkf9ePUaRUpJ8RGAvrOle8s05yucdZeysyg7M6e53aFsXG9Kve
Hvj884YEOUe7Lby89EDoH4Ts6g2PajLYiSsl/X1sabFgCVMdCtKcsrSmTroRRrQfQt4s3d5cWdmq
rbFgMvZjeIz0MzqlZzaTQQMEVFKY1bvCsHbUH+ZFg/aDxzMJ5uCzDwRE8gOZ3ha6dHGiQIkcplYb
GwS0Uq6iDmsnOraDO2kio7Qg3ctbX2iom4LtG+Xug5bZgDa3scILuLpm1oRKPmSIWZP+rOBPtkmc
D5OZRJzwJyc2VCMNR4masnVl4yUZTKqQ+PIDeEfMOm3UEfUQhO48ueXm90xztgPmjrd/lehnhetB
erZBN7OSyt6ePO5iNjROMd72V+y5H19N9nECOTL9LVG2KZs3BL/lLF2b9NW8wA8H/RzvmkcNPNV0
GDLul7ZmQ4tPl7Jj0GwC/X4+ez965p1Ix/y/uY9vr3BI9AJvyYFDvjpxraBMxi+dZsmVqkHiH/1R
jU38Ba1AfaFV2yso4gRLg/DUx7rM0WG8F7msdmw5ZzkTQCYs6iOeBfPmTFJPQ5v+Pjj6XY1gwRCn
5gnb8F097OdYkwUCIyuSbrGjMBbfCDatLG8thnqUQDVj3K8RCEs9oDAYN4yS3yb+rhjNvW3C4Mbt
JfUxZw5N/McJtyMOCblNRO9GMUy9rk0QsEujheSrgn9dR1wGKh9yN8P5BqOwhO3PK8uKxyfGb9aY
tgcr3HxiKf2Uub8UPmtlqmTqBAlvhet/aKIlb+F/duKH2+AxgL32qeMsG3k0YyAr5amCFhckYD6N
DFxoF8WNZGFXCAnSsLkKUUqmoUgYVxRuieEGADsLO4TGKM/5pcxrfhqKpbUAAMxJB8FLbDB5izT5
AkB//vYOgLlw/nM9lX61U0IdlEx8GM4ugSXRdisGI7IwjOZEQ9qahARQnQsIK7xteFL0UtFIa87y
DLxdbl3QFjgEHmhWUjdoE6Rh1co+AbYUnbmvS44cAvVHVEsEQIncn3omsLU9zgzsRT52QeUkPEhC
nIsjSF2Ju+mE004d3GFzARDSA6Lrx8fXFtSzXq1+IotTkMod1p2ZLBvSvKtE+ks1dJqRZlSCM9e9
Pl2yDMrMfpFo1IiFEEYpQybOny2NfsvrWUMCTMchBJoGSkbpEizfQ29UEG37T8+qGAB8lT2tQGef
jIcITNnE9gUiduYaLC6OD54NVuP9koibydQZ53EeOHfOCgq+IsoewaBT8WEznoQ+QDxfgqfETlWw
BWYbAmdHdkIk7OjIUHH3S1e5H4AM5gSOSvcI1cxD38gVFbEWn0yirzAOd4N5DnfsGsZB/NkHoHA6
X0tL/uEHD7me22VCoRXs6fstEqSkxWZMKQcmtLMM1mbaJDM46P+ffCiIds40dPbQVw5yJNWN28P/
yHySSU85jcF7rGU367PV/5X7jdbE5KABpReDHgQUxoBdXwcqyu4ZjnrOayaQ6pytLymIyR2N+5Bj
/6T21UjYLM3XGUqRUkm0KcxWZD06qjNYZzZSCiMPkdH+B58AfwWHvqnA7B+4PrCrHA89vdDEIEKb
dZNUPz6Dz50V8MdEx+pBp/dEYpsBgmhOHlYqOy8qHCUQBQkgFGxubwKpB2zAV74mzFy+l/oiVqAb
OaaYdHib4A3S9fpMiv/xrW+bnr91Fuuwsh1NhcyW8DrKF8Y3eVCAW4GIaJeX6A7SFrAQ/VTL/XPr
sPmqk3TDWxSl7xTzUIZKaiGj40SctCEKCJb3s1k/9/PLPJz246bF3eM1j5+GPxxK5wD5dAyEEADt
lWNR3pPJdQTf3tgYfDzpv76PlyqE9amWnCh8kfDErvwinaUEyYMksv2NBOtm+ZGoHpgzv4eiMYz1
oPFhDBdEfZpIpHbjbVgcxyFPkdsDYWEiKv/sJOjXt066xNxclfHdSZRZ1CfL3hlJ+Rzs5hVI+4gi
0t2PPtzojZEPjAU2+/xO1oRMSBZ17acEWCnPwPrLfayJcStzv9hoUnNWVoNW6cLNZS5rMKSOGCwy
LAU9KMMuzvYenR9pjXTu/0daRMVc5u3lcE43PHtCiwwyUdepPQ7/mbFSjqDrTHV13+4D/Rz2nyrZ
ReslI6lJudCUhgd5gSNMNp/4OZ7JSRL0ETW14X/KbeT78rouK0wzftF2cpWVGsg9L3sMQBkA4QHT
aadU8XpW7e4RQSEgFPqSJO9d8+vJRxFZf0R/TEDBwlt8g/PGtWCj73/++5ag1H2lTr9rgCFqNzo2
YoNuLNoi+HUcEphlfjtD4iJ46d+1D8KkdSgj8BxuBkZnfu0mf8QYXcwhGUEanwfscY+iKbHkXb8W
RJHIRRNrdXU4v0/XheWVK4oK/9lDkv+juYnMNG9EcdX75NJiC8ZPlxIPE/1josli+cn68C4xZdzU
qr+9sXtINipsjY02LM0mb/tcNdNm3lYOMH/3CpqMlztCEO5b+qatCsVh+I30rYNJdOwsT9IjFRx/
5bhN1/FjKraGxjtsOHHZum6rbRu5dSrfdgJHYJGQUmwejiyX4hdZoVmRfL7aY9yD4sKcUjeTC+64
F+YF3orklzPr3eJevX2UyOjEcJjxKx6HAWE0mpcVw9zIhGMMHjpOUgtM+23EoWyft7Vq6rNrpHeT
EOKSD3+TG9QSeqKQbWFc5hW8EDljDEmqDSSObGx5hcZuZuHYFS+Sun7DTq7Y5V5CcGId8OZrW9CP
hKGqm7Ln3Dd9E6d2392ANi75aK+6li3ySuzR+/r3CxZLV8f+jqxbIjfO2w+wzjuOMvakp+n2o/aG
jK8yfyjml912VPHj70OaheC/5FJA1+vAsUaQ40pEhH4DKnjtd9YHYTKA7Vy3yxCdrWji6DBCEHSQ
fjNcqCu7pdw7d6+jR6RQf5GuyDcwdsren3tg2mnsKArat2Nuo7tv9BDVTJ8UYfu4STgLHtpxsLFW
biWHu5oDdIFrFSaSPMah3RYaVhIxBWSJv472epar139QphDBXYE7li6lZVgKZ/p57IQxm3kcbe6e
UG7dEI0wA8V0fp8N9sgG52VoHpNV/4J1AFbIypo0kl6jV3CVGZHxbJD0vE3Wb8aXcuhqV3a+DpHH
FCj67+GPCLUsNVpC4kfh4I9uhwJ16gDkhAfVddbicJnxScl2DwFkgaJ/oowOt7nYMzQAlV7NLMSE
nzpvzEZltbxRGu0JqDd8LsUb/LjXvpb6DYhk0VLxM9Z42PP936JSp1h3XCM54hf9rOXv1pDEjs5x
p694rc6pGC66D5M7pssqefrIlXdqdE0UYfIQdg9KJuV5ZTVRiB6+NClve+2wyE8Yk/HrXpCOxu6s
UrbpuF8WhW6QxfPMUz6UzOyT0yicXTuzs2TyuVGyLR0UWaKp+5WQLnpr+KV4htSec7GmrhVC4qtQ
lJxykbCkGCqhPFSg1NJxQbfTsYiF5TKk1q5BVBPlDg6Mn55nLwP1LFQXhfNR7MwqwK9m4chgydnV
3uGTyQNiz892qvz61y8J1FcOiiy22YHnek5fykA47WY6b4fWg1Wp+Ujkry/udxA1v9mztOwAfjCi
8JJnZJsLvJbaDVw1rf5yCDkj2/ur1zVFWrHz17Nkyheg+x1Z3h54d4OKpZq7KJw/DWDi7LQqvpVL
jEMqLI5CcBpzAXkoS21W7pl9Eevw7cmI6Y9HN9vAKbXFnAG+Tv7XbDMBxSqaUe20WmWYfOCByTPw
kftcrZ1noL3PUSC1Q6sabnEQqwejLNAzkGU/xZzz7cYWgfBU6QGGPVyTRgBPZq/ypDzb7O28L9OD
Yia4lAzd2XVo0wuIe6Rl0oQLQngL+QR90x//qTD6qTA0FO/v06mIU04OxwzZNVwwmtjezP72dLA5
rmeqBH16rcJpFiDtHUkvuZotpjqP4Y6Gw5n2oTDsefS1q7/NEyojdkDTU6loeEsEqzoWnh6SpwZJ
TNMSnr32r5VxT3zAFuM3ubMVc7IU5gfDaTe6uVXm3eBgQbrinHXvPRqAgS6HqvIU/HeBm/bfaGfb
ji0RRQE6299hgEMkaTdMqRTLhZCgfCeJaz/o7/4GPxzrPj8Osb5xKng5L8gCdah6l1movPc3iG1G
sZB+VPUTcdQLscC5yjie77n/EVR87YrHTXWg1fMLc+K2yow8akuY48voFyFkXIvpzn58AnODGEyE
FpN8B7x/K6gz7YPR0a/CHd7xSs8w/Vy98Wi/LDWJqgEoBJB1V927UUx0/cus2aRemjeDME0Uxh7w
TqATZoYN3CzTqlb0yFdUUM80/S6yI6ZRJhMsecC53Upkso4LO5094GQHfTqWYvepItgenq/9v8pi
QAqr71ymOb9AHUlqjXKyYJNl7sG/2nYgMiM5kzuna4MVczCFh4prEyFHJvX3f5ayblvz6R4iuQV3
u61PdY0pZQTrBwF9HFu2xIYfSRVPDsqcgBmxXODDHrWbkvOR5QhClXcFKicOIqXu9g/gO8vDSccS
IM5uWDXzdnGqO+idslOhEcGXBFn67gBk9BWnQRkAMvbgXafGgmFLNQnC/jGy6o9uxxDOxJLklepk
RU0EhKS0rnFTOwFWz/iVkkraHDjnkjRiWBduFIUtl0ZD1rL5BE9RBD4uRkvaRsU6Tcy8UIKJysGK
1LFbHlUzlSkvHe8+x9lNgQzVTQct8wik8qV2AEKsW6CQYkQo6zaojJTVVuhwp2+BP/Kueq/la00i
nvYRQ4hosgeQq6/g1/EGY08nu1a2Kx55zhn0HHJR1fwrkryHL0TdQBUty3LpXSgpvnKqbFKho50X
1kkN7fDWrU98+hRPzflat0fuFT7WThbOg7X8FWidpruWLfeEHrKq7U2/adW7deABhi53YY8Xt1XR
wkOhdDVwBu8xfGsUKe8q+bF7Bjz6n5IrwwsS1wG+q6dspHVWkWjRC4TETxa9r0bLC90VFuyr/T4M
OxY8Tq/8WAGYRtmcAj3dJh82FMIh2cZOFi6SYvJ2Y+n6/k2u6wV/f1CvC2x53VSjpwBLFTRcePkm
shfFmkDA5B3zbLuYV1iBk0FbVUbdbopFrfa5Fjr7C35avJ6VwzI4eH4kEPbxrG1IMgrq3aYRWL9S
TAw5L/X3ypCvNciNNpi3ITXKw2p/8GIPm6rKZJ5peG9Fpd7MXKwEP8MdaTZasKOG0s9fwNTwsN2i
wgWoPO1Eq80rNkHhq6zX9xg8/KimM1YzEqpAOm7G/gSHcPteVYRa6dgj/2unz3ZnyDoqNitpYjt9
P8CdvXZRfcvMy2vzVFflxcwKaHnZRg/9PKVWcfYFYA8R/8CMBXtMkdlA2WqzS7kiGP1klmm00SX0
A+yumEzh+tWUBtLZQCX0V4QZMWazUcbEGll1ulaN6T4IU0jN76O8f/lJ+4QfZFAiKbYMwgdFr15k
RWly1GUMq4h6arkzSoiMzN0fuVj0ZM2YQ4BQMyBv6xz0SqZ1sbaRPxh/kvBBR1CMhmJXASV6Y+Dp
oW4kXqwpucHVq5MYn28MOK1altK+POICXK/tCiNha56bpmI62mquXi9NLLMt9ZC0kzAjSRgvmm6M
HsGYYvJy4wGmxPif4NhsAK8SWJSINXuJ9UoS/AHn07OJASqbNoyaJnpea+6yUbqmsKatMos9Q8X1
qZiLoOASwKqYvsFA0dboMYP0hsrXxMz9KoRzq8s3K9DfIFY/X+/lo8CZqIe8VsvZS8wlRHxGAUIo
E6POwEk22tIvNRaSOFEJvbfcL1An2M6qQEBswGm6CYpQ4Zgb2e99mBEkuVBxmRNDSa9mOof6OvNL
HjaPXYpl0iPuAL2n9ywV/V0n7fydGd/nJvZ69HbtqxMe1pj2Gnaxx80nTWhNTFyEuykz4EIJwWZ9
enhmju5s0w7co8SzaLeCptmARHQqCXEgpJLYo4uXYqY/MfZbyceMbPoprZ8emmhVU31Hq6pw12RV
ShoeO7SiNhwfbkqCzqOO1dgEWJ38mfkDN3QYWPsCpACvMTJi7dF1BNjYmxt7P1YfNBkmx+l4zm16
48cBlK3qZ5ftMInHCswKbr7KGaJrm+gF5YnJLZ+nE+0lWsHGTYV9JkHRo+dcMH6WTNieMdDpV0OG
SvNYBJRTsrp+Q0nuJF3D2yW+J19BAIXxNUGpAzNBrm0fMCF93oERr8l/jWPDzpf1y7/Di4eiKofQ
spLBnboG/NN+CUKdL70kZxr4vVDS0MDi/KO7h08w+yx/b+Jauh2q2LI4PdG9QmPNKJaAF6sQyX+D
8HRvQ4ys/k3SkOS7lBQJLv/d4yEmqX/68AyEZKUetU6jYmwe9J0hSw7aTXIQB15uW2YFFxoJlctO
weKmXBpUewJ+hjFEzBEmNepfn8YHMCvzvhH3rj4F+htKzvsJ64pP1oVpCD27cuyYhvTbnJNvDdJL
qlkG9ucIz3XWf1lMEzXzmsJcADvhvfBIQJ7flhfaYW7hIYg+7Q4SvW/HlIW/gWx5y+Ewq6PTwJYy
qUXGMeannR+L6yuFGjEv26Bpp5RVUR/aeEDVQ7G4MwqguAv4bMUFhMBzLV3R9QIhxDjl2854LxEZ
rgnEuMkJfaDX1hkTe1WHCESmUSX1QQM9lm5t2+w8Cve+GNLF/luMn5jeBgjm8eRpTRuZvDVp2zww
sPv4yBunfFj83shNWpgg7rIOND9zSfMSojJYKGuU7jG4j7r/0EvhpV3YV32b8dWGn/d0swPWb0jm
03eJtTQKKxzAS+Ptq4+lZ5036eapkNw87AJcW+pEe3Q5/TssSlA+YmHrOEjs3WTirgmGC9clx7L3
LfV43Ra7DGHkSn+L0OZ99wdg7NueUr9rK1LgtIqbcykSkSylXdMmxGni7q6kTKqh/SsSZA3OfyDc
2+JaDaB6SUK1FwZxlD07nQ8Ly2z6Y1uWCybcKcbY1hdVVVY35sjYyWWE+cLFx5CQhaMZTjzJJzXn
dz8fo6YJGUs/C/yIgJmdjZkY8syqKgylMUX1f1kjbg+TUczyDTrEvFITxohnCzwOyDOSY/xjIVqq
lFeg73/RpTpLqlaFw8VpCEDNcI3dKCnJOXOw6G26tZmxebooJ02m+beXsvEO3nav4rBY6/NCyQMh
CbK+wwbWRzF9fRR0A++3CkEskM3CpouYpkNK7mMjM0sUq43mJM8qBxEMWdJKd2urau94ViiINg9V
w2wxNSbzEvGJjgYyo7pIy+yYDTD5HGVLQsroXPrTn+ZbIzjj2sVfIBhx9la8/AV4/EWWMH99OOIX
1rzPp/l9Q5fUttnHJg7MkHd2LdNzhPHMz61OG8Gkifja2HyQN9NwQOPGGuBI/M0d5Z3eAS4lIddN
c/hBuVl8Qo0xyE7yhx0c4BRUpdarm7NBAE8Mbo/WyHTix3KANk73w0LKUKNUO1mqaNUzmXyscFur
Iwcd3opINJRscuWnfhsKemvxa8YR4ywJV7J0DtxFCWhBJNnuSc767gAGOTUjega2cC/onNMdpRKv
XU+E0/KNl/Fvf1WP697kRZJJ9xoRqszMkRQf7j+4filjRZiEsvgZi+p7FTLrV83BlNKpE1UxvG9w
Es1J7PKBc9OByUrj6GBpF0wQNLvYNbZ7AaxzXo8jc+JB1qw7qynHKY8KXGTVEWdNRUc9PRTV68ba
nHZ9xQfR71Ek19+xxn07n6/wM/S+ax8Y/uWdSmTbLKCPuZdumzVVCECVp9c8BVJUhzuLwbzyn4sw
eOXXwSahm31o8EfXPrAxx0V0ftoIVZC0ClArTOdQdzhEBZTjkwdlQ0g0rbsNSI6ZDJfLZtaSD1c/
durfHjcA405Bd5tMGuV0NAIKewMmhhWjIci6oIUv/I0Nu2GRlCIR9LlUfbBQMi4TydH0RGhvqn+W
ssTJmIezro1eMflJuqen9V4HPMj+deuW6tn1U/5l4lYPLk74Nnzpugy1vINo55XS7f84qey3EN1H
P4EQBvnCl0GREai630cii7zfqt20ewwrWZ7sdB/OCN1Bv1TAH9LjGxdvYK81LzL+7g/x7f7OPL5S
0VDwpytmyR5H5LeLRtDaHoVzIYihtLRXUKUw/k5DRjxFV2x+hhu3llVhXHSgwaLDQI3Gp7rkw+dB
XQfvFeNM1kh27rBf7MFgwARJ1pmbD3PBOnKYCbtuBPJXDgrDUlPCr7ZnY9LnNr4q/AnAYZWhR1CW
LrZe6KpgNP1Vs4pthZPRDp/HOXHcvoFn2Rfl1shgglmJXj2Nc1a0tX7JtYqf9BJncnokvvgvu9vt
mTwjyTtVFBqrQUD/g8VjuqIGipdr7sHnQlgkLcKzESSOY8BHq25/kyOWwRY0gVLTG35LtimYf+bx
ar+TVDUAoBVt2ZNbmgx7i43rpvJ8hKQOInFJheKJfyVxXcqI4+HC7BJH3ZCLsF9d/pQhvtdNaANz
HeEPXrIX6K+seZhuRisn+Able7DyQK411hiXQ/ayBQ0pi3BrCRTE4giYmw5QZl2SkXT99eHPKW0w
tzsXdJ7y8mGh0EoiDJQKxeqGl/67jQzdxJMNlO0RM5IGEQOhgrVxg7761zk9EKC+22sdD2t38glG
6Npe16yyYECuo47gPj51miM74q9i7uDOb8C2384n9Dz2NYYxly8AyUfK+jdosrtAI5im0gi7FUBm
ti/vfq7bTx0Pm4i7AJJ878oOifFc73zWNeVMNtmD7oRC1Hl6QYf3pAJi74L6NwRgii3OOVG9VlJn
7Y5H9mhaJd+bRCFZ8X0gKv+RcbbnJJHDyYzhy0tF2/sJtdgea1Xftuo9kmcbLp2RTweiklfmCoyT
ZVM8LAJ6pgzJxsfgmGcYSdbXIxH0Ty/rURvqX4vSFWbwSUFECXD8piiMaAsvUMohks4gyyZDcx8o
xpx5tb+mPrCKH/h0BZ2GznQ3P9Zv9W1Gr2OIONZWXn+oDKtZoHqPHGeFsQ2wF5Ul+a2ZAhzLaSqp
VIIDLCubPGgLJyeytb/DuW+RZdVHQ44ngR3nlr/L5qj+6jTm0IDHLRScGmJWCtRgvdMAJq2EyIZm
Fbbcin8QJftgJfm5NQj5BxOCs+ApsEkOv8/ls26Oln6V/NrJrpWVQAM+BV+fcTQL8AXQSbV0LZYq
BzHDYcOZd6XVg0fVNBUpS6MxyRdQsQQGc5wnwWQho4BXVG4wkByjpHXGAcGLffOgTXNEIfDJvsWF
R3rBQJMe/PjGR+fHK6+XaWhqto5u9CHMO3ZLWQWTmizn9fuVRNJ2bemFnGD5kehi8wkjYJPndGgz
3fktg3HC+2EYfeE1D1AFmjgb5t0A3UuG572e+y82gcKkIeiaP5b6h3uS+eu0y4tTnIW6Lw+rDPQ8
Cn+uko/nonbuTTqIr6HC4Lqo+izc6OtpII53rv+9NsPf85Vk5L+IqW6DRfIS3fuLZglJ8gF4Yj4j
xmH5DqwWU8+KPZ0ZMCQnPPLFPr6mCGo7cgGH1AiySgoGN5FN3jVW31QDI3lGHNFqYizo40ttNRAk
Mpl5gGiQCBAdUIw4pUKpLLroT52dSmzWIqJ7lwEW5qx/KI5JyAuQsvOo9ntVNiJDVmfw55F+6wsN
JGMvjAeZSkd7tyIWwaXyo+i1fByoQldsvG7vOWN+L+4A9VDKIIg4V6MeBa7Rv83OVFLTv62hCxNP
BsDe3r/RgH1wFnsfMFfkr6DXNxolQMJRvUTkEPH9cCxIFcykQvqkbQM6r84hHfhMCuQ9SmgvsbaU
h8kpf3i9RJc08rBpsHEmK2BsDycByMtT5PLCSMTx6e4+5/FzKaW/TBoGAUAA23fAx4+lZKPGxGTT
bBisiP7RC3MjkhF+57/HH16H/SUOV1OaX1HnAplVzIgiRN6MGhehoS0BJ/LAikmfrBeApgeGl5C9
Os4r4BMCAw4iER9WvGFAZUXRMX+aMhvNPc3lNIq5vbQCUBjVxs4BVb1LcVOtXyK8bbWWQbOVv5uj
MGve98zwk4kgcLENjYAH32P0YLXk98GzuqIMBONHz9TWjWD25ruAo9Y13k7jqOkbTk/XPjtUkUfr
hRAWf4nUkEPvXAZD4e1SClGm7TCn8TTWQwEftFivZ0rxanewcVCnM2VjX979M9YVlb3jMcUNPT1o
3fpKonFdlQoP7cr1KR+NeUxLmMAOxXv4bc6mfzoGke4Jpktx+/DSKh3JZWmQvGj24P295HhzH0JB
p2bwMz/K4a98jTB20hKI3kNZLJdPEqtw1FWoY6iCfmsUOGVQfqhRN8H6vFCYZ0/LReMhPxjN1XLd
mOltAabqh+SgiW/wy0rC9Q023ROU3TUQoWJZpcxZrFtRWOvuaYGHFxxLVAPJkk72bBjPz7PPAvFT
Ip7AMCH5IoK1BJzT0YiXLSJqTM+XYR5oPFI2j9qnwnb97g+T8dcNW8JoPpnhurwewTFh2MceSk82
KtIjnsct2vre2drN83PX9zYEs2dxi6GN+607/DaE086+QWFM/tv3txhMo6bpza8Zrlk54mG9bJgn
g6tLxPdA8ZHBbRhj+CmK77SqozF+9Y8Q+wXYk04pT2eMm7DzWbP9EImXFR8DR7NC5qYvqDbamIhH
95HjjQ/m5mKkYe/9op/37n3bxY/erKxgAZPtM9RL+qxIXmAi0GA6gRfVovtkt5kPF/21FLZJ04v3
+Q9sHSL7+1xz3kfFNH92AzxxDNmnpe/pIzfsBrMGtCqfbh8yeraRr1V+JmaMxsDcTbq+mRL6NO0h
8SA3P8Bx0GcT/Ao6gNnBtv2tiQSIf204VWux41smPTGM25GHDOVMXugoc06AxQ6S9euTP7JVAAdm
EA4YqXA4zBribwwgIcW0t0DToo9BbAfRT3tIhwX8Eo7Uv8Wv6IZSgWUMj4jaoN521SW31ORyOCzR
vE1flWJzQvZRv0Gz0jc9JyLSQhKArsAOVBuYs9zGizstCy1rOTJBB9mgKCZQGQ+j7V1lJeAB4wa0
gTiBPqZ+x1Q6VaeTK1VNXt/NFVHfpWN4bg94xWDnSZrULb5zKIeACSzIi7R9s/lo8sTSdQaDDwVi
dAQHAmWpGIlpCyqYiaQmlm2rZxx8k7+RZdlZoX/QisNwqHvvf0WGdciaUrgbEYaCQRMh1IY5Mi9Z
KyH9aDw2253H+30bILTsfuJ8ImxqaJblqlIyq2MSJuld7Td22OpbK1qfZr5c4ktJ3CGvgpmYU+Ml
2JgTyLAXpu6XR+OXlNwaTwdbIkbshOqeKFx/8YeMuHVgwUlMIObbTJ36QttwSZD6rsV+LE4ZeeEr
7NpDYyJfLnBnI2SQxB49guNMPuYKQxoERiGVKlN5qNzdmAGgCwuSuDfGD5FVSZ1daDah2sB8Ctdy
TDE01MdWtRPbXYVANhmfTN7ew2bTwUqdNoVSxbn70VPk6G0lhUSyQjhEp34l7vQHT6eEtJQTz4sw
SQmy4VhmA5acUmhFFuvtauoTdBMZcGpgI7NdagmVKc4Vw5zqUPce0aU+Z6VGE7zsX5HSXG7Dxz8X
+EQjcGvypHKO8JBhb2BNDva0Qrzz8U26ouyZiBTeN8bVhkNTejrHjAiBc62gAHBgRlXZsxZpAxSD
X8leyJg8Y6t/9+U1wepye7D/icD+hZ9TPxdGGzyDgGSKB6jQ8hxmvHR6pQQ7XNcj/2LhAO5vMfWU
emMD7iko7xMmPcVgBaObymvQ9bmeyOG4o3lCcuNKLwoWP07OInSFJk5ZXED2NYAsngO7Ng+1zvDB
k+2w5Q3wyTmd1lf5zVjHgUtY2LSd52QBeygziqx50w4i+vrgntJQM4sUvn5E2Blxlxho2Ylr8nIK
dRtHgWis2dmZJ1sPY2NtA+/1Zf4SO4nmEfGRc0Ia3Q4j0mSDqLl9CMFfDiAKeWHd27zxqk0acVNG
5GbSHWR/iN5OWJJlTHR5OlcdJdtSIudVcztKt9nRNUYOEuJ2to2MIu0rgYrnUsY+BbWpMhy/x73a
jv1fS3M7QXf728Nf2OEQLGpZILCzIEk+vGoNoA+njhztciHMCnXFOvb+4hb8ewU1oscy/X9JexTI
EErvYzZ5b6+dLP08CgLSUprpwFmmmSD6EVsIkP47nenQkAllT1X1/98qe+fbiPZ4w84GTWL/7S99
59n+nfRkMVA4zbHS0B1//5mfEPFZLhgmQ5tJ5ErcJqY8M/Djelxns1tDkVU3PwgaY5mf+NuwPNwk
mDfQSJWsVNK+JXS17Y9ZCTGxuMyAb2f0HYXuM7L/WP0ulunKYuRuE2iDPi97ZZ/bRClbUAg8wN7E
q+bCvKM7IMnC0TwKOcIpVowsvvgEG4kbhTzH8ioaOOszVBo2fQqNnJXnQIhoxgUsheDtdfpCztVv
Ad4oX5EOAGS8B52Rb04CGxCkvRhQRTPLWk73495cTFFjWAIo9N2YIWeie9kwMm/sWzInv5rkox9y
lajDLDpQIPflRDdaUsferv+B2ONpdpTObxvJ85Kv1B2Ui1HzmX/2+jie7u1IX7EFtx+3fHDm2N72
VMmn7PW8x6pPNlz/+T65rdHPqqxhLNkqzgv9WDNVX0OZ7dOeGVUcAv9V0Wr0cjVI4VRXWViSvysm
fvkcAztwvT422ylnpEbMc3hW4/vemwkfmGMoA/v9P/ezrim9Abc6yefNk+7HANNAvA79L0ZBzhNi
xznn4iYHctdGc+QhrIoy7y9s6bI2iZW21yd08KVgEBoHWEQsq2Fgh2SfZEo5D+vLUUr1NDagLU4O
d6Chb4Q+N0QOqc+1mmJEUMAYxurQKXFshhCDyvvkZjG7MBUMKZktjUtl+CyBQaqwA85s6iCFzxPu
rkDDATt1Q2ppNTzaRfjW7UjGPPoGw3TLJPlcgqVfrJQ23X5/74gpMy9JSZwuoNMoy+IUy/sH4xVq
Wz9JpKeTyjKtjNAQoCz1KxKN8DH4kTXFM4xVei21kcg8Mh950ZgH6W//hU2FCBG4DkYj1U4JeXJc
M2kFlWSAupCNsgn/p8fiypb6PLlirL+gJ4eo5i62yfjepVpA7D384/WUr/qskmG0zgjetHtCCfke
SIav5dBJgTP/2bs4ZMYw1VZ2JNletMkGHw56o83VMFz8WQvIp1nWmdUXvDrbk7R2mbHm2Xl8Mbua
jJE9dQyWRSY0mDZogZpGWtF1iufVlxTABVy2xaYuQKfT45LphSjgXUg6usBCHeGBUPFEWltpEWEO
Za9eu2uN2QNnYVln0jRwt+YfXrJneFSNDr+kwg1WF6CKxtWREB7qYRId53emCK69zGFwH/ar6LWy
PxkcnvxrZLaCp+pdnKImwMj68OoRMSVq/dGxs+OSEnfBFgjethTBygoZdD5kQ8fVu0SH9kUwkukJ
n8kQKvg/t0UDehMalWqa9pA+spQsZd6Na1Mq5IL8ZMYn0+fe/Am4j6U0GAmkCPMJrbXoTiazUFMg
0ZQLQUT47PU5hpp+yd+IP2ZIxKjkrO7o7REBu1+JM8WH2NigFUuDFAmf2RKMatdWvniQyFDMNZt2
Qd79gCrkyRqAgXWpAcurpzDxwp2zBRxypI+Re7jZeay1chXXxio1womPs5jvyANTXNXMCrDddDvP
Di2UMWl7XS+Cj1/4ZV9AA5n4yyAy+3ksZndO0+kTiVfiSN+1QiLS0Uec5opeodotSz49laxEqCVT
vCpZD0u5/ht9KVprRlmm0cxG/HQslH8b4/8qUnBA5U/TIYevoaZ+2GwPeg+Jby1WzxQYpgOZaolq
K2USP0uf1GbY3dDkqxzYqTySoQ1+31mjYBSdiynthmUGrwO0gvODrHkaku9vsvUa7cdW8PsEoh9d
+Czte9j25owjL7RWD326SyIdH7p+/2NnIz6oTBT2J3nxmIoViIWaYdw0tnmmmDJHq/5uwI0DK9q4
3MaVT2aWlUBJAWth5rKJDYd5fIrX7JVZvNtGEcadqPTXY7x3jjcpE/4mJtYScQdxgaXYooB3pEmf
+rWoPoXRBSqXYjOML163VeIlHtfi0Ms6gCk65piuxaGRCugQcO6NZhVrCs57tkFCotLbf4LcRDtP
EL5yT9w7mSpDHhP+98bGYCSjnLjU1AW6zWWLT5XXNm+EAF2IWsiGUXey4F1Dw3ZjFqZGEFIVbTqZ
C+VpRU7RONi91KoBWCK1eyHqlAdxaA0dJXWYFwcb99yfCtjlDPrk6/ZvUtEyqRaK+wGmMzpV0Mb1
MfWqCq/tjXuDZP9KTzh/f/vjFCAnWOf7U7eYwkjvRN42KyPqn9t5RImW/MkDccJ03yFbwWKBtiDk
jVe/F6zf+96DkPDO3WN8Op5QmtE/RSJePrqL8g36genK39mseUR2NgtYhTJLRg3ZbQ/olumlMlFw
pT70gv8asr+hD3ZnyYrRRT6K7cSib0wql6wsMEccg9kyexvSdy1rJ0rkyNbtGgufBg2IZCDQHC64
NBN/imv7hpJMHTn88MLwU0L5q5exm/QOCG+8Q/6yHmspU/YLaLIkgPYOPipSB/pGmPDUSJSoODCl
ZVzIALDN6h98sw2nFyuz7u3sWDkcEaj0jqsv/pTRafWzBaIqyIieHGLS/Czi5q2tIL8ubbXMKCEN
CUA7lj98fvOXCSHNmLYIAuCoS2ZCL49gn49zvQyankqth8HybKf06wkggdWsxjvNw/RzwSsJCwnp
xMvVN+laVOSPcnTAp1IVavXB6R5CE9gw7kUsz6ZP6h2H6eyA0FazCq+mOT8jcdW5sVZjXpsi5OJ8
qZbxB/kp15Q8D034iQrCniO1xpk1RglFroS9Ya9kjOiBD0Ghi03aUqEnYYacSQSDnnKmoUdRGLD0
ps9GQmA/njkuNePkWFss4GECsnSKBWY3FQ1KxD89C0pX90DZbDJpOidGGEvXbGhE1ACK96uk0sj2
I2Th8+8IN+EI2lPKwkp54ABczEz/ssbtDRhS2ASia+d3DpUAx8Sy6NW6zsZhGbV9svSpdGRv/NUJ
ViS+SaBA261duoI4H5ec/WRcgmSytzrXRdvTua6ZwLc3AZArBl/iXvIt13NC7L5VAM75EwIOmFcg
x79gF/hHhdWTenMqUU1zA4wBxmCtkE0AkkU/p8AkAyNnXUe56fML98oLr+J6xh+Crfbt4rcVg9KC
TE3+Hp2g1RZm+ZvC5Bf9SPYWVJdY4BbTOuNdjZWqQzCtQW+YM6voYGDu66isqzqotbNv7BFPQzTN
8Vc0QLn2ZAm4b7eLYh2kLEY+usnxPz/HaXke033KI6p94Z2OtfYXc+v72jVp2UcSQaQUqLLfeLNc
vTGTnzHkPK/NZ46UpKP7rNV8uyhf34ZvIssnlkiyWZhigxU/9aLeqwFesHcRbR0W4IqBRTMf8Pmr
BdlnB2TRikVdQIpr5TgaJe71KDrsaWQgNMN601p9aFNkvIo1N7ZQACNsMNfxrxUDL0xzq0gSTNtO
1ExDQaKMJ0Z3Y4VfaUSeP8g8VlijAwqpqfD5FJ6LCrX+pHGzoFPeoCn7QqiWi4iLD96lEWAajnVC
HUleZs3WXUr6JhHwYHjFbkAMA82PzDexqNR7zlrf504fJeeTjie9rrC7SO/yC/ljZ6NXU94IOMLD
bRCwCwZlrGCaYZOW3948B5zNR2HZXckJzn/KLdknqeI3k2L+W5zvucaF9pDsAL9pEvavq9egmmFp
ELeuYJGI9V0cH/8seI2LFrgIj70S9GTONZS3o+Z16LRQS7ZL9POr8wKRsE/gTFF8fh4ahpifqHiS
RH3wtKPvqH1RC+FBbKVMzDcncttOjCCA6rN3fmcZpMgXWmVOjyL2ADF3c2xix1/j96gFX0oxC9Lf
JXhReiRcYhrUZDzKfMEFBllqj+gwWqgon9CDpvqkVctuMqgwNaMWwsRumba2CFa5SkQfMk2CAa/p
KiodaM2uibEiCufqL18yzgiNCDYMlmVnttt8rMiv9PkJugP2U2wkEupd1b0uOYZDGsOGtwVbHS+C
9MzHfJcSkO4s1T7DOgzKBqO59EWuH0/Cb7U7QEaT5v5GupL5bVk+u3v4J0SR8h1hqRjJKXku/4Ra
h8aBWcD2xHL7UvZI6RGiXjp48+yGz2sVGVoevb2A1YlpQeOJdXG0AAJrAyENZPGz37HiiLH9Zw8g
xBuzA+2HJ+WlfnjIUeFTKP+SSFXK9RgWQdyLTvG59eXvF6USeJwaLPF/o7bmO5J82jwxWjbLzwuD
FpxhSbQOcAKfUcFa8CXeYrw3IyYosrAd+NfQDxYrN6rw7rt6Fj2yXqTeGEY057hq225cY6RB7gOK
PWRehHaKfogxGRfUdLoRR0LLt22eQ8raBv71vGtTRpJh0lATZAAlydnkZ6R9Nio5LEGBLt8MnbsE
+gLilJgYB+CuwFEHEg0yo8uNbKLttr1aPwqaOkozzerINXjXM1mEhc0SedABLKOt3RwrYcmsZHf4
+bdMdJ58neB+1vU8kwCMPjKVa4InCEk/k4TdiUUoi2zkQFdfr/DyeLzMtADaWqElAQKE2ImZlH5R
JPZzmt7JoGosIsnBTAOzDfjGQdZT0m6eqAGeFlcHoECjnrYzrFF9WOnSqhgQCdRhRxMhhjx++/U+
/pFDWXhsGG1Mi8QjeOj988W0Z46lxVSdt01wKxHL3k8mWVr2WD+AisPkXALqjQGJNh72fyrU4+pq
JkSd+v6niVJJMuvoG9D4DqGSO6HMqoMXqSi5RrotGLQA1bPeEC+1LKOR9cm4M3ka0jlcSmZKduvm
SCKvFx5dtfTY9KX6IxCp0uK0gWTdqdhd/iwigazEBQk3spHBlLzIZIW9eXchvee/IGQCTxY5R62g
I+OgUXGjkEQk5AoSzZx7GolvzTBWwN1yMXSm1l3EU+XuawNGpzT7ZpiLfIAE3GLbx4Jx2axIwsVn
i9n+pX4vActaaC+hlgQfxw5Z7TzglH94Tfvu7QtixmA8ViPrKg3vKUD7uPCTkqYHVGFHQKMeAPXB
4kK84UXjRi4EstFnmYRIZgr7mhm4hbD1ScEDOH4OgaY7CGOPvDcosBABtn79sfyCuwSZcNkOg93j
nrBPf5T8ONdzH5GXdLCYhzSFAKxBWZCrVs46to1T+h/7Ii37VgkHGXRyiahJf+EjPvE65XkCP5PW
xzvYhbkkMVrh4Okm1xtPhMhsYZn1TfsosQq+G+TBdUB9uP7KVHmkjO5ZGBBKZVXeyV43gHbpVZDD
hYUnm1OtXHGQOwFojN1426DSsHeyBrSgEMGhP4RWLANZeB1ByfHUEJZCQr1D1JPlSzFbTOd7r0sS
MoUe5KhI4CD72sx45peAPVqKwIMtII3s9sW+zdZBELWkTPkHT0k2lUixDLNnRgiwTEQRTFB9+Pk1
XhCchX3d5Z9xbcoQcW6miauG0hrhTDloU3gRhZ/CaBVcUpRAmAPJcVEBts9g2JhM+ExyuKQRvfZ8
tzNQ9R5QHZ0xSfAVB9WbVWS5unZ8wmdb22Be8xvUdHiOw/PFJgemNYPlQkUL1QsxfK+bseNJTuE3
BN9TUG77ljUuvnjx+7co+tUhQfxbZ4rw5YmtVWJ8tLx8U4Sy0kLSi/tF3AgT0uvUKS/oHCzAfKu1
lPAjkD/7JDmjy4/U+9a0jwdZ6LhpVDJkMC2bPpB4TyhTsrpzEyzVfJ+2qh0j7gl3WuYIvvZzxupv
xoqVYMMaUe22qKfmf/Ev70oMmhvk+57JTr56siKjr2vhEScpO93a0460NP832CS1VX/QYQfss90Q
H7RPwgQApCauWsEMYrNIuaPjC6bYOf9EFz7fU1eEq5pDt0kesd8hDXut43w1U6xNGYcRm4Bza+qT
U8lrknp3C3TIEbWHaAVQI6UoK6ig1BcBwypickKaOgAaEIM4JaUsUo2BOYVzVVAJly7uyMng1CUZ
dS3iT4/VozUW3hkXWGR3T3om1FPJHIBEDskllpNnuJ/px1FsfsvRtalhQ+TYFzdlt/feAvJ+a1TZ
ASWgKNMCeHMZG7lUwpBO+boTkScf6G9n2KkunDhyNTQC62bs2TL2kVK4pG9tyqsn+MpF273wzWZM
X/x1cfYQ7z33+XYanJhB9qV/maldOuCH/s0GZOo5aqWDl9Qw3BahM3DsaHR9KSZJFYXscrmb+s3S
acfhZEgjWTzC2eaz8ypt/ZPVLk3qCFRJM1xWyqPISoGgm8FZFtX83cUNhl8hLnYbVgyfuH1SXqSa
RYsGBMViv+Rs1Ft4JavmxQWLY0g0Ltn9PjzkdQoiXhI0FcFf8dNKU4HBs67JGIM2rDLDk6DeLXqL
HKvx7VrJ107B9WISOF6fIWAQ2KfhEPcG76sQBdLfz77JmfX4+t5LKXQc0uJ9JIB1ehOht/TW1io2
66RryBHJF0+z+NwAK9DhJ7paIZaBKswORT6N2hQOkgk9+tzGVjiq4j8DMHUJx+tCrijm3MJ+7E/1
sexkV1odSoM1fqEDno2SbPSfnhLH3KZoa6GHNIzO+7YEMXrMchhDTkNf56OlvmLmI8KSpWdfXzgx
VIbyRghCZYpzhFMs3pm1KxMs+MHPlUuk0Ynhstge8mOAUh1Acu4x0YdFVwF12S5hGw69IMvso69q
iNdkYXa2IaoHhm7hPywpA2zmJQ+YZqt+dcE6byBgQsLNeyciPMiMnnj6OE7AkKl0QmLvO7erw7EZ
/1vKjARhSotRpDPAKvHkWbWo56sWlcxgMX1qMLSDbY/2+KYoE7bMMYpTaVv+noRpY8DimyTFpI0v
IUYpRu/jTautxr2OPEQ/IyS5HVUtcVtiDzrOlgi7cGuBP4MkOAPGyimOn63HlJ0pQjoFvTFg/hE2
qP9ZQCsObgCixjFrrZYs0Cr5rP+Ut58Bw9o2WtvzKYkQR5lc8acbOCi9GCSS1VXM6CvzZoO/QwjU
fHh4cB646rbF2GwfxhqWQrG1+80RbKJDNGDZHgJwnr3YGZ3M07g/BjadOCR2nZ6OSZccdvkAv6ih
eVNJ249EgeJcUhqEqbZAAW/1JRcAEl0N6YX9ct3ytYYR9uY/ha2pIQ1DslB5AJ7e8AmTKCfg24iQ
w2Vk3RuKlK1Q+WpI46/LGIXE9Cx1fBcY19twofdO2F970jOFhjs0SeLdIYrwIb4+yKhs2v9ttlG6
qJZgIyypaTZ7/+O9X3xA0Pi9t7JcKBi0WAUtNQZ6VaSeQIqIjuoWHn1SD/d7qpdIzw1nSRGvL6Ac
RhZZBx/isBAeVCSToiqc9wFuNrtx7DIex79IRe5ZAj0W5VMawG1YhAEm/g4GK5xyS2ISM83/pAqT
ME6I0tDYB8zI3/JhawvRT56Vor07AK8HDFPW0fSJdDEVhQpCYc4iaFxsF/CXulk6iKlwOHuAaGyc
koFPHPOozt96xsPn3OWrO9IxLs4u8YzkWP0IlE8EbbveO0NOWjVPTc09INr/xZdlsBjhciqsABAk
dC9U3nzlWOrvPqBmb97u7YhrlaMV9vaif1IkEXx31wkMNYJeZ8WdCERqIUln/ofAHBCK5KhbohlI
GDG4HC04hAfCdjEpaLts3CqG3zqOKXQfW5agwM7lNz0BACyjdn6n+Q7SDPqTyWW6+Qu3l6YJxvhG
6q9qobot7qfO0Br4Bq7f+Fd/8XzEtRkt701E1iOgmh78VJPXahpQsUk+Fmq1vWIomM0zKIP53SEB
fwbIE2n/7r+hQ28fmgWV6hqOCwOtYakD4UhbaNVSHTXH4JvKAA0umyPZHMLf4i5oOSp6u1hcsy27
6mnk/C3v+SPfQOKcL868BmUfijmt4nq+5bNRDofaqZzs+Q3U6GQcPX2VBNM9ecqIeazPvzulqbIR
/1GE5CTVVeF9X5Q8AXXVcd2LmD0nOjh8DfenLUvkIOqzR3Xp2yMHsBA1RhAzZ+Qoda26bLtIXmmy
2W0IjrIZf8r3DRaSdKO8HMd/KwLfO0Lvn+AxhcPsf1mKUb7/w2/CXH46mhocW3K86attKHc0IsLD
gHiwfb/K8hQLN0ozaiN75jAbgsZDTwozdhurFKL8J6HSg/G5mgONHGPd7c7JLqA818f9zQqr1t+P
owRhjx2cB6g5aT++Q8w6Y6+4eapoIuWUzVpqBbRuv7gRq6/f0lVEPA7PCmS/TuTpi2r8/DkjHp7D
98obxlJksB+Qp4yM4zBM17EFZKd2VkHft+/8QRqVkImRU6jwSJ1jUhH/ZocbSrriUx5IRgCtmKSH
Gwo98Lgfloz8PxqyDhF5P7td0j+u1V+iB9HJ7jpFJeMmYoYZjWUAQMeTGwjOGfFl9tWvg+Du4l9z
By/PezdUcUVNog9eQ7eOtEgLLYs/vDfDMR3/3IEZCvBdpXROgu9OMp8GK61y5oIRMjmKFSnrQT6Z
kGos5xUwmybdFuNvPkpi6f4IipQin4gMVnd8sxvsJDIC6Y7WVNKze8wTbCRMTJVlEKq314vSVI0V
tDYEM6Sweq530dpFdjlNvAId4/EAiErx26d1Y+HBw6+RQ8IIk0RPdbQ4wyhTsYj10TNqJtEoD5+1
HLwyhSGbO658CDr/EIn9F5DaErPQXiwwNAuv9QUQAOnj8yf6eV3YyFXhU0OU37CDNOTZf3oJvymE
S4RkUpPe+Y7pIKruz96z149nvH06p8GQ+XAP3EpiQxMwork802qNm8LjpC+1JNxs1oKIKAHAaPkv
7U2jOTSvTe56fXU4IE5vHiZw3c/Ildc6usrtPoe7yQny9faQ0gcz0QEnhEKWZBKPWQc+ragPvksd
B6gsznT54TRbX3bBZ3stQ6WNUD+5EfY1hAh1rY8qKuyyIjflvTSHvazk9qIrVqS351kwWOHRYnPH
E3dXFG0NXwS7Yi60L42ZuVC03BWgyETvtGgYE7qq+Ov4NPKxy9P8rtsQ545MZrnXMxnsuF5j17MZ
a/JYNjFnFZ6GW5sjYRwapOt1MCYfhp6os9Rufuj01s7tHtlBmwiwFS474VA6vfecTc+AXqSibtQr
Vh1dQCzE9U3SaZv7KQGvt06OjQokwf4cbKGqu3qvYaFo8Iwnl0A5NESHwYspHkqf16PG0x+onxqW
+W8QxmXASa//GoEoF+0FtSBDgtB30eKXVkP0AS6envf4x71yKfNnlUOHB3pwigE4dN2dTEUvf6T1
BTC1BteInQhkszbZfvRvkg6RqaQbeF86mZIWkRFq9Nh7DUjqYvuVpGsExRbr8+2IgXJ7Gi7VdOYR
f4EE2Pe0ZFgHGciqADnZMLGNIQ2S4g+vGaN9/CsNqoSkkKBpax4ypgMR2yh8s8QsmHE/IW1HL8c+
+x0YsLz7JVIaW0TZKn27ChRqNikcxttu/fIOQh5U4eTSKNhr+BUpOIRGpYy/vMQnz6Q1yDNnJKY9
CNwWO7SbIoSMifE3/lUXD+52dM9UZF77FTj6Bro7xw9jlbXEgxsrkp2Z7rTXRYotTHnTyJkoguQ4
qfBUHzkhHuFXMBAQ9NWYv1/KDuTxN2oopY5dUHoYMqFAcWBGbWo/WJztVwk5PQfeu9S4e9Zr7ncJ
Mer9JCzAplmNYgKtGCrO0WtV3/yjs4pzZJYZ0vlXc27nlynCrxGkDbyMLL8KhpQLSpEpENN/pLW7
J4goiD29Tj4k00WPVLz0iIaQMUpzAQGDEcph2lloqhBtFJOI9cS1AE4dPHavZEnlRaRK0+3aOeXb
PG2IP/TodozxgM8X7zTohbj/ZefPlK65r1sX0+Br8FqqQkKdOpzcldhhYHdaCl/LjF8/Bv0LdvVo
lEJrkT1+YkswSylpRHRJAIPucfCV/Lj6RhRa6Sny789yEW4dps0bAnAhL3ERuJNP7bLURWyRRe73
VI4fO4ndn16lP/pGB1LW/J+kjKEuiXGpg5fOaN/7vaO3hqXWOGSB2IOuPviz+p6ChluPSPYZr01H
bshZgrn2BCebqbf62ebeDYp5IxSei6GITnrgS2TX5s4WyIFt+1tMPKmaA/0/HuoJ6+TSeg4Sx4IR
PdUsOVwAXsMswjnANfPOGz+IMRkBJTCVOAqWeCx+9qwutlBpcyZOVnuNusE7xbIc58Ox0FF/m98+
498OqtEAvrZOi/WQEbIejMdjSCdnmFKCROg5cm31gCFWnUHac7rqMbWQQO8fddWkmv8ZUbmt5P/B
gX/wccbzcf57Ayv3mxG8VysLELCeMsOJ6udmBfiZFllONgMG1y2TwRP3IbdqTIg8fXm+pOAtzPsC
ws0+tSgykdvDgBXMERRHflr9agIvOC4JJ5lZ8UZJUjvwfGXMA9MzAf+VsFxLYOKD8Ig1TqhqrycP
sme29eMbR6A8o6Pj2gFWcIXrN59aC92DGvsb6w674IZLPiJLUZM1rYGvSx1uIhqf4RSdPHXfrddi
LFIcBPbiQxq96trjLuZOkeLIzWvokY0bJxbK8O7G9qyDgROQHn4qZPflTb8Qmi+9W+RNzCTIa0wE
rmHphEWBXyW7O58X/dOqDoo9ok1ASM/GYwvzGHfcBs3FFVul2bagwG9TKHy5UnDnD5pBWwf9nMa0
6sac2g/LAFVIinhLsgexeDyODudP3tt/ipLc3POv1/0NzKMV1iI0eEevjoxo5AfJmvNgwB9WoOrS
/4b3tA5ZujCmLfjwjzEgbvUxvxQo6lfE/4bdrXZBg9MnPpwVt/cFcgG1AP5h2TDE0O4ZZAluCH31
OK8QKAavdSqAuRWBg+Xn1rU1V+pC6bOEEzL4oa2vA5O56+GAkJ3QmK0mX9KhQTEo7vmeh4nDwqfG
Ihc/QIjDbQF35eQUh/ae6XLurQg1hFeqdNtykmt8DpkctJqvpKPRmGHSpX3XyLr+PIXpkxX9l4/X
JJuuiC5tVJPoT7eaHh8U3X62vJucgPxC0fUw+RvGxQuNyrxXy7IqnS+2jasHBDxfFabuHgK/TX78
+i9wTUC6mvIavXmQEG6rUDJIDk3lClhVyAPWu2dBlOKyNbsU0aiIaBqJeo0E1zRj4b3zHdPX5uXL
QaZMFTyhSame3SwT9a+O2agGHQQ1kx0tx05etBiZfrOeQL9Ls1SFNpCTXpfVzYYPO8M+3Oo+cpVY
uMYLoo0UGkDUd1vXtqjv8nkA/GFr7FtFJgBrC5IRRusmGtjgD2YtCF2SkmSgI0EKtsa+y+wHl7Wi
v7O0m0SfL3XXZ+wHf0jsa/Y+9VzVe5PWWZJ8Nv7pY4kS7/M2Dx6Ey8bf/2CTa9la7qNk61gIW09A
zdfbZJZDRv1WN1SdpLRkHPGAAbN8ErT+hxR3aDQspVBM1vgICcQ4VfnJioiGytP1ZSsuCqagb8bB
SOf70JamHatgoZI0ZVnF0rbfRTOZqIsAZlR7hf44+zsdk5i08l0gZz+dYkSHub+rf17DYanKYRio
GKOKAgBgKqXKX8KKZqqgg0wGn2i2NzWfzj8/8bjrzmXn631NfuX1yByy/j52iUI0qW55HD/DZ4sE
FN9OGAx/FthW/1fz8RE966GYRBx5zzNzspjyu4DYNAWC6SRZSoL0+n4z/V0mCTJ4p7SIdwiBJ3tb
Gdt6iplAA00+B+9v1iXquFU0czgZEVGCISd68OyJeOS4WyPAPM/SL96aYYxJKPNeh1za4+ILCfFd
7ME5nf4FTh5Z4qiT0l0FnyWgRvrKPFPLej+f6FqbKtp7Yx7pku1kK2ciOb+qKn0ZUc4tjY1Z64Jo
2AiLbEVq1Q6jUBjeydGjPdWt86erNLQV9zajoc7abfja3AyQtgVUv1yjqVwXzMfMR9vsIRI7ScZj
LIiswFNMq3wIc/Dlb2y/+pF5e/qPWEIsvJo0id8CqmUd0lem2z5ieegcuWQE/FlUUSNrJ4KtqErv
La0JmI+JF318futtBu471qd7TKz4/8Bn0q16Ku5sbXfINMq17RW4n3ajqGH6Tpm8zZHk5Ow2inyH
DipKLKM8UstdkzR1UBQ8DS5XA4f7uenJ64uYMeFjynaFWOyf1cJNJuq2srjSZEl/VT87ggYLPr2U
5qwSfQOfUEPNeOtq+9TjitpP/nk6djMOrIqRPgEYrBXIAR6QiTCy56iuZ1zOJ6f/XfF5FsgNOFFr
/p0BVxdid9pbmQeGPU2qj2h7K/KDerV4xH9HmOGRc7Rby1R+Fx47Cj9K+YrqWIfQvRY0Udr7vUAj
gdcc1U064E8Ma+oQsugtCBfGm2gNaYEt/CJ/XwJKhNqsuEt+DaX5uzo+eUnlZl1gBy5YnnD1KY14
p9aTN114lcgjJPhXW5oU3BG+7p3mWbeU2L6k8pYi8UH26dX3A8Cq6LiCbS4SZT53lxuBj0xTRrEM
96WTFEZdRFYznqrLbh0fP3ufYn6JiWMjI1DiUYhanSVYaWTrR5BUtSHP+EcQKMEqT7rMVzI3G6+S
15ZGY5ICxHxE/HYEfFPL2DSanesEQRIZNMf+TzXxc8eZX0Ts/LnHMvfRE3yL4ZwFOjJXxM+eY76l
Z8RSBWSL1bQ2kOfzRMoY/yQvaxeHK9FiXH9g6Nv3OK2HPFRv8FFX/T4UlBINLDv2TSIXJUEQ/PTO
dTC4LJg563o3hUHakhBEXaYf6s2pKeU7j3M7eoc3GJDOJs5rKIJZKr+sP8cl8/UqHXzQPVvBAdUZ
6PwvAbEeDOxrBpy7NbKqbgo+gKgMGU+EIODV1Nelfb4PFhvFSQWlAuz7Cb84IBBhV0j/IregrFzw
aD+b5+GaIKvge65/F5gjPcDAubRpwd/cCfpuYAteEvtZryDDCq1lIU1qwGYKIx4gDHtUtSgpkzsm
q1NsGHqfsygPd7cn++wf+oimf2CwbFBoI5MZXncmAw7TkTYtdAMf9BplbnUWJ9SdFNS4M/VNkqH5
i+sMutTLwgolRN9jD/kKDLP5IrYndgAQ8dKpx6NR1gAzq4JWQ7u2eX6SahV5a5RARRWbNe9Z0ui7
pSvTTVs3tJmMH2FcUsx36YUuJFhJsU3+IBfYLyipn7eUb52t4aNm3yXNBlbtFUDURK0RlFh9r9k2
oJV45/Na9r6OfYxOUR+9rBO+KyQMe+nGCF6oFsDsEISLetTuYjclgdGv7Jq+jbyVDrWjeNoIKl8Y
eyknEsi/ZhdEh9HfcJxm7O610ioJe1xm8hSQJ2stizI/T+W54A7+ARVJgw1YT0sTvdbyROSYUa6v
1CJ6D87KrHeQlJlEU2luq52T3VjKhPyuPmn5m5UYYB62zlAot+kNqOJjR6IcQAnn/KFmBlcLkZvD
0s10Xe5IpyDti/tiQKr6qPPmcxswcAvZozNkY+5OMJ1C2Gsndu4NAIwoHHjCpVorcgojegvo3qgO
NI9LlslldCTskCBUf8YEWL4pUKJ4JO1JML17GJDfJTe9xuPSHKCts0nAB8/trcKQI7V1BRJqg9x2
vRAvLGVDLjrm+5V9cioMjL4GB2ZBtjn/Z77l9ZBbtf3/g/OGZe1ZZXxGTtjXyBb2C6jkLIAjP1av
piCSKbzDKHLHyxgggMObCrzbLu4ePHJjK8gIV7cz47Sx/8oIuz8n72je/ZS3lCvHWrBHth5N4KwP
ZKhq4i1gKxINF6Mjk0vxEeQZX8QNWva/1cI3e21iTV+FVqQN/Vw/1XrLLJD7uqPQYebfFUnpvMro
5/35NMYAHrRnIMDek9hEpkT61cVXpU7bp0MbmCGbCOs3aTfvryxqSGPz1rhJNt2CAdssF64Up/eT
WP0tYeN/TIanyUw9P1aALQLz/LbGhjrPLxXOM+Fp80WLni0SNV6yt8Ctn71eKHVPgrxzii8Z674M
nok9YWpOEAblFHLTbTbokt9DCZ7ODGR2r1FUUdMnYIMkbhS33k3dXJmOdcuPaHAnI6+C38POvWHI
sV5iTqYTNbZBzKWjgHxUPEpDrmdl3TOrW6Pt/zgymT2/Q8GL1RMFQ0occbXg42sPcgOcksWlWwwn
a8Q9P8A+TgkhlfGcpTpabtIgjrrGz//hH1cLi7/yEHKXf30bKJpzQ4f2cpuE3qW7/s3YWO7tkXoo
CsSLfY53rjK/4Q9v8/6QtHmC9SJSKUbVtSwIloK2Hoy5QW+qElzlBDO4JUr+ZylzsSRS08cQheVp
C4ZEVljFPzLq8Ju6KuqLKOc4rDQu3D29kLdngQ1orgW8uBNUQ+QXjxZdrIIijN5m6E15MD42k0o7
nI1zfpJYICTvdzBd6HaqrpVThVlGvxnHb4AH++8QI5hHqE90YEfPNx32Fa1exJSMtlmzM7AzUSrx
+RLrlE6ug80QuYo00sKCHh/+n/+ShGlqw/bTxqTXa2IoxkhLXdeQwQ3BRysCI/K+dWEOC/ipHOSw
wc68ozsorthBdhilLaVHDqoMeuPv9eZBNgOS1pxCsOUutzpmCAVC5DQGfOPq9hwYZHs8hBATEG1l
9QJPS7B81CHgPPO7NKcjBnJXJGBJNNKNnwGpLw3n2qG/gKX8n5+Q9NlT59OIzUiftQA484Kj8YdB
kUiuxP0uCEafMMrt6cJkog7G/B/sOKYB2geH8IlyBca0vAb4FxbUs0hhA85goWch+R05G+pXJ7xh
7XDeGXHvT2qxHYRcQdy6CgtmHJipNbIOb9EAx3dIUndRzgzCz8njiDov/wr759vbDpPM0HczdrmI
ECfyjPduprO4h+V/0rntD6pGjjbgDpIfgOWvqzdohDSjs1KfnnSPuH1iySLLv/uvHEOQPXBs38Q1
DXNtfjBaIk/jzFer8zY+yr0uvJh69plYCak/bC7NS9daAaqngkDjOonPnkKpxhJZkdPxylza2tzf
IH8SdbAH8zoK8IBYEszSAln4sVv7+Wq+XSOjZ7WqEBeLkWTBwGOstLSiKoBhMGLb4SBEulUwBIXM
0C/sazz8JeP8gRNxDAzoSfyFm+HKYLrkVb8D3C6SdS5DVl8ALFYDuc6RxUcfCu1sN5s7NA6ldpro
bTOvd8m2YwSkDJbcWzZ1PFtgiL1bQgR6FFv7CO249QLgb2BEkUoxlEEdO4Vyr95xK9ZpbLLrcWlI
br9VH2oA8rBJx3SEGbfmJnwYZw0b2Xw1uJ13QXzSObhQCLsbPKLHJr7gLBy91pzc5PuKJb5faANs
S+XyN/6Lt7iT/GvTcWmlUfyYc3X8vItUkYOU4mfHzR0JfcYBLuo0YaTxYsPPHP3vgoIYb6WOZz0N
8yP5z9uBefa07NWgaCaxr/FomAm1P8qna7aubtlCya15W2EH5VCXRMi6qk3c/t+ckCezub+2p5Hj
lQEjdhdbEM1OCrZBhyVUPDkWfkjjKTfEbgeeUQrZZ/XNlsdceL2ufn1mY4xzo0CbMBw5Jh1QuAu0
6R380bbHfEF31Gd+lDSPkgJZ8yEf6zJEJZLu/7nbB//4qgnmNioL//DevGc6mhYmfpP3OiHbHrH2
Ochb6hX5skq0kevJwzG9gQP0KH8GVPxypf/Kww/+2dP7s5hVRzt1HyFPVuBM46WzzR1PFE6zJQdT
FRPzGcDdsT8YK1Uaq9sew+Gr31pjGSrvAJUWImpKy0sv5G73u5KkSHelJKALIQVijzI1VdN4ZR19
I6ZKhbUPR2O30jAjpVu/lP4k+IBYAkZWiXse/01ik/feWEOrkUPlCfqK/6OL6gLerjPmqhEpQV8B
+b7a5lt/gcedriNnVkhRg8f2iRYJf3IPYMYl9Jk1vIZyLQ4bmQ1G9mnnbyXbCOKprNpc9S/+6YjV
V47pl3FmDDBJxH8EBmwfrz54tALjs80dULX4Yzn1kn6sLvJkT+gIipUHHIbWNHV/GJ2vmrHfrUmB
W5XD+9GG0s/OsIBId4aWQBe+l9PfzlCxBSYfhbuV/YUInuaaqt3xGL2fdpX7nHkElr0lqOzxlVQS
d3ak4KcA3Rik0oKZC+1m80VoHI4RWa5nkVKzeaAYm5/6U0pe5eOx03OqQfghCuMxE2eP+LO2hq9j
zWu4mGRew3hcYoucIURIkjq5EkfCZiqxTsjO2cSz1GFMqdC6HKAJ9rxD2tcc2+ymh/4kfzBUJ65y
rjV9x1EIkiu2+78RnninPGIwRIuwZbzdskHZMfkLy+P2chm2apM2PDG04qNZbb62C0KBpZ9vUybR
27UBZ2TGzGfrz6B5QEnsQNUmL2GSqzp6ga87/zkAN1PWuxMe5V+dbSZkBkDx4cwNkdSu3HbxkQMG
A/eswwcxm3NlbaI5bnznCl2KJK+cATZqQO8F8Q1NZzerF4mvLjgzatvYJeh2982G8bvBqtir1f4b
z9+xt5TDuISIvGG4c7Q3gAv95WsCAM93tKMyRyq2Dv23DQlsEX+OryZQfUD6IoJbyygZDhgQMkKo
ayW1O9y9H+EZSv7KcO8lFAuhw0GLwv2LZGvcibokRXYCIYKEGzY28K7YgTYZ+vdUC3FPBJtTlZ++
64DVGKP+QEhrE4WtNkOJMYG8nG/eCq7geEb2NEiP/30N/2heFQvMlPrdHh1S9a0gm1UaddjFegnU
n/TT53b6WM7zznnLYYw9QevDcdwLy+Av9ZFxk2z1tgzNsL9O4B77OYUnnP537Ak8SCsq4PFc0cn5
whFsXZDgfYeggQsEaTUOJb8H545uTCOyBLClUlbEf+ZPbO2qPsuo7Im4IvguAMtBZqUb+ueJtMQs
JQfVPhRXZHxLLJb/6qURVdHpVng7RsOGOU4Iz+vLlRj98gb00hxzSX4u7BX9E/ALWXLpBgiqTchf
H4QGO6tT7IIibDIequk3lGXjPR90/29enzzyswI2icFvwFm/zYR7YpXqLcWqCKYAl9UlNIxkrSgV
Su/dhYk7ByFWC56/TkdmwX4XGJrGkbmXWtdKnFGCzC0Ekvi2gJLDIjvRUwqni+yKK9uel7npJJuY
sOCOeHBC0KDTxNdEtuVGAglO/CEbNiXzIgOvcPT9yw7p+JNsf51Phat5vOzFACHZ/VA1AtqR7lgE
12rRWEvSNQF9++U3zBuyrZeG4c0LcUJSu5BlYw07XB6x6/R4BwuzciBQ7aN1mZBVsKKJRGkaVsvn
C8HZOX1afDVV0iVJX+gyksKFlBCdEIOdAWE28DyDFB8bdN+exrA9odZ4sKiUFI5wU6WEExAqCWXO
r1blYe6UyX0O6ovLFMHOFC3jOlq2pspMw3MWd4A/3fke6y2AgvQDOEeOnLz8MrXAmcmPo98oVSPk
Sb1MAI20gaJzWInr5KM/fEoFWGe6UcBVYcEwL5++ca44MBysSoS7hLycdNBv6d4q7HW8/e+aA4H+
j82ddEzbLdLdyF/jWvbvpbhyvjGPuDTFDY7d8CRblSdK/Vmhy5C08VqUXiemXW1fPpV3VIr2HibV
oYdbebZmxnBYvcOZZvvEy0DBp4u3K5l2MAyv6nBeg/VNRMzw/SXOYfEegeT6sFPZCSukPPVi6b1P
roD+vaM+D52CoPD3BdXGOYnvWyhTwQq79eTG1A9/2LUXQ32he0XJNi9a0r5qo6FbKvz8tLtYUOp4
RZTutA1QGDTRVRLTZlXFJ2xn8ani6SqMH+O2pr3OzRukPk7Rmhb4R7n38x6qS/9xqzaUqVOlQJUH
iGEjHXGre8djD9bIhhIJsf/iA6SrqvMDsALpmTuPtAEIZIXQDWBBJc1SS9i15Qf1fYT06Gkosfgt
Z9v57x1vtGMJQRa+8QK+JH9AHA1bqam9Kwv2d1aRHNd/sO+4/ueqizen1SoUyMnodL1wm89FyWtB
i3BYo9IAJCa7hv1yvROaa67wy5l4H2ZTC+OZr2l57LZNhcSh22vXhVNgct70SMosw4JomE6M0UsX
epkLk3cJhbqttKbqGn7cIC99XU85uhTVTDJYpGQ3qhb6yr7PHILgvR4E15gmYkP3BMFyrPHpdd41
Iqpw/CxpCwdJ091dnjAfK1R0TLwphPsVMSmC5bxueUfGKawZP7/2k5ST3oPcY28t2jC+FF3D2ZtI
kRjzbZUKVB2CadEchvuu9Y6WQGOP49UrMxBu4L4j3OU10VPvsq8+3kt5JfsgH4lTmCpzuweW7ebs
PgEursMYqamhUP7DbwjN9PMg/0dZsbxaA5L96HTTfLcp/Bp95cMSsf9tSJBpKXlmkuimyJBHkkVG
hCn3nN4YaHNBos58ZbzVLs7r2T8+FtpnPsrgv3astzC9PO+GXkJCYXXwRTQyvJFdyc/NF7qCnpw5
gw0bQ0U2Y7NfedJ8kjL04nSwl865AO+FepAlyeM4Is9HA0atyaN17M33xTY57TpfgJCzf6EDBE4T
Enpyhlznf00RuIekGK8MTNsQlnSc/GGOMRlJ2uLw6hurKIPMNVscq7Sc48cUC6+ynRg/ZE60EgkQ
FyhVeVRnQM1gO/6V2vjfUgPmS9XYT40QXgku7vT6J4q8xDFjXkdwBFAYBfdHeACabtd2tIxqbeOQ
sZlFBB8Jl1AM/+udCc64th+1dEucq4ZqRczfE9CPdKZ/eZlz9O0gkpLtiw5j99flkf4x1bDgFw90
tP2pDHh2QPyG77yzWrR8XtOUoH0s0PH8Vrqo5X0WcCy/kNd4fz9mYGb9+LnwsP/MzQuDnOdD0fJY
PVqGXCJeFwCjvD/HR5yemauHnMuZIYjg4Jv7cGk2KAzp3g3jKxVMA5tMiGt65ps+CzJw5oAKK2Ln
UkK4RyJiRG7gNb83dncFPurT4aRum4DqUlWBe8hLSVGcjrmQczuN5l2zmBOivSW5mXOK3EPMknOq
C5lhVrmx5sUf8WiS9MnnkNmFWbOrmyyisKqLjD3INui2SW/fbU44+34mf7mT87e6eIcZRVaPEsdt
fnySACnnZ0DzWhI6tMav0O9QJ5OCUb5XwXYq/mY8iYwi33pn+0LgqIlQAhoNu4Hmu4kHzWUHNqUK
FREMHZHBSS0V1UBXEOeaUi962jYyaMsfdHIbUtI9XpGUkNNx7FlHibiuxsUKSJUdK7MVXKxGQRRZ
qIeTxJL4E4mZ40ifhtVwvQ3gLxWMR/t4ZBLt3eQvboiAQ/j5p2INevLw2h9jje4Pq3TZbQ3Uoz5w
o72ewMkeioZSA44MVDoClRJeqyxmyBME3co/AjzE1LQ62lKo2DvXhxgZeSLwNPvWd+r6i06WLbAA
keBtj9Y5sn79O3rM+v7Dz5lkda+oIYb04KjpKuIpIILakfG4/yKdZuRh41VihbOPxJgK6RSXGJ0q
9eLocZOIwDsst3wsC5LM12j7SG20AH7Ir0PhxYZYbFVqU+3Pihqh7QiNlwxYFo7u3ES49V6bqk2g
roJmGZ7AtR7435c7r86srm2FE6/ROhv5eIjELXWBWfFvetjVt6yY0VvVkpu9R+AjlF+ZJxh8d2zK
hCbbyVR6P3JwPW5/Id3J/zCRL2tEWDupnuxMSDt8Rp7Mv94eq0dGajJiwz4zOOimyfdWzbAsXchI
Mk7BztQiFAL/zbjfPDwYWuKFq0lbPoNOgKfauHE5OCxEDXGe63JFzk8vLIOJ8A4us3vy3QdE03ol
lnqCMlJ5T8kT7y96/yUwspVh0WvCgrEEDzmAZNHAqw2P/arlr76pBgFtTEWVwkf/6+V68J8s9DwD
lP/yFliNc/6xjwrRyquHJmCb1Aa3ppJdKSORxhMMS3/jHWPBqWz+K5Ri61YvL5UxVfSPAoRLAZsd
rHNFORY9OlfuLWxiVNq0zMKjG7hipWkKCtNwVCKmRFwLuaaL5x/7PMG5y280uHNXB1Jw+VczqbNb
kSWIyAjg5X5Z/H38/6qnNrLXAx6C8nvuqouiW+3J2SfCfvYL9RjjpIry58SsmCtQG+mQ7UutlOyF
OQBxI8oVQ1uyAZ4D68N0+vEsuJKcZWfjsqbVFPoGSKI6NK3//X2mHOvG9M7oXYC7Xl8JY6tg4OJD
AZQUUPhONZZebtPxGXnvciYQpVyM07W9tPA1qijBQKS6ZHb6p692zobHW+JkSQaGm0TuMlRQ3Bc4
4kok28IWXE+t5IOAeGILoop/EU+3KBY2flB9xc39V1+mJlP8LpM2yP+TAQCCTf+W01ArlbDLrIA8
TA1u0qs7ehmWTnpHXxMWU7/5T4hqDmQK1ou5TPBruF5dzSPwkvz/X4Zdw3uqla81URb21AX8ZLHr
W1G7QITtngEaG1CXBfrwWOUHpJ6EoKadp9DmPp83VgtccCUi5yyYzmtz4P59eq+yjqRw+xxPE6wd
OVwTRocNwbxTGA7rrOuD6+R3Pq6GffVSysUye51mcyawWJkRR1CHMUkpieKBehHfAV8OA495y6Dn
HwfiuusOAazLJsz88koVGZ7Xc+77xgABasTFqZLLPS1jkP7zWY7ODYhndXOjzLml4Z1lDN34vbQQ
5K+sbloC82cOdbFrSmXjjNaAu/VlfyIcRhrYcNVfHgubiKGnmAIui9qHT+EyCvIV2FC+Q5dLxP7p
ai/uEthvcfDnHZflgAXAgkQwlQ1nLBP6gUhIU/p063qiKyTM0E+B6/F8P/+CmrKNC0uVM8TXQJ0l
hbEFw1l5UvzFdlGUFNw7F22dEjlnBOUAoadjhgqE2Q++II14nN8xhCsK7fxTBzpA7WgfHcYr7OVS
g7ZGJj/I4XT47kZ/apXhO4HWbj7wcXuGuQc0qbbnNq34sBgL6AhRrXIST5PxQSTYKBosXsXLqlTl
Sw1OMeQS9KdkoEN5L+jOmXyZO85pMjP/dmBGv0l/zgjLsNkz2o4abbP7VceFDTaGTFeESYpTGWQw
zOJ/krrnPAtQjCTXfFMwLD4zl2sSuY1JtAPqloSFnE1f1Xo5dhOf6W1LDEjEqQweRTJernqAs34m
3I+HlHGs4zyL63t1UXXjF6xQCaWsvWiTAx5e7dVXAKHVo5QwPKwTcUa+N+UEX2v6fWB4+HCtfFgN
CkDh30rzosfZa1tVvl7SJPwZVNOKfdEiaB2i8T7RL8sqUqr4Zg6p/MVWkyKVltSqDfNXCu4ST44k
BQg7pD0vGAr2LBqwFzlk/c7asi3xqzZpaGrszbVp9uYr2/TTEiZNReKfPNy/9YXwYhHW7U7fMlaK
Ys3UATbVCw4nk2j2DLDF+Oe5frAgK9iZKCGXrM853ZNgL0IxzRx8Is+xa9mnQ0Ks7/Klc4y2XrmW
fS4Nx46SKXHbcGTc2s3iS1XptU2NaX5C/IJHuKKiQCrbSNBIGO9vplFxgaQvgDYaV3fH3qdF46wk
peqdICx94WU/x8ksstfqRP46ra2jxmCTEZ3MBgnV684TfNYmw04UK3nNUbs20YNnZHetshl3MCbf
MWWqz8hA3NGYd9nlg9ksFjWK6bI5oD/ROApJWcQhte3rQtUh2o6d0zfOqWo/BgNgWGs3zsbxPW7e
S4Qnm15+mpcT8TOoInRm3k7MgYCn2gnrs51BsOn2Yr7Hw+EZ9c1gYck/5/SbP57XrjVEh4UuEbCw
LI2yf0rOnd66HtpY8CCBwQuzLOu59HD2rNGMYzeRzIP2qXeJRTrz/YoDOUZBmTpyauD264n8QW7O
QDAhmQXLWb28KgyU0ntym74vHVNfCnCAVrh3BF+PSUIVZ+msB3Z9SOgoDGQmEM7Mflyi2JOnw/8z
M+tW/3+AfWvykkAhmIcz8/ZjwPTzyAGxaF8xK5Di9/5eAyIfczMN46DT/LrR459CLBO1/C3WtA00
RpU9SdgyAIYPEfZbCDRxDG89cPaAeQbvh4ONdUC71Fqb3jZ2d9qfdUC2DtEEKdmDE18VYA8iXpGQ
2NM8hdgu9fGTLHUKRcFGJ205mvKXWsD1Q06YeRiS3TVcdjK/L5d4Cgx+XGcyVLQlpmzX5swy0vBE
aL0RIFYNvPU2W2bojG0jBbLWDpIf7pt7t9fz7YjVKVQv3/Cb3UlZEJgbtpb1hizulUdD8at4fQcf
7DQjIac44XIex+HnNFampKzZIhMqDS+v3Z+rdc1KAXpse6a7Slc6bbn1Q2T8++Y70frONsUoRXlK
ZzQEp2zgFQeLFf9M/sr+cxP5DnAvZql/F2m77DpUTt9tHnZQfOvV2fQxONx5p4DlRFACUwOarJC0
0Pl0I03R5HZLS8iTmONee3PGPneQOuLTSR/Re/yNIVmNDjSCR/vX+1AHBDEZAsjLpk3m7DUIgsvA
C58biwRB6IpD3Z13krp20fzEpnRNO64c5+KZwRfMLgb+hlxROAxDGbmnQsP0wXyLO8IlDaWFmAVQ
jYBcGM+6vuJgwZ6ecmFy2MrzMhf7g1kueteg0jF/FhOMS9n9N5/s5391rNyfuVf7v6DLEOvUjTme
3fHwFEX2ChNPm+YOI+FaXJxMywvdgbRtpCrjOi3rj/+7NPFOzaK5sDiVZHLvn+l1/2v9yLYSWThG
+g7C3YNFxEuuyXvxdNBOffvku69+WtoL/EcbGJKN+YxJX9UWWr4A8XLZ7419iUD0BkmqOkc53Vbb
sFId6iXHq0eulwC8ruoFo0PIxYv+r/O9GKpVEdDlSs3fjz05Ff/Q3oHbzqoxDI0+xVnm0gEC4t++
D3Jh0CbRwu1nkqhKvzHSQjaaVHi3m68SSIE61g/a6RdTfl+hFZBMS9idd/pJ50xFtAzPLnCifD4W
jA7VjN+Ctj4YwT8rnyqJOEGPlM0/T100cTYosYm6YHR448oFo+oq9aI6CSFSZmIg6WbhplIuEJOq
OkP/qBqJB+BXU190USkbwRRzEEGXa4D5mZe5E5XppggLalIlRczll018vTUgQG1nP6UKRxb0EEpz
WnHCD9SKxUdQdwkeWHo+a5ibRihw5GQLiPixndhlYpb55LNY/8NsfAPSlQZtH9qhiGh9b3qr7qpM
UkTYva9AXpCFzCYYr8cFsPthbcgydKg53RfSev1Jh+92vNUkMwK4wVqr5FJ2Gmv1v2LISzKlcAYu
/pAmlb4IGfHz7P0MGh+zZixM6pPbo8xin6RvtsflfcF2a+ntDKJJOESb/IgILdSHJxwe5AFdAhJC
Hc5qmbdz3rQMDv8wPDFDwh1zJtpKoH8Vh68+OD5MDMIf4xG/N0cI1laKD2rqb9CHPyQ8/xrt5VN3
elNev9IddsWjsdw5YxMDCAOnIzUrCLRqbtG9eIWn96IBvfXew7DoHQ/+nEIJmKlSVbQ0XR/jpm4T
IbZuKrg5XHsjMuH5jmqrNmoY0JokQRRPUPtgx3WKgTcQD93s4/9CXXki8v9hDOYGfU6DTmROjRG3
G3mIjTUUaM+N1rE4SPC+yyXfNDH9E1fVRznxQqzSJxTx34+n7D2sMSTDinaZMUNKMTnpKATzIZE1
/jhun31BXYX1zlriHt55WrqX+u3rUO9VC8LximNTOqy6w7Zz5Fo1nhVL1F7wcZyd/YYQJrMTocEW
VuwWQ61tZ4Q5LDI8VqzoSMrOPtF1K11L44hlf7qQoI27+QJFLItuJApWeW/lcSAuD9mTgrFxWcYz
BxWfHGeZWTqBzqNnpNPj0wzGbVmQ9JVRpMeVidI575X0m8yaInE3tTIRN6fjxY0CJwa7PWZfn+y6
sG9zj80JLMxZMQ6bYtxXVZpKif84TP2qNH/gLRHkCL8lXGB5+P0DMmkJ0lnaXaHPioh5RIBuOt8z
aT9xGBXouKY+P3zCv8VAoogmnCD3eH4if1ZcK5GBBTFMaG+PH9stIWLUff3PSt1RRDu0HndlC5UL
LLOVnA909zy8Z0xoDQQclq3d8+Hg5nie/blaGStpzLXBNVOTUplKt5BiwLn8ReR2gwi263ygJ92B
W77b4w6qb/X39k7h+Agm3dwTb/MZCe6RrIsqtpoGr+h/2OGEJazMx2j8bAPbmXZaItjaYVkIkaTB
E0/ptw/9PML9wQhLHhylh+njoEXWDJIyLn3b3dSkqOEXK80ECeb+D9cz39QnDqrKNwbbnGtAxDTm
Bb+LJjGE/QO0iyfBj1kdASIHT8Fxz+oEBzjJoiJLV/GqR8THFYLR/iVpBLI9iZA+CfryitOD0K6Z
a8GtF5VbfvFxTiDBldO2G+8o6X6uvlCKPehCrz+oVaWCmpSxX5bsGw89VP/VbRcyQnoMZn2Yk2Gv
ll88P2mqE/pydqu5KbHSZrjhPQ6sRsp8/PGU0ZjOKYyuUySNz+moyUdygucjR5QK1sm1DqDXg0t4
uUqy7fBnVa94N5LAykmlEnPhes9XRt2sSXPdr36MrRroCP6dy5ZCnpNMl/bAQCyoaDa4KVeo7dqX
GA9FIn2NS3MVaavu+sjNM1UAWK2K3yd141FxUDf3wPyTbDkeLH6dbttXMQMB17uf2b43lWhESBFt
kXMGunUYtLthKgqmjsTcNBVRclFLX1qL0qSyqbf+2WY5i02QLtCfxtB/UnPCIafpeE1ZG3q28Fdq
WrBEYBB/qliv5tu2XSQP0vUPpuq074iJ5NrTgIcyTOS3Z2l8q0+ZabFOA3FqPIhMs9kCo5NV92Ae
pR5hid2zMBwqHBi3jiV5aDqizdzorAIGaNw6Pw6MyywsLHBwYwJVNBTtt1KIgZaFEXwLaRZaBS3M
3jujWKQNa3HDGEL2cpJE9YcOMkBAJ54zDE+u+W9mARuz/JJ8tumL4HQJx9JxcPxY+wEG/VWqs8/B
J5q7+ErLYd4DcwBSPqHCXPWtdHaRju3HoqmavLECHDfbkT22+al2ixygb1emYLPM5Aj20VMhlQpu
K9wqNEbCJiBL/cP86CMOLf1ow6NJymC7aQzhC2OdXMCCG+VVaVqlO99RdorxTtE+j2Hd0Xv84KEA
0OtfMA2S/oAsO7jaOvdQqB0mgIijM98jZuPnO/V0lyKu28FE89B+rjbfBRm0GZ+KSNWYhdzPQ6t0
bB0+J+pFZ0TCb7FzMkziEKOFJjs/3hqqCb8Dp9o0FpBsqLGHjL45tugjRVIqnD6pMkg2G0yFfAoW
KRdGKjOfx3NX6WqDnrypEoKz3iuxs8j4Ga1L1iNcNXcmFDxJXfxULTeZsXgLDK+MaVkJguBEy/0h
IPxHAAk5pFB9e9K0CH/0y3ukXt6V82BeB9hFE00zn30Q/VNcRInjnfawe3HqkBXwvya0MEx4P0Pe
rPfhC4EyR97Kw1Cl7rDsU7w3Qj3l7BIxJDMYOEm2q39fSVdK7M/vgT8atAbwHQhoBSLEcCfqyxOQ
+/Beh024UCySkFhT/ONt760F8gfw4UnEbdmugEz8bQJ/9sqKaKASDayos864t3im/o6Vw5Zb0ouR
WgCfAjJeKGzPTg7HZIvG4yUOoi/Q0NG9C4WVQTG7T4eKbuJMsns4fSzXpGy3EOn8ieyb6Hvrv7OW
ue4GTfAmdnMUzhZk6h0Km0shNiBi2eksuxrmgZOCyCrfegMFYZ5km7+4EVAdzD4PsgsoratNcfZ+
xIi5cuSmAnrO5tgvSTJern+UXAE3+YQ4W5T2Sr4iP9w46kJORRLm6HN4KH8cql3VquhLKSxkOhEu
vVEiHLzRNrme0KE/2kd7shxVjCjBNesAMb2/IshWsHNY+ELSNhcBI4eceVpKq4/ldSvBQkMuJjw8
koXdIDVZYAan3yN8odrze/cMPELJaxzPVT8yulSfX8OPQ8mo/PsOYQ7LYVAYEFfJibo/y+7FC7iJ
8B8gKPWKS7sXaK6NfX6jD5xaPlKlZMA+7hK9REMun6nuTzTcyMGGu34U81rSQjFTbXsVBRzvAowH
Cc0s1kH0WqmpumYI2M2zuH0fRWBFPLLptneAo6Pft6KLOG4BN657epjMLj2SXKcd8kI59ppEi7hL
QtDNRS3spteJeB8vQKBGHVeiOySnIRG0pOYjhAtefI04Txn4gm0vG3RMgiTpp2wpCdXbhAGeAYw2
Njk9J6d/kV9NXizpt93x7wiPRueHNLwZmPeCOhyIXWzPyGW78cew+BvdZD9ncw55LQI5563/FCTH
j3agmWWRmdazKBmtsuWPtvKC6NsYJxx9bd7Ap5DUCZWMADffbz+nXPzvPv8yy9XDR/LJW1G5Cy40
+/CjaI/t/7E3IudjDiFNMDc7Bl4DylqGramw9h/ubw5q6AnLWnKsF4Qrzv6K8+rFLG28gV9x2+tm
SbRXXbB7Z2Z9UDwmbCG/A3Rvr4VhzM9AB62dEnSni2F0LQDWu4t1V7qMf4zFn59ZM3yhAw1BDJsN
zIWUIJ/DKKQLUaXqhqeSiGeQipLdYSc9eFkb0FQHEpANxbtpKGfZhIHYhwByvtlkkWfv2+O6lHD9
Ld/9MxDwI0hOVz8NyaBMtWr8TFoUczd/1Oqf0OLnPRLH2t7ksIc15JTsaDLLRwJ01iT8VK7Le7cB
RKaKQxJnH7wISTlzfUeyQkQfqMlbaongrzZOtVbHILwnM5UWzT0vG2XKfm8SWkIu9S1qcoCTJrZf
QAx3NyzIxovM+UQrHq2GSyqA6u+1v2Rh1ul0Gd/qukkYvPW0OY/eyP2q9kSBPY3iGcRbotXu3HDD
tJeNM9JW8N1eotQI/luk++KIVq55TJG71aXZTHUNlhlaM0EnczIqJNQyEnH3Z9K4EZqJPFHT3OKD
JyXlgJp7Uy0Zggodx9fQt2Ibq4w+UlM64JOQAu5NVQQVjTy1HjEwzEzc31lt68eM+FImLVraZqhl
E0GPKrqud8wS3yJE+uh3e1ofg7veHIjewWvYZNJbuQMfQNzkPNWCd9GDiUd6SDnLPuLlZ9tXSYlM
b646z+Fnv4Oztq9ccOFnuA3ZsuFuj9v/cEersaK23P74DsJE/dD+wavD2L1CGkSGYOgyA5l9NR7i
6rRLaaXC/I3mM9qP9QfCj1uvvT5/EVtHhEmhsUzxBmAafSTBWbiwYdZoQpXxrLC8Er2wzYf5dZLo
v49X9RIRdGi3Z1CWvEzieuMBkEKWoQBkSlReQ4CTQfs8o8omkXzWQ1GzaY3dK12FL+WF9nHkR4w8
8kAFtFTiOax7YqEDSrbfOqKK0b88h3DiJxHdF/FIgrmQB/3NDEDB2J/9+AKEexXBLAa1OfeC6y0e
qxiiM/vSyUREO3CDzLtehO7/N0Jbq/9qH1mx5SQIHyLvtLqTO7ouxLWx3v8xU3mpfPNPCwTR7Mae
H1v8a892LkQK4SWa1+c8J1UowYsrJ9LCDiaeCYOLd1UiDLqwXYHhPZ1VuQgcUqnmw4dJ5BYyWS46
aS8cIYbjWtai5TWSZrkQOGdPYDmklKBHWSobCRQQCu6+CEuOujXHP/9wtq/4Qb6UwYtOiwK+XtpR
/zk8Oat4uix+syiuppM25F/6GwnFXuHZ2NTBsRpv2kp5M+fCCIy61L1Eo+C9ZsYPxrENj2aaXhhA
+wUq+W+RwvEalkAyHm8xUQ27myzYyaCR+TxhHesarOL5q8oCE7Zet6RIaU0VRPRs8FmM/TU2Lv0+
TfcMWYxTJLjhi0YtJnx913Jgrkq38CpiPC0N4yaIPSKfMFGicD1K3Hb2RkdCY9xa2Y9wsFgsS8v8
YhH2N/250RqWE8TulrR5rj6T34o1FE+DTDAWjkeGN6rvZJM1rce+TsxeSl72mvevzM88oEISlz/d
QZ0ZycpNBWc5nodAVbUyt4m6wiMyeIF1zNlXJuWcCYIT9Uj+1PM1bPJOO4FiwGQtngUuBchobEGB
hVJAUhr8wtCS/yloRBHdeYQtx5kiSRn4JqmLdutsf08dklPdi+Q1Cx3re+sPUsdqkgX3LHhD1lGQ
0AieVfEgLjjw8YiS79HeTSZZENzlykDuxMpiIvSNucfOJ15JTrIlyLpQNnR/ulZ5KehcoNW8O7qk
9F9Lg7/+BDCrVQVImJcUS3jhzJ9+u/c4DiLBn6P6MckFw0z57FmyVJutd+TfjZP45EqST1H8Ecuq
Az83Rl/7dnH97K7Ugc2pKCTcsU60M7wkyiBEkq2iOrT3fnD9UjEy+UEGgYPz3FgyBjGYAGKLGDGr
kKQGdjv74T9TAhJe7HOn/hRaFs4B20uGkPBEMdCErRjoHIkaELRnfNdq/NARzj7GWWzRRvKH5vgV
8Z72Fp6wIyHHkg+Ur/5Jz2vjF3VAszudO0HZobeWDB1g4LXeleMvUu3sV57/bjxp8w8hYqSH2hPV
JaiEDIEJ1sytcsrVWzP+J0gXcj2uznc3p5CZhAcF+DD/f3+k13WKAbpP1/qCaIsn1vda+E1KFSoZ
Jd5xQH3qidQZyYPGnyTD25hfKOOZXJTElD9RTSca46KJtmtiwqYEaEF//F0U+7fJMH5GOG6KLaA9
FXq/hRvMWTSEll/D1X/wmdCDGD2qoyOV0vD5qfyTXjEAIoMxciqGUEStM3JChlajj81IHjjYXdFN
gpfslE2kvPOKDS6SRwtZVyza4+Ahr27WXWo2OR2FHYqhCeklJw2goOap0rumJm4x7QMBWqxgAN3O
c+PryiD8tZIeyK/BPHhZ3wqiXKfRr+l4PRiBEg+tQJvjjAp//VrW0tHZHyu0j/XHJHhYkg7tB3y0
PIXIIx35lunby/r/wIek4fQApAwKIfR8m/mYdfjoHWERYw4QLbSZRw/uID1mSzSnuLiBoX+Kq7FP
cLdKs03gl0BZGbSQLmANZVeHKf9ywofHW5rYG1ZVXaCvC9Xf4GGkjV3jqv9fM5D0AXNHnWqnlrIm
x2vES7CuDX6/sO5pMOI1w7Cv7jEeDzMlUet6fCnZMzeTIXbjcqNuqKWGqB4GszSSxHYfs8WMF6pT
W33nmBh7LpiZLatlrjnubB33tDuA9vuOFyDOmZQHPILkfs7YAkuJvxDiHFq1M83CwY3UCeI/GD3B
M0p64nmh6Zd6xWFHL68wFpLGhMQW3/STE7p1GI+Phcuq+379zHLL7lzhVePQQQKS/ADhPdTmrIns
bG4vYpxmKDDR4lBZd/y69a8ZIZr5vFZARQq6e2WTdjhE/+fiPSSyU1yh7RZsH+5/xbA0dCw6gM6v
RxuUZCrqO7CVbg6a+oS1Kpo6Bk2fyP2CZ8xNVTjHEhAiuouAEnsViUVd5ndO5Q1WjtG4FAdMqydo
rL/ybFgt4wR5Ni9h4w8aC6teJKIFq+U/1+Miyh+HtZz+GWUHC2w71o8rdtEX26nUVfuknS6NkYjd
D7isTEOBcCphNHqDDL2Ha0FwK9yzSO9rFCZHkymKBv032O5gKxwdpo8gOZQ59lt2xpMtLILz9mGi
eLM536ZptYF1MpRiO8RSZ2ekWB1N8FnzsQBgSQ0XxaEn1x29l9eBScDXc/axViNYxohXcbBuqGuR
TIJGDMPPI9sfOeNEQtYMPIboiElUzw6jdS+Si4OCJbUeqI+i3ZA9xhqz+uDqRx22HuXT91OPqI+2
UdwxmU0uUWAcZU1wX1uF9KynIgyFjvsbMwE+PtBu6vNQl1oe+HJH11a6Rx2FnYVtHWUC19OyGRJr
530HWz6s1xdFBGW3NajZfjd0BP675BQU0PNxwpgrq5zVqwWCkqDnC/kXLpB15j/lZrUSbEc+n5rn
ETVg7AAk/+QKsBTzZmPJfo2Q+ffYPFWJMorDPbgG4Ca1pmSP4HVFpXLymBG/aXEaICOAqlP4DEkP
OBN78rXV+2JqO2yVS/HQyt0q5/hS5XMZ/YCnG2OGtrvI++J8WDsBLG5w47TjbrLe9BYey9qQ0K5M
s+2KgP8qHvGx4o2m4/eQJ8kHyzx7CONdBfzrKRQJRDgGtbukwup8z04BD3HfxjvmgmU8iS6zAgDJ
djrYGR9cxgClhASVCckFSrbOpM01779TPA6SXKSRqv2kQp01ZMNOlLyrpGUUynvKq5HIt3ZFMzTw
BQZgLuZTQULgsCEW3MeIY+lYyQsELMelNSBjBSMhsgbq2L766qv+eWVdFxaZqs5aaJlnxHCMwxvR
7H47i7Rm0nb6g/y9sH8CUxj+Dea1ZiDXUJbYeGPoDHI/popNgC2EBBdHSNZMwxJ0bwuNn8qw4UfL
s/38rpBivBQSJcqSyr6FcXhBfEU0FIjba6DXxJ3e5FrtKvZp2vA7Pgks9dUSE+alVhJugWvYsLM2
Tf+l8C4OZ8YK8LVrJKJgQEdyAsEUA/W5KuzLh26R54uV5kH9h4s/7kgcCYAiLanRrdY2XlX6b8Eo
5lc1q0yZTWHWCU+3zuNmuKxL16TKQClS5zXiw0H6SIJbG5bOebDzBZZFSMdFLEl2TCfbQB9Tqzbt
2iFsw6tvZjCYoVdHppBe+btBiK9rnQ4lt5dzqE0Q8WA1L7mHfuq508g2p8rYYG/ogNT3QsZzXynk
srNybkTjhmeyvWdYkgCVpfWy0EjNjAlicJscSNMJSu8rFriLTOHTn+XQWG7c9XUg5DpiGrxMfFZB
hdnwxcW8+dynL8aGOXYEdTW7NWzqTqFh0db00QiNxW4yUanfeYjLqjeqPVztNFzps6k2BA7jczHE
99uUomZihiYUVHRnXJZR8XcjeTSi86N+urybqvHs3y1fYSE0zWvmkklpVFnox6HCAZbS8r0mB8pc
wfMFgMKRDzt38PQGBQFtDXkxmLGt8S9vFEx/kLsl0qElJL+uXX2gwMJY8I3LqPUdGNF2nsXaFddj
rLmCUJ5S+agMaP3pd2fNx0ZL7cMUSL3Td2L0QBU1xxoXSWCf60VD9N0V7WGRY2CAYsIn5SKd6f0X
JSWVFaqPjuQxAJGhNPMqAb5OuaNiwrRYtj6g3s1c4ED6asl7+kNoi3uvR5CFxMRuqrx7wYXpfeMS
9hwam1Ra91kh67lqt8Rr+iKxqGVvUXYWF1A4kf6Bxye5seBeQerlISMthuYPDOtvynioN51dTbSz
l2IuV9/aDTPz+j/QULMYaGWcPZCV538WaA0IngCndz9Q9dWpGmganb8xbooRWbabQAWjJ36PKJnC
N6+gGld7oKgtEqPJWOxtG5+XbTpOwEBTmZ4tBPIXGfLOsD+2lrZJM1GSdPYzEWJFaiYIHaeWRsXy
NXPGOqCw/L1SeueGq+pj4BDOqm4Ehynw4BDjo+v+i8khmKpMH9NyiexoSwMzjfm9Oj42K4JZVwts
7DfDiAz/OkrG67v1s+dvR5G8WWMvWr0Rs3ieuVaL2f4s3eYQefy3G3FSh3Sv3fMgU9wpSd/cqVeT
HMNTA70pYex3Z+c5PGwMpNRt9JeSqB8+l64yTf3PCYDhl81yx8Lepiy4MXQ3v/4qKaadZqreZCzC
tn05aazBWccOnGgOpNJrZvAkXgM1bm7zbAJeDXoDi1LBqDe8m2ZUxOpvGtyZDEFQrSYUTGRXQ+bK
T+HdFlFNvL9FmHXBLhcVvJKnHh9MRSKEtO1RNL6MnixFcDR7oDFR6rPYMll+94fMj+NGnp7m2Mbu
l0NEb3PSq0holitWanzF8RWpiIlu+P1pRkOqGr0LpajLZ4yIKp1LcMDiNg9ipHcCbzlen5Er8rtv
rZFSXGWwQ8lIKI0KXMs7H9PgVJKl1qV9wUj79nPKV1ZHg6YGj8ws0/aV0zDwmu8UZYDf9oE1OZG/
7ZNoC/GIUgZo9UGhRAtQUzvUK0LnojWONAXYnM7/pCc5lZAZkpzFh7uRvCGZe01HhY8OIMl42+03
0dEEs9ScPb8wL3m1iEfPONO0tFE554wAYVZBXWbDNYBdkxPleD6PrbcDuYZVPbN3hiXkFNBODvee
l6qLql15j5FrKXuz6k1uHcP1N+cCxyHdlQRTnumaYlTDKahTUlBZOtZH2q4XTbmR4w5h1/Pwv5wh
vi4MPWUkdd2WuwMG7PXZIqroEEYPYA3GAM5AZC8JqEdr0zHiDNpd3iro1j/UXV/xsCnki2IiWoAj
4MIIKXBxeG2RnTvEHZIZpQ+ZX/B0cKlXaWp+tX6n7HorajXTCrPithNkGBt4QlMVT49lWBFleHCr
dXEVtPDfu/k5Fn7QvT3yPs6C8kw2BxluF2aBS/PZf7L/xNicC/OfKR5UOBAyn7gkBGtU6z2y2CXv
PY9lj16hd9k+qhMxgwsDsWFfFB+Vjx6chIC5sZbNk2EdtN0xHrkBJd5wneugDN4CQyrDFdZ/uOH8
zs/6htBmFsWnKqwHpQGKF8uzntBKDpUkw8EUThzgSoDNM/4A2l5tIa8u/0J8A9sjVbcJSP1YSkb5
8QDSQbaz5WDKAyH23HLFb7cgGDAeFSNXB2xgWtBvRes/17gGHNsfKfZ0Qybf9bKfIYEeUUsWHcOd
1RJPqrYZmYZUMZF4+HJ2d6zux5ZzVzUxyVHAQwS2fvktRjB25lCyylUK7s5ZfWFmuAHxUZna5TZA
tAz1HaqBH0dZAEB1u8KDq9dLmEy+fEpdjK76xga/UVvY4St0CSogUGJMq7R71/Q4plzfZjBvPy2q
iqIjQhah2QzHEdqIlNGgZrTAaSJ6Xa4qvLUjcwPp6CI1wrY4xa/+1DGlQR12b2c3SCoAF5B+Wres
0EHGhWycXUdlV59E0GrfagCaI+D1tBcwldGrhYzG4uexH65WRJ8Zw3rDp6Zlrb4Ay0g71jShIXb8
B/wFVSbHLeCZhLZE3YDoTTZe7+qHpT1I7ARQWnCeTlejU44yG2m9k2MAlEweWRQmvQZdf/jbmJNW
f/oqnlQSOE7b6QpN69u5/BMdsNgu0kC/Jv9RQTCqSM/UdfiR9UV5hG//MNsitL+pspKCSIpHeMRz
1/v3X1p72cuDbgDECHJ1THfKV8rce/E0wpX+l3HyIVZXPGIPqimafV+I8mDfmcyQS50oCkoPe9vx
E/OptqlcobpzKYcG2wTAGmmNYI8+D8WFAZl++S2UoBwon/tyCUb6ka6aSVOP3OowjgTgDFL4eBNA
ber6eel3SLsrVXuCMfG9I16CWZotfWjPIvwFxs7n+xTkoIfEAkzRIgjfEjwr0+qS/zfGe5cF7Ilv
G0Ku+c1YlSSt8mEhs4ElSS7taz4/Uo0WXFiMGnVsFLYRg5SQ1lFjOSs0+dSjbUPWwxUpvMh42fVq
7X8TxU21sCgT1+XUyB3uc0f5HPQ/msYt9I7ipN2V5zMSnnYMQcehQLW0D7V1tWamJ6gDgoBhX99B
/VSMDBKeVXFYcF+I8PHp8VPdZPnrEY7aVUdfNKhTFy8XjdpaZsYMxegGAozngEnVev5DNlCgYA85
0AmR94fdQvnr37zw1qMCuhGzVio8fQuPn0AOu5uPpilFcaokI9Pia8Ik4CSpDdwPA4t7LFPwdSMu
kQLmEtYWp25zS1f4tcJjBPqNfTzxAV4LiKGmjDxAoeN7AQ40PHCPcF7TSDLSWGsec22I9d3+1Yfd
WIRwO9vgozR4VgSStbBRPA/YEM+If/r2nFXdC1pX1+lzU1pJwajszh4dBj0Zk6VnKOpgaIxj5wyr
SGoGfgLxI3l3z7DiYdrpuvYBQuwU6tNrAXQIdzTKLvlS3x8+gPUou4RgXpazTUCZ9zgLzQbhccPp
e7kfx/pl49Kpm86SiaI71HJObJBCuY3BesRlcoEYcCkzbZUY6LeubmW5Ta6uAREWR7rN3FG+3WSp
2sUF6J/QEnvy+rsSjjZ9k76pXXkwNysnKDJNO64Jk7miPx4EvA+M4NjotXibjxvB1biF94PoWZAR
IX8NOD2LmXmLaidGNr9y3Y+wcB21B2DT+W24r21owRyhB8tFXHccQtb3p+SuKJiNAAElNg62VyiD
zT8/ODDI+cx1LLXKQl1PNuIsuTMZjzuRqyKAnxkShxYNoBLnOVPihN2lYCRsLO3dVw+OjvZ3caSx
RyuoJ+ngq2fXPsSs+taFxPnZbBm6wn5o28jyOLxGZq/ggyKBAceNXcKbQnkG/N4vCmacrrYWo7ck
Vr5j6WnI+Gt9ndIMjM5c51sIPrX7LePkHxHY1IrrE5bhfM16Jb68KsD8HpFo3CGS77lSBxjuOC2Y
LvG2bkz1cIUYDkrQgPf99iD0fj9xXiLwdEyl/O9tDOvRTudi6rfUfK5m/lTPS4QPsbbvepVkioAy
WabS16QVvnN/6GGlEJ7fDIgettACNC1Rqng7dfjP+yyxC/1Gr/VnmUzF5oCWQ/k/qySs/hUt0SPS
w/k9L4Yj8xj+OGxzc6sxFpqqfPlvuY07E4MoCMafV1VD97M0QZKPJFedXzApZ1r3EynzQEYGQBqV
vLiRqNan+ko4iX7lR3ZGcnJmBXGPPR9W6OFYfRw6PjiC4RTMHN34xZoKBaL7reDkjXmUa6ZLNDLG
tOsqZnQbXGGgaNwgsz52Ve8Qc3CXyT81PiHQPn4Ov5SNTIW/Sjcjym4D2VA9Sa+Vpz9xiIEZsG6g
qVkae1hADxWMInuZRaLFEYIKeymDrbqs6RuBwKvxJ32fQnREO7b5gBnp5zA5eO9dsc7YsqaMiY56
v4lBsEFYE7TH/7kkt2HauOklCiZ8P/2kuz3k1QO3+A9+W71XwmrUXk7uGVxGmzAL5JFGayIB0fH6
9J3GD6/4S0oOd/e9pIi2SPoUC3udHxXGqyt+caoQh59JzlnDn7+EU48NcHLFLoveEGG3c/U5vdRY
NLzgtmGG364LCvTdCaX+uh84e1RD/I4UDrbdqYDSbs4bGT3QagpGij9DQqxEhNrKnurs8Jc3joX0
hilTMUImm26fKiQ7Y49id1l3t5FZfY5x1cHLe1PZlronxIkOnThstP2jZDbWwlG7YSOziBBhdMs0
Qor7CiQKtJlkuAEuoyfNua9NwkMdbwIq1Cdis4Pnb2YjTv1WuSZcSlFUc7N6O+eGX5AI0iNBmAja
0DoG9VwwZo95rjs9ukvOylA1bdYYBcKBIf1hUwctdXJx84DfzGFH4riMof3eWmqh23ksXLwKZiID
f8/a/n8eMgnPrcYG1M1jCMDo6Rh80MmcW5QGr63zgcnAoWB8doIfn7ueTw6NKAV2QbZxy56hgIGl
wfjDpMGo05GCrJnx0cu2uO54zxVNx/oHvvXELmG43oTq9xy96sl3zWOiSRfmc8K0jQhL4TpQs/Hc
C1C0SnYwlrXhbY121phOYEz/rlsbRrp4E857Ij6/RbCfCUp2MwBIhLeLNpG+qkDayFPY4ds+4Ur8
gOuZLamHxf6ACAReOHEItk+pkc2+aW4y+kpsTJGYwVTrHba6ddHK11Br72R2U2va8l2XlyKOOx7y
XzZUi8CLY2GeJj7LEfIrHueKcdILHzJVd/RmW1OQh9vZ3XjMgGugOwS7zUH3rQpIgJWQqohvEfG+
mdSStkhxpeRNxXsN8NmcmbLOqCePqi/m5XAK27eo2Qv6xmJ2p0BOuvtEN6IgU9gNODwOXNZhq3BR
ESZmjhjpyi4uXY2F/NeQ2WToirPMVH7OqPMWigLVMedP8mn5VXNauJ37XxedgmPdvx+qCLShzJlS
+Utb2Z746IIrrKaJKgwTOg3LHIWS7gqv7ruZysfn/+7jgrFO7GXLiUq3Pia+pugBlV3mrXLdsy4K
QV3oDMqycN+wYuK+B5vrlfwbEk9uo+AR4Swmn51eE5rZNY0xHZhdwizh1gfgbko+SXXIhWD7sGyx
JPlKGVazrJc6jbkCoucouB5euFdhvqAjAClD2lCGWal3+Q4nRFSVp6FzIDOLlg3LAejJ1kHGUJUl
AgECacPib2/8szO9xwiWLkLy62Yo8QMlgXL9E7hCGO3IKIwRW3FaduiGuIif09aSjs+4oIoB8ocL
h+EpFFPOXrHniP28/sOIouD2lSy3eJJbosjxv/fZj6ypa8mjE3xlGkR3MpYeA0qUxLZ7NlaVk4JE
PpCTJc81eWYFO5ZhgcfF00Vgx3mxR+N59BIONUQ/DOjQWS1i2jkYsBWdVdmOQx3t8jXu3W84k/Qq
qh/cU8xKnr4SRTECY6ol3M2B15OV/5+WiWbUJ6uQ/pPhcDBs6eiOlLr2gpDSYvP5HS4SWMKipIBn
xVKCd2OBnu5r7TC/yzuhu9sb05mp9xrLy2Y9hbcWlHCDtiHykD4czS5XrFM762z6y/lyUJy1rP1N
eUKpZ1HRTeGzaMdKZ9bORIuaVo/F2XoSD1MEGr1vCdv7u2flmj8hezTVQgzd10s3s0ZvGnkNvFv1
AxnTHc5Gv2nJLX/cx2jBTh44KwRs3GO+NIVA6gAFEG4eytr+6A2cUVgqXp9Phobwun6ajYpJEjwi
h89H7TrAohPLQ6XzqIx+MeGe1GKBaNxGymeAZdasWzwH+YHBX8Rqz6mDz9IJXBjpWKVKg53us+gy
xtUuFM3VRILw32qgGZrMfYWLQPLIvfcLNEjiGe3QpHaydknLH+7TB4gyJPxg6FN47uLYW/5RmgKX
SFlhAifjq9g3ER5lnuFbfF3BmnPOogp93at/ZLcOAzN1JAN4qX5hoi6CPfgtHZtvnTjOM+XylcVz
MeanIHLjMXy40sKbmDUDS4NtLAaK5ID19cx4uLI/80pufEWoTYfKjg9D+8gt8QiQO2BGMLhanCuJ
xKUZP0RF0+Q34j4DQaOPcorVkMqbKxbxIRvGvV2AEm206dVBTLA3zvtxS+x8ybG7Ao+1n+UjGvoQ
VrdtFvoEtuc65Uk9T7JK1DWuT0UMm6GOgoPk/9sygNSKxkMZIshejfKcyP9lE2qKbCt1iKBUuzOV
Qhm4zOiCcouvU0gfzuhM0Vk6Arzzm1aA16z6GkwduWELqlqB7fvVQrJSCYaT7XovOcWtBvs1i1QQ
02WBJGeNS/1+nnxmqNjif+o7obuk1gvtDJrcLXGORf9Mxc3yyjmTJCeqYckzah8KJo/xQE97AAg2
4U6k+x5yjDbhg2PPwIiC+CsRsmvSmzOgLCeQ+UgC23d0MmfM3mHLL+xKP8/8FpS3UdMNvtJa6M0u
bB9IXySq0ogc1u5Hmhrzd8tJ12GWHWhp55XkybW3aV8ji/u8fd0/jVfbKGnLA4yS6359phqHeM+n
MvAtZI9gnrvMUegkf0xDP8NyVWy1SscAs0wtPJb8/YYgmKg2y5YEO5kHS2J6V3/kkVhISB1G8esH
nYTJLSiJ2SBbdRdv6WEGWip0x5UgKrtpF1OCA3vqnV7k/IOx9mz0sL5kfb7YYhyb+YrPGclrynPa
RNKWALWS3dJycHnvH1+S0IVe2d48cTXHeRM5Aonvo5ENpvrUMJfaxX4lgYMmqy2VYsputX79SwBd
yENrb+zF06gyGHD1A9ma3Eov7s7oUA/Dxs+4R7yUvWOfkx2gphnJks+dPErtwi0RTXKOHqyi9hhj
3qVaVLgC1xDZrZUT72oYiT+6YhVX2FfN23MjF21t5jw00sEGNFazwY4Nut2JxutgR6MpC3CbdKfz
1c2QWXF45UL7ah6ZqZ4GsDYiA1XPpy5ubrAkqaEcBNS3wRkZ6wG6qzLKItG009fUg+87+4r78Mtu
4V/tlCfM28EANkVuF7soQPi8Ww5YIOKKcvZCfUOUTdd+Xw+k9kaVMnuUr2kHhRZFc8zTNfzjGI8D
S2TiFPRLNbxLP/Pt0/YoCO8H5yMZubO6mPrD9doLS/uDZf7kc+SN6tkzDxVQOPw2kD4FFCKDnAKQ
9jOKU4nHD91/smqIA4S26GS94WEUpJdG0Z4qYWMPmuwHEh1ULKHSvwRMdMm2Az8kP98Apy2oHYl1
dxsovdZXKBDylELVtnM5/QirMgn1sDte7bkQR6hvDsq8dk2oCf0dEBE6zZwG7NbGdLRBMkwWvdpA
ooJbjN0mMbHhWuyNOjnLxfat8s3PbUkTKKFvWVdE1myD+r20RY2crklFAP8hdH1u0THxhEk8Nz0g
0mvDdav4E1je3rmOyRV4VBngQ86WRIJGJog9qYciK+q3vn2wr6bdMf5t5yIZd2Rc7eMIwevL1wVw
9upqoJSTOHbINaXHBEsNdZ4+eJLVL5U0S6/O3oB3GbsAF53LMRUQZ3y+sI5XWgFaXfuBvj5SZhqJ
IjW8MCQRg6isLEEvR+LmKVK+T7BylytNCxlL8fAegLw3S9+o2mZqzPkOzp8oqy99mNFZZUCIK2W0
AugGckgq0XhuKksAkviYIRvdoyn4XYtNQm5/rRcGgz5t9BY7iMvuuxO8ED9qcJjy804ui6MxWPcy
nMGzH5oFE27FicH8CCCV+79egfjvoGNE4AIjIEnyOO50v+S9Qlgx0pjSToIo4q11vFEf3k73WXTY
kucazJ4SeygrpcBuG2LPfgpqiklv7gcw5O3UHa7Jt9o9qyiFdMFIMSGMsZkRl14pHMc8NnpZxppC
NGjSnTvDkYS3BEa1NEMK5l0bAwwsxwpvIMVaiXuikZc3h5BHi2daQ8X4x0zyVGOCgeicuSAEQq0U
knaB0vSXBmgDKCwnq5Or2HBlupLUaXu08WMqg9f5lFZOY1G03MASCU0cvMnpwQwze1KQgC8zlN3l
wra9ziFpIktoQdtD+lQikQN4CqhPkexZ5/qfuZ0TJf4n+pZ4Q5uOd5QltDG5IoOFJGU2epoZFd3q
6lNDPA0qJqPU9aXBAOxANbhySU44JdSqvH4qTi/JTUzKsJk3gwCvR0y/CofAsZ8hF7GyWpZgwdDt
OGO6+iEeGkdyH1njHDhYwu7RMs+2N/PJKxpPgyXNV3CkP4KeHuwWGRq2kwSbzoLm4jyCsJ3sqUqY
rKXYaDq08k54NmTiwFPSHIXxfJk4NmbjW+PxeoeKYF34HUOOd0QPfre33j5rWXTarOY6TFJjvAi9
wqHZXbOotdLYdDS3XrZ77j6/7Rexio/0ldb1uF8bKUOXhDc6MdSHhy5VgnZsjEQYD+k57+kFU4d8
7awgjKlr9uYlnbsS5OYpK+eAY++G9gWes13gCz9SNvyGVgkpDz3FSKaxE9UKPpJoznia4uV9oYfV
ze/8cvEdN9bsQAp26BG4l1yljRD5or3mjoRx5owf8Wp+AVQ2lGORUUH8uo4xqaKrbp44KgPH1PuG
FA0SoJrb1lLQMK9023aVOM9K2k+J3Tpyq9xNciGKNOnnLv4OXnHF9Q0XG+u1pNloEQqFpeIlPYPU
IdP/yGABa/V1Go6/SV72Vjz/GNyfjuBq+7abW53p1zdaCL2enFhy5Op5JslJA24QQQxLy42SWWBy
LSvrul4L3xwI6lL3mYqW9NdSAGMu9dZy+r5gBTP21RLqXlRz4UHofbdpawa/kPDREUjDPqlNsh0c
iZHrWBgqsqzXMr035S/JpMgyOFt/v2eiJPX1D+7/bjuwkoByu3Werp64eOzNGeNMsOZp13S8Cj7D
SPcdgOlC/mQxpQiPuBgH31AZc09xT3UyA1ji8KtFEhV9kZeUkwbYU84hhtDMMCtEE+zoFeirKO6U
cH97QHC52+FZ4yMB6EO8Q15GlZAnbyuunQ0BW6OduPGdvdsv8ap5M1T8FpcSWw29OyiX87Tgfx6O
/f3f8iN8uv+I3U5saelci+45KJJ9J0xvWIxIalob6n8buEAWx2X3OYQba76CS21IGOu0i7ULZUZC
d1n3ZNqujDdOIx9SyofeEbSMuGcLo2F48/ZtkIX4gXuo+HleP4krdU2mICRG/wQ96/vm8D/gDI1C
9GX6gt+bVRBZk/3arX+VSJYSXDOK+BlOYFrAhaW+kWsvvBExUdefBRRztmhspXntrZZRC9VcrDnY
jJaKmaFh+fKeCPTi2Oqb8jkrs/7AV6oxN/LA9ilviS7t2hw01MqIM/OntkZumSboWRuyUqYjJ68r
ch70vGpgkB+woT1aWYpMu43CL6DKnRTo3N4L4S+9/0iQjlgDVYMLmfsLNBVTOJlsc3B+VIgbV6dI
prH3Hi+oroOaGu++m7HiztAS0YhbGvViT4iK4CcXRAOLqrfJMr0CiQ/V1WMf/epWsDcXYLGPq4wP
RV6TwFdj/9nyN9ahcZiKxF1fXldLx++ATcWW7nY/H2f8UeozhXAiMAoC4KwTczrZ57C1PZ5RFT5e
8eNv4VX72mvM6Q9i57zSvQdcAN2dPuHlEMo5LP8S0jTjoMv1hu6mgKIwCUKTWKGYd+G2uFavUFK3
NjJY6MXJ8M/R5/Zfo233nj6/CIrUGulZgM+5RuAKPGSdKmk1c24vz75K1P3E6K2m5mDXP+e3ecd4
aFdHGYm7y0VKMqpuG2YdwaQx6cEwjfhLiUGR/Q6k3DjD00oAPypQd7F9GuhVHU+N5AyY2a+7KfkX
4szd/zb+X3sVa003Ei6eUhKprnpI8gAmG2Y4TzV+qdFsz6o6qqK9yuqXAkv5bZ994nU1/GnQDEFP
sCpmHzogOhyQznbTTnFv9XTKCZoUcVlmznfiAlKkD3yFBDEfr8ARz/5lopTD/++rodBIFUWWnWGB
usTUSkapIKV+YczYAzSGV7LRDPMQFWbxQJ/C2uBKxyymASszt9SGYrewmt5fH8/5YeFrZRkqnMjY
o7pgxpnhjUZWex2PFk4BReGpRs6Jr2pQkOhQsbxVB9eYgIbeN62KFVB2SHGxea7KehoY2m95yvIc
R1CKJ1mzlVWPaBj+isj+iCx95OVH0taoD9sBN0Bv+ammubhwpYKcMHpGMQTekWixHoW3d8OSLt9w
zVrTj0PbRh/djGfX6FZI8uFBTiur9y4biB6Uzwjm5qNm9CBQqIUxozLwCP1Yf9y2LomGo79Cm7Xs
wjmUWVweeeEu4A4P4zmf6ZIH5gCfDAWMWwR0wxO75kTzk8mTVnwZrDlsfQ4AId1b7jF9nM7ypaPg
GXYCAgrZxN+ovNvbXvbnbSQE4FijPota2Apdd4A3zNgil7qp+1+fStUGxKWg741pgX6jwxGbg3nc
PfUakd7hLJ71vts17Qo8VIsmfHHiQESV6SNrbZYoKgz4xpx1oPP9UfPleXdxpwMcQAAH8h0uBq/N
d/WR7RdCrnhd83y3XMJO+Ewh78KMtspr88DruMHGKq2Crvx5mGpEMZ9P1KeuZ7IrUrsWId7jtoYQ
CRRNAvT5gxIEVc5/lEXac5xw7Dk9Ze2tbQWbbuvNyG54SeIl+z5xpAcbsisMjfeSdcOtvyG4oqsp
oIGxzr0Cn+t5+Xqm1dhiwW60AoPay+AhMVfht3ZNhk3hw6yVDW9+GjBlWNBwF522rYr4cOrUCats
K5629q7n+O24yYp6IalWBMwIDsjjoGJOf/bzaUabkL8tt6LcxssO65J1q9RoyQFTG044h03yQke/
cEppkewWRDAIrn7yCEkrW33mDnwVcWNCdPU4W3kRT/YlFCKWnklrAg8jAxYFWTykdMKcIfEO/2QV
4QA2tZMA/fczFjZ/1t+rBAlidz+J/LS7Vy/k/QZuWSuDa4syB5YEwM1LKmFh67zTP1xML160RV+A
BxXWF+9NU4CM960UfWSxKNsLPSw9+7ZNBt5m3xt6pNCDIN0ZR/C0F54MGMycuRvJGd/a/JHHJFjB
R5zX0uwH83+S1XLw3ufxT72tvGVkMh7BpU2Ke/AiIclv4+tAdvcSVxti1sRSnAYrkt0AD5HKXEr6
wJeqen4aEdf6LuR11OVbZwhsk/BrHZXdszI+K7P5wa+RK0XAubgeTXwq8i5eE1T3doMk060fDTBD
PKi6c4KrH+pXYQoEOvJLcRt7ifNQoSZQWkWOUzijwFf1vS7KF8AkYldfs4IG/yfXONHJN8wh2XKm
du2d/bRqK2neP01AoGajmonCnD6JXcP708CMfa4aGIZoWi8K3lF24uHUgzAdLFNGosmuJHKWe6n+
cVGnjPgxvO27L47okkB6zGiaShtTst+tNExwgd09idyOWJPlLoGjTaQvsTTKJO7G9vC94FOVR4Fo
gvYrQiD/lWkwmTAGMjPOWvclI+aTPlX+QGY7YJvzMBa2dPiQtvLfKr8aaK8GDBRowGvC4AzXGR5j
kxMoHx/V1H0m20oaopRUTDccfQ+O7dNJBelQfiTRxiOCUntc54J3Z9d+RqFXc61reHFfsFcIW3Yi
30Brssso6VGFl8rv7y22/eXQyWqvx/XQGm6YTHb52ZvA42y11atf6pGsoy/MmlCh3FwaYa9g/j0F
giKREwI/ufKvqkdxtTmso8r9nEW0tZqAFN6lFOCZ9veYR1gwiBCOOJBVxHiuKI5bSKw37Kz7BLWX
mv1YheBWE1sgjmAUyPPwzo5IQT2DBgMytzAYUU1DdlT7y4tAsTuOmbsYl8In/UoaXSng40C9QRBw
BCgHHk5skGYaR5oR5puZs8uli+Xw2LzHyYJt2oHWrCQptIDWC5Wo/M1oRTed6GLXi7RSH9mTVc0Q
m2yy3HR+FWZJm4nvFxM8gAUhUt6p3+P0bRjMnEgD3PKL2IFv0afhLDOdW0NTqwFHTdz93UNaIKlU
zaO2sk4xt8WKU1YxgJtc9UosfGYP9ijmU4UizK64SmMMOhTfdcpogoGazBCnFtkKe8vn2ZO/xVo6
0ppmQWngurOrOnYhJLzQfOldABeh5I13ehlSxt0oryR0E6i1bq+PKAlkSYb+OMCO1os0caQza6ey
bqCeLDiYh/LYAUOWn73Yky1VLBWeGhMPmt8kQo1aK66srLdo/JwcHCGKukS41e25rBfKoNdJXQPI
oN5oHK0iQOu/5GYosvRGxyXKCCQiCvv5wv4qSYRWwR4jhXf5imoPAPXYfIEhrwJWwK33kyIRGyJF
WmP+dl72uXxfrEX8P5cj6YLINU5PkkGa28eGb284a8+YyxUV97AOj3COX0C8fpBjKlP+VCuuhBAk
Bi1PaLNO7GslZWlpE3vPjUnACLSv9Zm6oEcFUabcB1QuSoIgyItDNYAT6abMfC0QYw2ObFEeFkYi
BK/NVG8ujwHOQfkgF4YsNEAIpm2Ud4pE450XnMv1XWtsnu0VmQWrOKllsytTczxOikWXF7qLi3c2
xpKHXxs1sZKEnBkFgw/gAYU8YtqqgpiTuuHXWTh0axGwVgXpVs4Tf6GhQc6k6d8UQoFdWWze2VOL
9cDDHsQI25IjZPjK2NLQvTgKSbAi1/vL1+hLW0ahfp/ei5zOFrcZpW6UhgqSIXFHTsE3RvSLPO+7
hYTc0LOLc0tnM+oHwxCWdd9Ay+4gYrrPpSQUcjhN/ifJcPd61mP45SrFfUO+WE+HDjkM4/VA4amQ
UpxQ2EBP9STz1kjylpd3DftJSMmtmeaMmsxfFNbSGnag/GeiKwgxq9OkK2ThOn5i6aK3KNCxMqac
qBeVBl7ZLmUQjCAFqI3+lBSF12IZr4lk6yge6VagGVhn7TuQp5+uFVt+zlGrdubIk5WH55x9dmsH
dhrkqH3YFi5I3P3oKEV0DYnoWgGHzU1+rR/tvwkPOc6XRBGRlawXrKl7JRBIVxMz0mdIOjCYSPHs
y63U1oc/JaqrULD0s171ACg4mOupUIowsZBrx0aybD128rb8VDHtPTDEJy/1dGDvb0Lerp71jCIg
doMew5ScaqS2BDUCV9EOXkBo+GskgvhpKnOoQT4BT7Ld3GrEpyLRiOpeqZoNGJxQ+SQPdjS1HlAL
5X63FHjI792Szz4fuVqQJasdIZLDdNKrYlHrGV1EOyD5uuBdpt2dImcsznvcMcA+LxikiwtF2Dc8
0xR/4Vx/5OvClNN5uGyI+TDunuLI9Cme5KxMmQej7h9hqhpAEJyyfZNPkR9yDB1RmOllO3VJKlfr
cWc1Q247ACeUz/FdZrgtFSpE+zfpIUpnkbbYM2kq6n/OCAdgWVGnkwWXeokfnCV430dmvB1TL/B5
3zXBuVQ6/SiXwXMLalYgJoOHXac4oHIO4u2vz+ui9V4YvTwgxdIj/UDhKjO129If8lorWDSVgfNk
hFWzJR0v1fvULBWm/HxY+P7Wu9R4hQxjBzqYl5MNBXndI4yHxccfaXPeK6YIFVzZG+O3oz6sshwL
J5zG0Z0PyfcwG8x9KTtzy8CRdrBhx192kJZhi+Qf6Fk2xjb0pMhEYl2EKkP+nk5v5FxG5/Sror9w
nJNgB5xGC0cfbfwTARACwlfTqeQb2f6Mi8G487U550c7mLCz32mm3T8qKXayTZPbGdzUvl5uMtW1
zl98S5MVUwDru0Du6HNItXdVT5KRSn2pKiingaFa+M2CgQkCLOR6WirMPq7PeQa8/HCsAZDznEGs
FN9wAwBUm8TPflD+DKrsLZtorT825hDId7dkzoCi8qoKT96EuaI6Gdwv34SGNV33ooE4p28JZ5xJ
IDk2yWU7ygpMcvzC1g92lMLVaZkHDunGVFBpA7MytPKQjuN4XN9Cd6jbBjbHLr++VGsGoQTlqnWC
dBvos7YkJVC7K4iT8ZJ8q4SHX9El3MiVx0F6EzpWS06IeDsGZm4aZqqlxOuN5gMAwxEH6u1fvxua
SKrqqQm0QJ98yurJVC7bDayLdcFpoTsKkxZekXmUi5QkLuoZhqCB2qugnxVL6xwON3njo+t+W0rI
3g+yiqUdoQ6PDC/bg3nVxVcQMAPLP1kfSqvx0d1DwOCXQeFfW9woMkeDPuFZjzmS3xCpglOTo76F
6+N0+1v997Wq+Dqs4t7+ByQhKuDUxx8SuogPjtD+pMh+gYC2st38/qPzewJSeRFavjIOmwxr4fUE
+aphv0jpZ1TUZIpKjcvdUo5hoewTGyMRiuNOH1yJVbkBtRD/9JI+vEOmswrE+IhmRy2B3N0m3c5T
dyQH6q9+/hg0U+EfP2UsA8bbRKQyo0FFPJl7DPNpfUP2Q2HhHjD1IeF0I2duHgiyG4Myr8cF3NG7
SsPm+ahHmdypypW+S+pMWOZE33FcORwEI36H5efCpxg4Fzo/s2AdzKppxT6LkhH+fMIY9BVvEOZH
/kkEnfXJKLpsYD0o16NTDyRS+PsHbzuAm8XAFbUGj4kpQFY4+FNb32/HQMZbOrkJCn5fAMrLEnPk
tr203U3KkyJtIEI/BrgwB+1ueBXOlod07G6WPqp5tAqS0fQzpjtQc3+r40WraZNTeGxoxDA/7PhG
2KKei+GDDOACyBCK+PGbMu9o5YUBbQJt0WdhrWS6DGX2I7jJEjr/oJCy4FCCwSaR6CSkV2ySqdzk
h4YSGkbS7KA7/0J+uCyzWV/uwEdVmaXd2fmAL579yKGFjn16Nge0G6n8Wh72ZQoG7dPygP75LQjb
dVXpPX/cY7pRNHg9aABYlLdJTB5TlG3x1sq5dLm69iL2ENhwThdR1dVJvvQ4x9/WDEb/3iXtp6Kg
h+EPhK0BLrPG0nknQZl8SGJPt+Dw8LFH/Umjuv4GfyXQNuSoQEOqZqNyT9rUn9klarkbC8/wUmZj
GV89fISagozv1MiqZj4EiuRBnMd/O/SLceYb9hEcyxwqnSiNEix8eblqVmdrQU8zG7VLMzzSjcKl
DLp07+MmUS/rggDWwnw0cT32tQBO8T+QaHahZGmF6bpPwC6AZBF7hLdfn3KRCb/xm3iCOt84fQZz
jVskx2mYMVXYLQ7ayM9ruWjbzQS7uuj6SRZKM+tXliVNCvLuyzLnF5vaNJDw77lh7gZddOMfWKGg
BmX79XC4euMJPCCDx5fPZIpQb0+gFJ3KKKgl6+uNeqyyGFcAVkG+UO2/SV3aeJyqCd3heQJhZk4s
CpTvthCcJs0/29M9SxZejQAfYNrRZNLGCNVdQfP5Z+Wvg/IQlsX5ApCi0oUpARdIg00go1gvM3vl
gSDLdtYYojTk8s7hezZ2L8H8hS/RUfcfoPAzYF4IxDjQyJrmBXLWw4ZKMmIodquBX8rbcLZTVUAy
9hC5W7EBd85YAHEDHLtKxZaOpZi1quvSK0oFdvKmL+TQthD1H7K94WxjaB6unZk4SM2HPqhscC8A
RYdmFHKTg0v4k6j6NzxcQLVyROtXYn3y1/x9kASYSyCBSph5tPniIqKoDwUzNZg9Lml4wAAQHD5T
dnUzAdwN0mTzUog6jnp2yd7lUTEeE0a1SsHo6EP+cUWxYEFljhPGniYKYul4kH0y4ml9MlkCFwr9
naMZ/ttBTGfHlIjD7Xyt/gPnvZwWWrYD8Df4H1vYOhhgDzH8cWo8muyfMX0CPRTcEkWoQoOhRge/
ZguREv6y1ER7Y+0+J6Wnnv5lTfHK3FGSmCEENE9NzbX2xlRrbgE4fCEFVg3iiOSW9Pit6VIjlCKu
KVbisUreY7/7dvJO8F8eECgtboDZW57AkskgG3ApMgnHgUSrQXCC53MWeEmk12lo6oESfsuYydvO
liR9fPQcmnKXDsaaNbybix28Rg30EI4i7Jk82hnwXq+coVHadp3xynY/ws/HgF65OaFJ/dDy406r
iGiDwXN0q0eWSlgeNnl4Q4VL50g9SIP3ZqYP0gXk8RevRJf960U22JbZm//TzLE66c/woRPmEq2a
JvhCyGvMLqedCXSrYpiMiq8ZZ3Kh5vPSUCrjLp0moXhVnGQq88ULAgMlzzfZ/opVOMe1/IJNSl1m
EbC6mfECJEMDFp1HMg7O02aIyjRi+rZHctpB0Nni+C5pjCBlEVmqo+rKdlulvspU+AwxWhwnLH++
6NBdHr8W6cOYbFp9WwLb3/iLE1lc33rFLAXQqCbrrvryclVSLOmCIvc6SCayUJxIcn0Rut8m4q6A
WAhmT+h3ye6MxGsle6ZlY/dXpoDQJ6G3FgBDqsh+AU1j7y9771Pm2M+XRjYROb32g53giN21kAfe
lMwaXcxCCR7P5bdLnUrobUZQKFDqi7bGmKahQu239qU5K/WIDDM92ivfu9BEqNUEWnC0/33n8Tq+
iyIl8rH5rWxs+6iJojlNcA68CkhItMLtIlO47dNR+apGJTZu9dJQgch8jhInXbcl5V9mXRrZK2WP
Qk87Dwo355Xr9f6+nzJHESl5HASIEO0VVaw6ovDIbnxXJm923zNnJCo4jCZ35F4hGZ50NgsGuJ6X
RUEuTE6pn3Rw5cz/Tk2Nd0O2vzSD0u545wDPJMAdkOijlOmL/kWjkZHn30MwJJdsX8diBMQfi4Tr
W+Iu4LC6fYIcDXQY65MN8SD96kZPGf9BQUaK6C7zlolRRat7+Gwb9Z09uB3JziUffJ1JVlCJFxZa
Wmus8wPvo/YTxeL/VMj8xt82dPQvNIp0QWlb+P8wiVCPvystC722R7nBI6PmVco5jP5Xz2xSg9Qb
gWnmP2OWAzb5yk3fFIhE4chooilSRSlwY/wliAWat9TI6WlJi2I0fQ5hFsstIGCsetd4Xjr8aAXg
30ghYiQFUGNyoEgQdem4BvgrGw45n/FfFkK2JDB+8jCo2ltaAdgm2Qa1m3mvITWV/p2+Crahii7j
JEqcxRirbFKAn3p+ZI2tOm+sZXZ1U+jlJcbBxhZ9D9ymDpGRueznKWP/P25iDn1E/Ef7v9MJQcdV
k6Cr4ZFx1eRMBPbUVHgmhjtchAY/DxGuOFdumwvO+MEluK+AMXK9y2TFOikWFi9X8LLzln6zuveH
IZNVn337ZUXcyywVsHBsPwKEVihbGzAo6pJt1+jRLiqHeKgdyLRf+Z2JVF3MuKupiPth8Tpv2KqI
cir2B7TaYuzd8yHUCnrK5CsByP5eLaU/akNL9ZNuUKI/yaLjY6zqUo/poIV0EdpEpFA0wc3xZ0r8
5DCmxBrw1q5ugaSAZVvye/W/UtNyVNntIPNX0RPANQcsC9Cw3fpcKGc1wosUI1HJYXyqByFuests
qXelt0y8ToAJZ0tug78K/i83DP8XV/GOzC0WDEyVjhYU3x9aaSeQ7tDN+St21g/kaDp0DpQAiwJ/
pDpFQ4er6rFezC72WZGpjaW1Ev/EdqzTKzmJo8wITeTtIDt5um67fT742t8nF841rDEv7zPwPOdA
dj5yh/TPVUKxaFfV12qPzjduA8YIGhcKiFNhFXlbZv6FZfw+mzxcFr8J4zJTykbhgcHuGw2nzGB4
aKWuCpM6diZx8TKI+aHWwAZ5GOfeeIXciwKPBA84GUVWsEba1Y4Gc8nzznFkiHlkcbmHN4CC3IDD
/AyRmQ1Rcj8O8LegiqSV3rAvEcCBXIi0eWgxffTNQXqs1HvxKZIAwdxozRMVYZKyNhJjiQgqmkwz
OZqKiPZM57yQMHhlstFKTbrWX+WAn42qBsXV8+tg29oFgvGTWl8lL54R+hhECBorGvIkQNU6UCp7
52+VMogLnQpp0z+TTnBrUJI53qCb+qdjds8EzuuNiEl3YVHIG/PGDCSLpucZe4MH2/qh20Qs14Ey
XZiot+tl9xix8G1rcYB2lpjid2oSlFOXzKaViRRscK2+tXsdy8MCwFkhwOx0pE7g3nhAGhT2xyJH
1gvKj3e2lhRFqpWjmUnYgMJttzSe3owMIw6aBg++4YsK9vxTQOl6DrKnkrHJk5jaG2TbjT2CGL4u
HPxLaxGK31rEuog1xRIgqP1veG4Rb94QBzZnEcBdxonCAHRNcEzjOHyH2wmCVaTVQ2FgyIVGFrE4
cs4UeGWqF9aFlRTrMbUoadLggGLJHw3r+g71e0E4pSJkR3J19xuSSnkmueLJaqeUQI9kLXpOUZ0U
9xSd2Y1j1SDMw5lH8Q7eJML0NBeCpUJeV8Ht7B3VOIOW0yVC5gBKFggwCchO+/bA0EMDE3u7rcVt
mNuoWGbZYQYBezbiW07bRZNAHhfCcfWD1Lf7qKmufEnPiUIdwgngkEC9Uj4f044MmWxw8sMrqXie
Pc4aIsl8fVj8JFbH7Tx5Na7V556g1u7hRwR8VW2qlPQXSlSEwg7vGbKVcuCENic9ZhCCRC4CjAUW
rT0wVq1YZfJagP+CLFT7Y54h9BNxVIGk7+B1RLNZHSKNbNJPkPW7bm7rnkeg78yOd/E0Rvvzc2Qu
XUa+fgPuaot05ogrLKXhUEGd+o2WspR1FltD2xhkNkg5fGssymX6mbv3h+2jVDlrapYGBTXsemr1
WgM3Py19p9q+GqaYQph78qWyOYXPY2z2dJspbR1k3JCBbVQQVdpXFnUNir0XzXCL4AbUgAwLGwok
KX6d5K3SMrDVwzAQtO5tUvYIHiILDBjpRq26UMzsC/RY804ddX8UZiQzP6kPfOWDExCtRa2W8DeZ
KLi8f2DrqbCodSMVz9ldzpfX4wrXwUKSMWGvaI+2+W4WeGOb+iZAtncdyWCu4iw5vMUcthe+42vw
C2Vp8euX0yYLqN4DGEW0uE9pD6bivsaKpv+cKmSjit9yl9deYqgdVzdIVjuX1mUm0VnM2G1quZ4t
kR2/gDISowxuIJtdGWIZXmykyEXBg+2fUWGjwWG2ZkUAR5os34ugnJ5YTPEprOEh08CzITWGNAxr
+Etws5/4/pOwzDcJy+KdLhlmuSaZF3iFGuVvd+qViaayjSjnCgB348HQPlYdoiM8NnTCazM6wfaY
LNxrsuCv5OXxHs5Jl0BMXK+U16aT3fLwzb17MmMrAYD2ZpfytjW4eVPrIg/A3DkeQP927GQa3xmZ
+GbOoXD0mx7V/Cc7Y5e8cGoPvx1Rb6sP+cSQpub4EDmnT+nRVqAcG13D3odPw1wNBBS7jqugAysg
doTIi0N9/4u48zclx/jvAiaBk8NtouUZfzmAuwQS0yWePRDGs4TfeEQa2jSR1hEiP7hJq2c7ZnR3
8pN+RjU4wIWrIJGkQpfY9xb9hBkicAEUccE4zGATkjT3Q+0IV6WVsbJJeHUPYlcOZJOCVR2LCxrC
GZBoxJVeZRUsbxAH2rNAcPEVj+/wuboMJVZ6KLjwBWy+maNmgPVGRN1B4vLWbkq/ewSnTi9pl3Sf
Hfu0Eqinjwum7n/Kd8Z8IiuTPQ6o9EPc0mSuiaYZ6hp+9fqHcXlnvFhPWaVlTOCUnwBJ1AksXlE0
yw9fGQPeDhiGwJFsxNQwQdFp1NIJdLkDkMtjiMTJtBQb6tO/OMNN7wq8W3wAvVhc3R/1iW6tyanV
PRsoYrUMW7M/e5838NqBGFranyhmdLuIvIO/kcDa6CXGMvKdYzN9VpfVc9lmIdU2AYX48HZcM5t6
nnOjY3jmuZTjMirNVp9HvUlkSt9z2d6RKdjLMCXAgQVCExR6dzbr3yetYQrmd2vBQI8WNxiyfWi6
6yqqVfic9f72I0gZ1ciSGpiT1p9TrwxcLcGaJwY5NfhnCw8vCNUrhZ/jmsH5DVWZH+6Ej5uRRn6Z
Ae1RxIvpqArb5w9jwh349Mto1tNReBGexpUhMb8st6iHy20seAzt8txZ64IvaNOGOk1qY/cqS74+
h9CXT9UX9zJhL2bMkHB4ToV1ahsTd+30otBhvE7efhJwj52BnonwVVPZmLLTe2+yVIMfCVeRz0uD
iRVU4eQzPkFUDrDjgcSnAzCaoNJyjSU3M3VZU9krVcTmu/NcecxuCSFSvbGtbSHgqM7213vPDKZi
AWymXyaJwmZDc97KJ/ZDIo6Q17UeV1D7HyPR7H6ecpvBob7B2s2PoD6UIcKuuWqn656laqORHRPG
n1eIdl7CI0ZXwKeByDOBc7NtUrOO68gzH7ZcGDwiyWrGxvWO1MKRtjv4MVh5HYrFMYjstr8LhBxV
nM9zeefx39GkwP/Bjt94zxf1K1z+SQ3ShIiPupkjXg2/QFM0jf15TcqElHh4RKSjCs0SIAZ0qePw
xXxw6N14tBkO640Q27mX9J9P8ZSSVLMSPAMg49HqPn7uvGnSY8RBu7clTnF4PyFSRLnHYXp8MJTX
Fe48vobezDOY49ojad0CUo+TMSixR0mB5rXGtvsM0LC1yGExCLWzbwRlhQEnCnXyrLPxCjcfsyNW
N88yGvFRd/7I2RJZn/+AdOVGd+SiVYQ8hkQRqknlWCCL9OmzyjOGsnlBj7eNQp2CYXErIv2Z2wLP
8MCkUycQaJSdztt8osSao6UECLdnTsY5I/zLFdljAgMs7lx0QcsVIzYwp9E75o6TrQCQN6CRcgZv
XkNUUxhqZYte7ZmS0EjP4E4Qhn4+UOBBkH8OZ94fdeBuu4LsIBgPusFBY+GKS/k3NCyFRMaHmZt+
DJU2az/RtjqAV/0P+Kue+pSC1MJ/mYAcS0jx4aUc9QFMagkePsnUjA9fZfrebclwN4qC+m9LIP3u
0WA7u6aMWmc74JsXMlY8iC2CtczS9EO8GZmeIj1+7K8oi8OC4TVY0J8dM8IyyraINxTWfuEP0B43
QFnxj7zSxaISv2QKM7NgeCUZFkHGwxgPUP4NbRS/YvxgM25971J7hFEpn/lDPVMYaRnU86lAeaW/
qYnSrEFRKlPA/HBNvOF/yssyOAFrnxkMG0AMinRSae96attNrNZckNXUpg+yy9iW8/+KB+W61u3z
or0V78F2aSGWrgPC3NxuOUC7UNPu9uID6IvARsyidXlKOYuZVB0LaTqxqpJ5ZKZNd5XzGq3/t1q8
x63I5X8RWFCmtrsuhe84RrPi1Uk4G8FVRQIzc1zFcJiTfqlU/FkSvM18lsJ29E9uQ5CWztasxkNn
nxYlP8sj15hA/uMZLUEzrUWjlaPac6ItN6Vso47d9kA8R9NI4mB8o+lYizR++EsRbFdGtdTiSfSo
WGDFgyMM5JSZsJgZDrQ/h2lmepx44pPzYQ9AdvH7XfNBd303nMIyH4tXzIJ/VGANE/ajCrBzyotV
sjx/ZYd0qrY7DtZ2ChpinbRmMraOK4KsagoGnOnqP1J3NI8C+hSexr6G71+wFFjs6G5vn0Ni2rcz
jUq12ZdFnPgYaAak8TlbvLr+QkOeueHvml455j8RVs2byIWp7e6ptjMYGhSM8SPZ5D6yp+y4Vm9r
bhV4oKUqFQOjkoaTDbHLw78y6WrJrACd1uxi819ZAyVpeq614sGcv3rCAFCDlkI8snnhT4Dz/gia
GCqHRzvdhuUiQdB+3CnoGOMBqXRAQWyGEnMuEJXYmIFs8Ml19HLURxHZWPPtqn1EmhY++xiwebjE
dCcs/Eapw68kT8pnCOT32DLR50alOMb+vvH8DaXv/X0z0pbLbfP1b8XCawe3iHZ19l2K0UBz8vKV
+/VuPWwPOyG+udRc+FZAOywFAnXG4yJjBPieiYEcs0bCnI6sTTQ1JKZs9OqXKSyE4wrCI10OsRct
bJWDVFNH3ua8XNv2QZ183rw4NfiyA7zr+Cq+308jfNcOUTSd1mtVpCzJXD7YjeSbYTFvpJUnZfKj
jNU5lJNnktaRiVlGRKnnmQS/Lmq1YFE3b/GJJo/NM4cKkgBhDubTAR6PgcNZUspcnv1FxYI92B8h
UT/ljSfDcfgWX4TqJWneKRFokjYmGVvwoNVZ8ZpA2vwHFFR6L0S49UmbNj07v0kH/D4bBxU5grXQ
JX3z+VCA7XC74KwpAhroqeO91VvczHh2GnD2pmxIuUku2V54eaP8DJVbnMEk6EQ6Zk+N7G8Ypaca
oOOarxAIUIZP0vIK1GtPmODeU3UQ2ThWxr/tUUTylo88qY/520i6s9Eonbthno2MQ+Hi1+WphWkf
GZ+EXvpkBiQfxgUSsJ3cHSkta7R3jlZ+3eXybaDdw8dtE6IQHAAhjC7H/x0MyPPzNtNZeDKUzX3f
0Td6k5vsBl1I2c8iIgenfDZecXtsAeytaDKK8Yh9c9JOv+KOzJ8B6MisfNNrs71NFrHvxWpa9HZp
P1ICNRCLlQZtwAKQeJLxnXH9KT1S5bIxd2C6q1OY21mudIHOPHrf5ow9XhdqIBlw9BZ89Wb/Z2Ap
0vkxWCXxCcqZbTlZdqBz3eO8xLMbKkx95od57hRQalLJLT7oRXID8L12KzdvlmxXxixzmSXL7ZKD
/kC42LQXEkeT5tG8mJEAnl8p64Kn5RtH57IEQO78QdnyqXTi3aKCYyVRVlxlBTI5Zkdq1GStVQSA
a7+pEuFyC5PonXT/KNKCjYUc2Dcyok/Cm5hPEh8ux+utvGH4ZMo29E5EG1jUuGzYr9aNv0IJDDdD
hqydlyilzR+Zkm5h0vnNZOIIfndP6Un/uECwVqyItTs3IiFHwfiDw/dWLKmOLxXLo1QxDfjiUgFa
tOSoR6Dmf9Gid7uycF4sNuI0G1ksmCJMXAntYHr8oJF59RLArCPpio4pSZ4ekLn+qbk+7AwJpvsX
b82/WuSa1S3CJgl/ENEmVuSOP36WS5hZ9le/nQHVsplS9uORxMFBcNI81CWaR22yxZMQEm21Qt55
LfhjCoSU5h2vJ2p0rkQYGPjoovQZFWMlspB7IUCrOlDS3AxOphqWD4efxLekY8YV8BHkDNeKmeNa
eUEUmMwzgD8OVUY8tGC6rO//JpZj/rDGqa1RO9hrtm3f9RxwlXNpc8FP4wCXYWfIDfdL26TofYt3
R+sDVPYqUH3VLKGUJy+RKTL7yJ7F31dpsiwmAPlbx0yo1HXGIvg6ljvSTr/9qtoxshtMB57TZIDB
G9Z/AhdpxecjLm2bjFCmxqxUHQ3dyV8DnSjkvGXNqKQBi4XYZsvvHe9MkMuCVFmVeCVaGNRFhCAt
evtag7+d9lFRcYv7kWPqk93uhRn6KJQKnis42apNdezgh5vGP+/ht3/pwpxhFct/bmU0Wzh1KqrZ
ACQVKbL9LDqOElUxGhjuGUz/m69/TXBM+UiRCAcUPxDOU6wweHG6LQSAN6DGkSXkYT1fiC43vt8/
aJn7syLiXcgh/PZvRKvXW7KV0tuIJvu0MWX97fmJv4tGQWyiFHb1ZTCrZCbjNzaKioZwoaaxOv74
Lgc14nGVIEbR6hxFf3QyrsUP0C9TSTF3tyu+8w6sNvcFoMYfMge89Vq4pfkwmAQITJQVZDx2ZPjV
lkYYWOZs+sRsvIjLQtz96deI+HkSWtCFds0YZJzOpviDeNRm1tqelTsHzwD9KDHnx7Q53xdfgzxx
FSwaeybyJUpFTWxtFExz+OPh9nOyVgQJhu8Oet37truUvUzXOijmFGLubmbfjrA0h/qv7oooE9V/
Yot2pBsyURRKkYkttycCxuGcCvlHrlKUAIPWUZOVpa1yzrENmEjxytkxdbf5Hi5LosHyPjbToaBQ
kosV/16I/usOf6OYqzsKmhSvAr+qL88uO05uJWdor+wROn/xwFa/7Z4tn743usNh9BLO9SXGpsD0
B5sGUBtzMlYFHeZ4IQkM4OwsOD7s2hkZC0lrrMKHH2hf5X7/jOOaqQYpjKnvKwFrTNf6dDiHiaak
Qkb64yJCQXym5pUBPIVYh/0ZowwxxOU4R2MDOprXA1ZorZbufbCNv6eM4YxGCT1AVm2rOwguCMpH
2SxQ3fexRt5wu7igXdQO5SkmrSXU26Tq19liW00S2zFUkIzrQFRCH0jvOoYXTOYn/jgwKB3KRkpe
LYoVSLsJvlELp212U+tJX0HXS/iGZoIUBskaIUYm5Bn5kPc0oUbUbKAI2d+4/aeXL6o0q8zcY/p7
OPcrAAUi8UT/NGu9xKMj/pne5bcqkGlqkPZSIBDu0pmbBXFyIRrVfEcLbC5hL93ik1ARMXPZJcaA
Oena5nve0dir2wC5HDwQw3zs/xzl0SoXlzVK5BV28aHSMqxf0lvPBtzf0x3Aq66VdAQBRSn6TxyJ
qdagy33LEZRpjm3LOaxdBgBD2Dp0voq1NLgZa6LfbsQHlksG6GEdMegGji0/xLQgfeqI04w7fPpd
8TVsUGctus9IJ/KemAICvnr3GrttgSs9sEAg1MQfC6CfhyfQtEtnXJM9Yx/6iJChGHwdzk0s5GsD
TIJHmA0iFvBIhHSn3OI/4SVwBRICKzeoVUGKWc8WmdUp7WpbnU6fH+szhnCoZrXMjkasbi565r4e
Xc1nlTSDV+QhbzbUi6UIfrY5v9EvaHDVoHuolTts1PmWyBAmcDvfAD+bucFNXAw03P5g93e/HXN8
CU+UH99jh5au4jXu9mlh0b4I8z6pm+QcTJxzuU4yO4rWPRricoJW8p80uE2EP43ik0SxLpxXFq1p
iBKb6mVqn4aQTe8dtWbkV7fVkaZf/ubCmpfbfn2BIxpL2+5sfXvJ8ZQD6477U/U8DOdHA3HbH35K
GlGvMPzPf+CKCb2tVcl/QX8vOQx3yXIvfuJaClqXNB7ctgUT1wtHCRAncNyeQQdWamv465/o8sec
Qt/sZQBHmjXXP51CPTp/mEtOT9fJq0ngP13Gv+qKS9fcPVbCaquzPxX0lFG29Y4wcKippvnvKeIV
dYgZgF4/nZJXPo3N6xacNZSWHq7Ibpqy0X+UbqT7Sz5cn/2+Vnpp4EoT0I1sb5acgGOR+0l5+ek6
5PbfcU0nTlB1KEDmw1W+wF08vveFtoA8okkk8KHH6khtFH+tgCdYmQQkUyytCUd34QqOcrVnfm3l
K/ICxmtEXXVJfoY7pGvzcGqdnh3f4dL9NZPNjoWJPGGokRQDDQtsUUTuw7f8vRiHNnkIamICNxzy
Brz8EK6MYSrwdf0ijn8XiG/yiY3A7NXPZiLVhe5naRrWAXuYylVyYXWrrvEAXAWvwePxKfiv/dYW
tsjogDWVUlG4fV6qVSFrolz6Ow7HwiGM7QXbZybbsI5J70NxIwVxZCunC66BxtO6GsKOyETweNIm
bfBmMaXEP1Hf1yKnBDcXXygs2T0y91i1e0eS/V0WglC7ZC5kPscYrqmPOsfvPb9URPupBcuUBAqO
b67QBhRVWF528KLflGFDNVeVhxI/vpw6gVhn34whaVPRzv0fVPAWRP/I9rjHgWoqeX1E1CThzvhJ
p75O4FP6oq2KGM4cN9Cg6n34+fwelu0S8JNatayoegzz1crX2/sVjpTIHh717OA8vEZn9zyy+aD4
54VsNWfyLBbMqzqB4oZBR54G/4fUEs30yqUNVh75Upj6NIi41IbjqbDHd6Ar1OQQ61oTveFVhsJb
XclPMRiXIDdHxPsayp8lxEKh7/vwY/6oPMwBw+dgwI+8oJvDcUfc0UBaZPpjNz3yqf+8SbpgyzHH
XWx+J7j0a1sKsXGNE97jIcesVyXMLpHOqJAYitZaO3U9PNP58h3xR1pkH0VV/5d0SfN86cr0XlHA
dPpAMpDIp1FphU81tplp7hrPaG2yiZFzVwgPh9SBsuBNPFpPp8UuK0CNWyVKBJbGgoqtKxJdQhCl
Ah205V0rWjh6fe8945mB9ok6XH4JuhmU6N6O8F+1jM6qmHC0VS2i4tVR1Ykd7w4C0NIC9pfVD1By
WKoRPt5MDR/Hz44fA6YJ1D4oNU+3AzGGdKObt+77IjT4F1bP2nljTJrvaoquUPUKFz8N8JsORcwn
8DuStkf/5s+/ro4uOCI9VHPkdfdMzQHfQw+WsxgvXFNspW4MNvjiUAAw4WWdwnO+bXdHVnuuhzAr
5sENhrSXaH2n28bzRTqH2thvmsMXLZRh95Olr1o88vK2iMzXNTZtW2a7ZVaM4r4XzyrZR3GPY0EY
2rJfbq/76Ji0VSUN4WU90KzlaSuLjsJs03SskmD0hXZmK+lflpiGOmmBASAetHI7E4J7ngBUgaqA
G0d5gu7uAVOUABLe0P9ZIPZiwZ2/uCGxa5hJz83j6RjQ/NYJyRHcKD7xc2hUtkB4pqJFZDupFDyE
DOFCseQqI6oAEyiS6DiDdEmsTcYLolsMrdts8EVNpKXWrlF3nf7Qji+vnTUolo77BIXPQoWV8GmL
R7yFIg48z5Dq+l8eSD11fsjUXtuFKsHY4JA//i0E2N3t7iO5wymZ9ojf/LLVirQAdR8qSVejO9Ci
QJRqSaJq0OcfSf/TQAKx4b+fleyWuZ9z5KRHYRwbSxOuoDbPMqlI6/gkxVyTkdEghuoQhhmNqzbU
7tvr68qerO8yWAf87DMgeC+6v/pF132TTbYNIUyjB8a/pErzOu663Sxiu7kPxofgBnL7wvFbJyZp
EC5kUmGNvvCbmcz81OLHufF/Cm4lGq2QRc/g27EDucdNwV2ycLcp6GOVgR3s09m3UDrPuG4oD491
JAVdJMCuBlnBxHEMJrSdU2EH1KGDXL3Qq3hMAIghLXe+3VTvfmYMnj2t3iGG+KwSLLjWt+2zrEW9
kywFkhZxtUk6A4VKNJfiTgTbm6JirZSJxSu0xSm2e1gStlIEG9fRbfh2MbD63QUJXoxkz9nC56aU
83W/YFXmk2q6LRFOnuHjGGaWFNSOTIdSKG8U35RZslUveZEkhq3wKTvlNU23nh4nrJatHMCxM5or
5S8nvys2mZeHjSGYWbTyYBnTM7VajnPHF4po3Y593Qxzvt5iM/79ATTsZ7cIQqF7tk75Ot20DNdt
+YmAM7SNR9aArU841xbfRGCXYKaYggBWe9kihe/hTjsTPUiw6Z3cNCr92Zm4E7dBED9frtG6poqc
a2Xic6Q/+365/K2/n0uqn2gy7v4qpfe0KtgFQT0PupdmHicgbIuYph5PnONooL5Ca/rG3iQuEVt5
YFzkei9OHlTo2aVVscfHVHU3hwzo3tR7pAWEbPNCXpmhdI5QmnoctmLmZQImrJ/AoGcf+IdEPbHT
QCwCFsom40fMIjRm9eXajvlNy/d7F5OjLaWzo6P9rmJE93e6cJ7Ntmt5tpPjhDDvqbb7rXWQ/6cU
a+HBkSbwHZtXruvfJijFzkw1oCIithOAT4znwJ8DCbPddRiSogeJ4sakvuO17LGcHLJ5msL3tdTr
bhhJrYiE68YscNabiYOOLaHr8coJcQHH7q24Mfew9NbzBmlqfBKfS4vOTVIkFWCvMShOj061iEg1
gRM+n9k8PUIrZZeVByxdvALKre65Mqk5Wk3l0rAqWa6pU4UL9fjq/O9mbwViL+xOgK3DAlfZXVH9
xLbat4AbLJ9gRAx/dFCgUwLsZZnoKFQ8IeMDK/gMQxY4FywfnfrXFez0GUr5/JZwYrPVMctP+RYf
4E7UcjqY7IpSYEdRjhSPiV9x+WoiWfhqBONC/Jupq7I8R2m2KAcgpOY3C7vze/SVKn3Jmg0GjA1n
5hW0MbnvN8FE2vYGIU32Q5bUR/XP5Z0ukzN6/OkK4kj1RxDS+cndZzJ+g2Zb5I3KDDRrKlOjt52b
PDFLUWTB43jWAGmT6Twu+xfGOjNDZT7DNctEiNyrqULgaOHjIDIR+ezzY/Ep/z5LpaToN4ddzw/5
isCbEdfb22XyagvK54xLdFcSdavNS1S7R+2vgpq87HzEQQGYLTINMGQUdskrPtrM+QRz2Yq0Pb1e
XOFHlnnELiw5DtJtBWZJ13DEw92rBrqKE2IWhg4QnXRdhGM4ldzTpShotynFHQt7QJGwEh9VxDV4
ZXyaqqA/V7CRmYRBQu2zSePRIZSfwuH7vITvZeM0yliUuZEB24/iShVDZfgalhDT3QX6okxdChEf
vGGMr5y+y7bKWgz8F1dQWnI1GukRvoKKVx56GgMtCZLo3VfjDi1FVRyUSGVcLQ+6mk5bxobZYNcR
JRFKdJ0wwYfz0UIBpzu7GdJlr4aZgIa1hJFDG552pwbzuShA8RR2JmpdyxSu5IyOO4W7tNwhgdHc
9Rzu60bxyoZaAji+l8a7gxHw6d1yOHoyZsTXDyqgaIAQRQTHmEsYbXdDeytbGoNKlZyGhpWy7z57
bQ1CcGfgPnR/YvqvilgzbKFN9VMf1s62oXP0y03oWXpD137zBxE0bZM7zmntn3rxNt2uRJ+yzTzg
9XvSrejMhbciapbDaBGnOfpNopkRvlJoFxaBG8RgijL5szXqQBqLkDOIpoIrMR1VCS35M7MixhZw
anAs956O6b5lYZwjl/eZw8cyw7jQQN4PQamBI+vmpkcWDOczjpzGOoWD5z+Rd7X5/b0nmGPvA5gO
UgiyqVQtHZ0IHpRMHBzA5AXqRxdKVvUY1dsCoCnfQVIqWqJqU3ZCWUgbSybKrjSlF6tFgUAj3u/3
yX/YA9Y1NJtRDnJF+k6sEo5mumNcdnvpc3n8SOVGGoX8btkbrk6i3KGAY/UYEI8908Py3YQC8rWD
IFao/waS4uPSuLqTJUdJlVu1+usmXmeuFN9CjLty5sCecaPaZKzP7wda4evTjHgAYZRZN3QCWkfs
ve9AGf3dFTIhi4ZzNYRVsVTb2dipSORoSLxNrJ2yKfZIpZNAXuGFzXg7NaqNhy0ro8lOtxWBg+kK
JOcn80QlaJjaN3nOyNVORvAp1DX0nOKhNBedL9Zci20qyDKsc0YXWU/uHLmxRjCV/KZ/CW2wM4+H
K+evGPVu5Up/hRcRZT0GsSs9954w2bBdF/f9jUX17p6BwDA0nV2zPugwX6w6rYg24WEgPzpnYyag
vb+WbdxlVGtIxkBfTnpJNUZb2eNIxcdz4j89vReMxBhmzWLEGmR3xvpBfueSIzDjiQcpV+qXLiMX
icCb4y3kg7/Pm2QXWRoPcQBCdGv7IdlQaUSdwTnWJFSBmtvC7QciAN1DszrnyL0Z2188S3zmsrCe
Y+y1oWMwcsHa4EfkZwjRsHoZH7kELb41cTVE4nBvRmcjy5aK1S6UHDt+q1KE6XT1xecv0cMYcPa5
BmywNxYXJuy17BrkZX16YqpC7aN87aEw1HeTdR6kcf+hWBqp0V4m0n9YvMXX6pIJeTqOyZFQ4xTJ
eR/eFdX/321MdA2IKHJHbIa387YPaVxNPqnYfJQiW3GPRXfuJ7Qwu82aintmoSobIO/zkA0WvQjf
52cpExwYorXMVByHYHXcDzO3J2x1c0QhNJ9Pb66O0xgi25M2vBkoGu5cDR/e4nhZiE+bVS/Ub6Lg
S1+lQrQl54Tr67XCJ/ZtzORPwfDvIgbl0jBdM0xAzRrf/FLGOE6tE2BO7SE5fMxubA0YYKeHClsE
YHZTNf8X2cDTEK1JXG2Eb7dLV8NW4xxQANOCtFLbrWH3P7mry3Vu7x8lejgGFLjTm4n1F2dCZW7y
/qdx08L+0WfT8QEMbQjYEJpPwSfvZRtO7EaTTrUplFrNWyx+IeAjjW4M056BI6EEQ8gb52zRmBQc
qV7TqPrcr2xfoFZsAiZM9pXV3y1HMEf4K/+n1baBZpGSHnKs65DkAtOoxYMDG+wj1qPGXUIIwQw/
tRtJrGVLqVIWNLu9KrHNZjpuRTuGJi5cieGtdsYW7QwNEomHaj6a6Sg1nLfyZCvT/yLzOUCp5zkO
ILQDMGMPMVnsRFTNs3zPigIGFgOzLc6O6DxPXtH37u6FWzufm2aio9ZupGkE8rqBCu1MqVd0XQwi
9YY3j5Rf4r3iNX+/iYwCkikX2I3PlzDs1URVaDh1a11wT0PK8DyIrhTujuFXpnE3aLW6B5BDHkSw
FSfuYBSo2sufVUAP4HeMnGvc2SrfZFep0MZCIUoFeYM3OpWiAWVTlhSunsXdIV8sCerVVB2C5eCv
YYpfeHvjwxuqYnjq/QFWL/CLT3kIkGMC3OqRrIybTJedzMWRebeCK8+ywUfi/IMyM+6DYVZxTW9w
RcecvrTSqVmYtG+ZEaBO7VWFeuNecz6hy5CchKjjy9aTVVy/qJLwRjTBP1B4A5aBmnhm6T/qYtfo
Xw6qOhQShWKrO/stNBpqmSkqKITAjlvuC/6jDSAjT/7tVg8SiW9aKFPZqrOaKOkSwcnpp6JmuOgi
4hnkRnGjfYBe2OtOrQFoTVVGhdJPnT79js/asJKAMgGgkWu5SUKyNr4LHETq+InLg29DzxJIyFwG
/EjPD6nnwHoqBMB+BouiOhxvLpmGPNEo3IoJNckdzFFNwIc67ucRg9JvIOBiT+iSiBps+kCBNQ5W
k1HGLy1g5LAHxM7sjS961HMFA3e/Vme/DO7DscP3X80+5yAbXCX01aVBarnnyYHwTSDZ0eVf94sd
SQkbUNTuPMKhzkz52ib9jkNABagAWJG3jxOYVj2/eR7nopz6CPBKWLFW9bfBnxunfZkl5oI96BTb
Lfzzl3xV8tJNOkABnSOw+YVI9DNAr8UQz69xa/FsSFGluy7QV/YVpbcUwa3vkwwKnPz2S2/ceuZL
84teHfMEc2s9eHPHChe/vPFV+Z/FgcXbaADTYFhlW1BTYA+rDJ7sIGnL4b3BjFYebLcKg4XKo4f8
kk2pzJv8bhQL/vA/UV3tUJkrrgrto6GNVYXgQMHzDhHP3WqbdSZi9DCZx8QuQlN1/EGqh8rld/uG
srOulu4rTaTVFw+7TeAh/GtYV1/sC+VrJ45FWdIzhwiVwTgDEiYmZwIYyo/Qv7wfj8AMNwtBIpnm
hKMjBpvQdp+AkQQ6hOaO0v/rfT6TqvHS7HMOvI950BinH2V+nO/mDf5t8KebyFj+G3LYV+7E+C6y
wp03nP+cJMj89QrSnQgGC+eI0uFo1eQ/nUVjaiNY0oSUxij4FbNIm/qpdFy9gSlDdki3DHo3CX/Q
didd0p69cFyr3jTz2z15TuI2kKQK4yOXY86z0iqwuftfqoNnu5R23YreNd2FKKh+5epS1JRWHQsi
XLYflxtjCT9ID/Bvn/ZwqvgGbpL0FaNpGjAwAHH+sDh7+F8d/B97n1S+v4u59NCtXW101+rAvy+Y
rIdRrW4SF5gU4iwSHm9oxlH7KWD4ek3BKk467xevlp8mFmjyap9JIiEFMJnFZ1WqaNGykbSrs8b7
5lFzEUkCLsg2KgwsmWhE7f8js6fTNLTejJhndJgmtTknJux35isDAYgn67hplyVgRW0hblk3uE27
ao1rcEF3N+EQ+mzIUZ83QAsonXodtj4L+29h0p5C2ItfU+Q4lBOmZaXskr3y3D2rc4fZciycywKx
JnY79z22H8PVOdYPEam9L06DsNJKT81/OG8qT38gaQfRcI1fWg17byngxJUgqhbLgzZlB5JmoQJH
fz3+Y9seJR6RLPKTEutTfUT6+BMdIqBs6y0ljGnQGSykF40q29tSNx9nO1fe79KV0yLqWiewvMYW
QBq6ui5zl4RmFDh4wtTE4xjQOtZYIlzooCHqw3A0iqQygzQl/Q1J4UjoqxXQ3gMSwbeVVfABffUN
6zrVFPP+ngVeuFU+klNUdXgxm4/JQxc2zVCpmTvTa6LebOO2Av4w0VUiPuBi5uvOlM1hcZafpwMU
cUfxtIo1rmCO6VVLaqoaJVXjuhmRpR/4DT6XmQOS2sh6Xpv8NWzTLNgyr7q/tjf4UpZos8y6OrEZ
61fuCbLoa8nXBNO8ENQSzGOOX7EzcyR+N5WQ+uFnKo4SiY5mpenxBv0Qi6jHWfXtofXUIJ4oAAqv
DTfhFdchV3iGsfim9KEhnE1Zl0DwvnEGcdJ5vzqWmwDRschyE15gJosedFOyRmVJPxY8Fh9qHsOE
LEpEOm96VcKttf2EmGM4P8qAEf8fpcj1Zzl7FhrmO5za4gwrZe0uZNCkbr1J+hgXkUw7Y1knhwMD
iHWiS39yFosf+YeqEmiFzXymxm3H2oIBxUIRRWocWXm/QO/A6I+aflg3An/mjitf40QgYcymoM8/
BmWDjHi31aWQpVsfd1dbN8bMvFQD4jqWJMQ79eVxiBCslVQKPYXZkYp3mEb6/soyb/9GD4mm5Zx5
aSuXv4/0PevzZsO7jAJ1Yjdvle2VRW+8kpCmBnQIfs7TB3+/tSqnvr4jRk2C5/6Iu2IBGYDLHwBE
mBKNoT3II3J5z0chNisfWt0jxI5Ze+USOGgEpo7OUA+j9Bl3vbSvMiAD5vKhFut9LWY4r7HmkuDk
JB0cTBpi96L7NL9L7cIZPUUbEeHBt4ya25tBmtA1sjnx/Ks9D2tki413xkdfayt0VFaiW0wuDa0e
B2TRHj4N7juiTnM/O/1Jwlg4eAKN0SoF5wkzxN3/Oajg5aWsYFtk6wa6wS19nYqWW3rnU5duY0nn
G25O8h7XdEmxHkR/neFNaja1s3VYVVTtlnoUdbrBDkxVjZpBDoD/3Tr+cRK+3K+J9N0iuQKgJkQF
s54FJ7G9t33PL6D4AnnPoXFTyIWYhAExtF+Z1NUdLud52BjfPi4Z/xxaHj3oDGwVBY+xFkBvunVi
LUBXW4SfztiJgs/TyPOPFEdGdqA2SBWU7bUy05PwZwKvfwGQp9aAd6E5zgqHIFWz8oP1E8p+W6i/
rhx8VHFND98bXzije9VXTreCLB0nr4husdk5mQiziWjudXhmtD/deCONtF1be4uJVbBGIduO9Z83
gBtyKAEfvFQu5hq1GFPG9wKN27GScSUenk2Im5GWEzti39+B7qgMOXIHTPgEbmVQm+nUaoUeyLUu
gx5+zz+Ij1Imy8sdKAmTPGzxl7YqPKlgZqW1WBVZmm+TEjJv/5jaLMnYcjOSrgsKExh9r785qZNk
BfThTxRVHqPTAodSu5Y8uTP/d5fvggeC3T+Bc9EJI30pq6QEapTHwMdSha7yShwDjJd1gFg6DOKq
Twe0DPttyrwWNkFitugk8hSrPdZCop3Na5+49crmtG4MJHAcLWZbOfw9n8ZhdZXtiVhpI1rOb7rN
6lhssp/dCZWDWgFlknGiP6hOMraq3KxhK6lgA6UW+ivL1dPpow6sG1Qbx4mfifs3kRirSYHIVHXG
Y2wekHGL1xe6s1Sdw3tc3aaYw/S0YqBo9FDOKCjnmw6KZZTw1SfpcrFiCPoaGUh6xEWiB/h7YlrT
ZETKl3LDki6WbG9cUFSADRcgFvQ3uyomngJ0QDymFu6n10FLkJ10yULHSkH/77/9a4PfK8NidGZr
oMKMS8E1OmQ0EiaIz1V/9TWeaJOjXTG6e3Ahmh8WPv/FpsuzeVwkLlZv/5RMY0AkBH5Bk5S5SW35
sPVeqlfBYzovzi+h6h5ZkL4jyxtYxUef1OBAmd9CHvQ84hkDjb+PX3UZZPYvfhSg45IhvrG7Bek4
YUm6h+lECkcq+vt4ILCVNSEr5xeinj88uANTGdWfny2radBsM6ajz3X/l6lSgw85gH3bDmcyi0vX
SweMjvTcyi3p77mNUI7UtKZXzELj1wiuYUZnEJaz1wGb13q4yVeSAODnNyLNqS4c0+QU4Nde42wA
Zjk92UKmFpTBE/ehDjkAxsY7q/X/Pz55PCFvuEqjb+CzRbfyGUhCUVt170qo1JLiqwYqRU5Iqojy
3IO0a5OZ35VNNnwnSyoQ4ZHSqI5uJsJGTuNvignBvORCoJ8Up5zXQHClQ3RIiHj6ACvGH7/Y+ICl
uQfOh1zKmnDgp3+d20FQVjL4h1CRTwjnF0JeuNOTFBb3pVH2N7Z2ZeTTNkY4LTLhqkgS5fffbpZu
QW1OP3A/IVD7Y0nscH73G7dxHfbd/EW6AEotteJQBUJfdAKJy8OVmbKQd86/5AkomU4cTSUIH7IM
dDY1IuqxIg2prG2H6l45E2GCJCjxefObVjL6uVRs1R75YY5Lndk0ktIkrP2mmfAeDPAfYr+g2dRJ
kXI8EdPmg29Qq9U+TAyefIfNKBm3Ztrr7Kb1Wgk6J/8WmPU18Y/uJRKnqcW6PadErXkyQjYnYSQJ
wSNHJ1n8063+cYahsfaF4BcbMdeo8OaDvTLq5rUzTC5yPvsMzSNrm/yH7WUQgRryuN51fBnkQy0e
XoLDpjDl7pShkMwpNyLWHH4IslpzkXSd8SExwmg4KHIgi8abo7lWnUC+li8/wmOxl7lybtPkJ/bJ
j+g2EZayNY+hLu7PMgbPBMK4nSJnit+dpU1UYVFLss6qMVB/Uh3T+MfG7+xYH6MIkoY8ZVd1+B4V
WGPGQdopok7+6/sjqOIel0lATC1mD4BqHk20Vz+VWhetW0Rm8u9PLVKv3kXwMqf4U0hXQAWB55wp
EhXAcDujJNzUkIymuZdzo+qzHdMTAltanzb3K34q5YmlMfORCgQXbZt6F4NaIu+InD80iWfBLaMJ
Vw/FMcRtOJkm3kmBcUxfDjEHTqpewj7WfZfMgz8CzRQ1KT8pwBgP0dGnPafIyTDQ97OfXygH9WR0
VUj50FgI6A82swTU8wWkmvmPHQyBBIpuocxTg3jwdkx0uZZUHo7vRfN4A0FEfHPD/xGiSOUU+rzR
A3BrMQQ1a1/HwXXrYMGomjjgpVCYXkuaj+KBjv+d3sidmj+hvc/adm1vJldM7AG53Q6vnv34+FMA
zLYajM4qGpEWiMz+yulSuv1sZy2dtlD1CModMzEgJFESMWCzLZQQSEm9SoGYB3baXlCyph9o0Ctm
D6othEin9b7UEIys+iqvb0c8/jjP6KnsY++0uakNsg6kT44vdu6AGrcnQgbl8jHVv5br0hDDLOrU
lmc/GXN7hvBoIjx2LQJrRia4phnjX/SJ1x/N0ghzkCc/m5indSRiyIqJouCEUt7Ltyxm4AjmlYOw
XZPpsqn0Zpj9Zr6cYnJpmcHwJMErUpwP2Y8+xUlkBRML5sH35RqO3eQdcgzgIEc++8WzAVttJ23A
xJDqlj4hNCoDHvPZOBrgnr9pjql2IU0P/wmHoh+OXFebt8tZLJzGgy4bt3z2Ykr2CHEQQ1ksHA2+
AuxSDf7CkuJYdsBNNoyNozBEgLMo/fB/Yo/HZ+DBw0etsDdh4JW4eSMzRcdaM2Wydhoho8lgJr/g
6Iza1edS3em2mGDjLv0r2G7szlSp+M+Ld51bIrVl+2VfC6QqisK3rxT64yi1VZw4hz3C/C6HFRxr
5y8jxG8ISpRailPGB4O3NYzuhOrU3o4p8Dpx81ImO2VFKVu6cKz0peRJlCh197NnuqZQtgYT4A0B
pW5pcfp5J5xQhmUQN4sPxhYUbm48UParL/bIFDXNB0rO2ZpXRXZuZr1gHFpnjnUprlWUQ+X9QyU6
eIh2z/LFPeIKdQfiQ2WB/03LxNQswxCpOjEvRdS6oH9mSZcI7AVacUC/9i+TKwycjOiA9qF6rrX5
NC/1wNpcW3dlp4Zx6zWYyICWZY7mRpievHH7HHHhaJjVYAmJrxYjnUTYf8ruPJ8JZqgw0D+lM6/w
nhGSbYFBMHKv/f6Tm6HwpdiAIM8EZmP6+EzsI44ELQXoDF2p4wuigM6WXc1JWnQQdAABxa28clpX
Y1ZCQ0XW8Gsp5DKJDVNPYxbKX9UIbKMhLUN50ymp52D+az9OWiBvPl+fN/BoZy52tl8IuNRsbvnc
cgDw7dfajSu1COf3pZEy39H6q6Q3NiSa9LDCt9J05VI2aifNy1ldrXb2rIl+BAw97FamfveMPDZP
MBQn/6NZdiDU7LA2aShn8Kcri666SLkPAhrzhXN+RrVDMswh+ET46sBBrRwy3q4XpDe9PsN8dKvl
N43o9O+ymMA0pdtiSWmAmWvLW/LZtoPjPong2Evj3hUOVD8mMe4S1c+Qu0bslm3kfw3R3knTZ1Z9
mWwiBS/Q/LlSlLPGL+9++12uOPOC40jyRJENDtrxLA6BDNqQCcx9Sqw+Jlz5ywnjEAr9PLzR0T7Y
77O4m77/GwfD/qqEtRN5T/e3jgpmB2wbyzcgcUobRyZbq/pbmAqtzCqjszN9lZHiqqmMtf4xGdrU
fAQLWTT8LvTZ5Mssnz7vYqb397JP+lSbFtcV+unZ4TIHuvZczfPQQhG3BrR4FfXzs3pRPkbYfZW7
Y+7YOvw6ELl7Ucb3XR2pZvtReZbDm8WRC9jnmzouaD3rujh3jRsFO3iPQqb5XhXkW3sf5kxUXKZK
ggyea35X6B3fG+Agfx0euwUjDdLlfm1dSwZCSbt25knOwfnWGlFiohuL+K9jfX4hoP+kL+L2BhlS
+ATpf4YCWTgBYtkIyzcAzyRG9EQqT0kdSfabLg3utDn8eVpfazdRJazNfAHDIZPJgnx+xH462NUi
EW8FexeQ8nyKq3TG1e5D2WPNeTLlurIClYUEH//xGRnOmJ/kNEcKBpwJbqK8CvBb9aBCzwiPceH/
9fJkLGz/q/Rhhxe+p0e1YZ69fqjG0mzL7Sz2TqNowqve0o5ID8fb25QiecuJbyEdNpv/OqjkiFxG
CN1oPU87L8K/ZZD5JPnSYvN23ttS+TNelUgHV7huO02g/yOcANP/BYAWuflAJRuJweSUeZMJsvj8
8dPLVJ2OSpZT047jy0Zq9aS2+ppzm1+OoS/PcLZcE01QCfu+TcL1ktk/zsoy83VFXY136kN4GxWl
JN1r1qgSBzOOZAXEKdtzvd6DEndrKuE4ihqpbKzgSPHol1ika8bAZo6qyVPFiTDAZadvon3G2Jt0
IS+6pKCsw/btSRmYE1WpZbzVL+5YpYo/NjbZh/k2gvdDY6ERsPGThrBUE5u+FxdbFbgCuYDadRDw
KH4hsB+sBWVMe+H3AdpBluBJG5+nvvOXcJ+iCk7V/H8Uu3LdhngEtuQfMS9fA9g9/yd8C/LtA7Ns
xfGlrgC8e4h/PfJYQwWoZNKswYwFzuHUhlxQNgCPsGXVktkMHUICa91Y+g42XOsUUWgGyrUxIHPF
zAXTS+3k6WFPoMquRTnLJWkX1cQh8H4iLdbaI43CWE57PtVO+WyiuVjrlmnzLowYWHh21isxGzmK
SLfosMs5pkxqcTrC4XTD+BfgDdywK8JlrUY3WIvO9OyXuHkOYwGlXzmHB2Fj+87p4ZFJ7YU/YEap
KgakEbgVp3o9P1jSAi9wD9PtJPKTkH/yqlxo4xu0hAkS+kgCu1Mer2SzuAL8kd6t5cNMSzO9ITpw
EslhkX+4adWMEQ/7VcW2VBU173clp9zQBRr9gr8vpVrc1p7jn0uQ9mZXPym+9FQsbmHBjFUDoDZW
d8fgoYXK2VaLwOqPIJ611nC+1vQvcInyeRP3FOCEt+80pRDxXtZtdlSZtgIisrS9JPeFQ9gguW3q
qv0OHPX3NgN/wLY8lQEsuW8LRb7iu/et6sRLjatYeY/BQreI871pol7u4xRvKOvQ1nF5kgyHldJZ
o5jh4rWDaMFarVqZbFnPLpbl7DiVqA+bgc3qSbT/stwUaozhyuvAJsaUvH5+t71JPJjn9b52KSDD
KbGwN1unfsvWQdQya+0rYpy735U8cX6fFcAaNOfJiuVLGnX67EzNyQI5Tqsk0QXPSB4hDrm5oARH
0LL4Re0PcLLCypMYKZwx2vhlTN+FEqHFL52iLsL44k137HbIRPeBfvnRjpIA8g/21YCdpxLkn3Mp
RwicK3RijV+5fimep/YIt6U3pTY2Dsnw2y9AJJjIuoOpWoGvq2cNXliKpvYxW2nOxnAElhbWDP/9
CYSc4DXElIglBtrqcZSNd2MOfdn0XvIFW+10qZpypSnYQ6F3p83lI85VmkiH4wqQxVVR8XqzNki3
7sd72T4XY5WzUOp3FdxrDJ+yMcqoV3Y72NZDcywC2JRI/QqHXqxU1LNEHCgrAnT02K0wYluYVN7u
O1/XUUXbu5Qa4c2g6A/qhRKGmaujZ+9UgmkH6ay5jskGG7uIfw5/Y+4ai4WpWQACSDa5KYMH8vWg
ihHiWSriCno88UlV8fleyC5t+gANNcvFn8uaPvoUubYG9+w8dQYo+f9ceeF5JWxmf5mU1c9Ryw1g
w3tiu1f0fhtHXlYDFTGZFl2KtkIpb8Ww5wrhyBkshBy0lUIKqRypm7ndczFy+zlAnratpONMaf7x
ePqJkOdTSRXFiVdjYc98r07vfEJVXLzkyDdoxNgGiU3IC87InHmLXFIpyuqqR9w0Uicm7tcAq6y6
pMAG+Y6FHI9IChX7bzvsZT0RRRt9n4Bd6vJpEX0nAcEbtBBBjMwXngJF3AerETnMszk4viWlCccU
hPn8QDqCx61HxMIGFxkE/dJBzibF15aad0nCS3dq5/7RJlqWnBjFTnMX1iZJe/kBCaI4QtieXeXn
1fuM8Oe6AHgf3oFsvGJsGP37r/Qn/w9KIZnCUK+dpU1JcFge9VNJUf888Ym6xPum/7SMr6o8ly2s
VXaK+jiIHg8l+jkIQias2a+phnTek+9ixZXRNqezGtFO79bu4zKYC5JwhronQIcHrWikD1rDsQQx
nrHxfA5tbf2mgLA9WjxDaQdP6bmkToiDKIBmZ6pJCLCkqScrtFLSRSX9yH99Lekn0CeuERs9n8UK
/2T526PwHiOk+SygpdFF8XYLow75xATJ6P6sAo8d5M17/p89cHLXRsfqCM4Qy5tAPO4InXRYq7w+
RpGmx7qvJlBdxpaWiIoCEqBUL4UkJ66RawB+GXiUV1uAYK4ImYxNTqWzoNiICyCp9fjnYUztsNJt
IdzgjdZP5h/EqpNnmhzMR3L6RI0E00tXBEgz+N5VBsd76xy05154GnIKWSDtlj4UWJprv+ESBXzf
dD5/60k8y9TiyBaSZeFiyQ1zmoQ+TMpOLq4ahDd3jTUjABwGahshbILweImjzrCRtXN0IH/kPMVb
0El6RHsEE1VIjA7AqfG3MpC+DRzLeRT09hC6f5PS73WKJ8yC1FWVpuxt49nYccc3OWLkPLK5YX0d
5DX74GPZZURkUXthBRQgIySnIQ4noKtCKJr3RjWcmNd+IIhKeI56wVjPQznr7MOs3eLszVw10bmX
yhevenCgWNLvcVWFUCojBkiWHS5dpFMrsiCmW5omcempBMHf4O/274qybXX/ChZkvUBMnjxRH4yn
We2jUO5masY5uVmUAI6SwWXnjZTsNQE31Ds+Q4wwB7JGP42zyy0z5CnjVKzeHpPACubI30CQBJ4D
h8Bb0Dl3gaTTH8qK5+Hh60KO2jZkjT+mqedNCaXwrliGkNtSQstM815jLgwtwd4Ca6thTGS43y8g
fTb6q7fXpKCFpI92PVQYBkfEKoTVK4rHQ7wQwgAkze3KA3FYNNp0IKd44yPt1zHJQyUesxxfcvdy
Mh9/Qs3krdv5JGTAgoFFGFSm6HH9Dr+t+VcuklUOvE9MwDKC60DjxZgHVYv5H77rk5C3nTap65wJ
db1+P989W25hx/JtR4uMxYBOwnoC6LB4vheeKd3Fekth49lBe698lT1IuyxmuJ9tIadCFCLubOy+
VXQlSPqADo0/U+bGqqGoalaXwV3P+OonsRDyCS3RNxvWO/KWXqO0ow/RWb0Ty0+LA9JDWWdBfmx4
24avAznGOqH3Qpc1jdLJX1ImpZcbq8YqI9XW9TBOGJXcNGsc+qlBIqjUN2SS0si9e9I5HcSDKBPe
l5lJp4vuZYOxAjZx2+L70DDVYUAAbdTWYnrX71wNxUoyA5k7BOIXQjI8JPsL86f+SdcIQPq0ta7l
Zvxd0V9SU5BCStFULIIi/i9U2oo7cSalWV3JVJJJOdKV9MP0453njE70NrukHnqHB9lV5tuqOAir
KA1fvGHTIzjZEqjT4pcVeCMY0Y/VgeTbr5/HW/t13Jw5IVSY15H1OicdqCwy+Qdcfj33wgMlWMxP
8tZSb4Yks013TjjX0uIYS+WHlAO8CrCTn0IC0lTct3ce7wOdBZHZofGoyesuw0806e08xohx/6IG
wCpGJEwvwa/TsJoi7dveqNsHa13fGjmoTxDhViDW7VIw10E2mcjnIU8vKTLUhns9GOIdk/9LWRlw
ZMFnpBMCJJujSWjgdGXxCiHux12XEdwaHxoKWzi/1cbJh46sJprjaZx/G6E/bP51KBC3ltz2xnqF
SBYaG2wBAr+cNHQZc4G0EXGFHARDbt5FUTfD0SzR7OHfxhnXNxkmbefJdm9GJel8ri3HmP7W2jLD
N1C8F1fZtm/cNJG1sm32DVh0e/rCjK8abBqQSTOp3l63kF8hzuQIDJcU2twHHWiwxHna73Mi9R8/
AwOYvwtub6psUNFXLg4WOclRMTRqpZMDqvQMH1fFV4XPQCZNRQHOne1MpVTIFbwo83R1Y75S7j+h
7HyPbwXQQRyoBd4uhg8mNE8W6MrITfJv9zUzY1A2oh4YMOAF5EK2+2aVgmX0ZXLY7DD0glSJpvM6
yB+nXWKfl/UPwZoSJkzt+/oLRtLvU0OKGjJrshG0cIIleWSANQh3WMoSJTjw+9hjNH0e8WddZ3Y5
mCqX9MHMTBae9Jcy/OfZxc8VF7ewyqXJniCw/OEX2R/UHp/dDxqMfZN0nHAU2FBiDjilpUT33Te6
MwlRmZN8LE760z+sZ4K732zJeDI04lm+gvhJF/DZaKPrGmHeLz2o2ZEOwPoUkSNzlk4vfSn6HuKI
qpqyIE3nVTpZYREfwTcd1A/JXAPAtZgNWKDeQFVSA0ZzLOryg0XqE7MAIpG8oWNJhifY2jQ5LiJV
gKD4RDCp0cxGLeyq49WfC1pMFjKcRIJY/1c1jI8Nb6gPYwqO5WvlcT7XKhw+bxsdswqOgvUmZDOO
6/rEBLEM/DEXwOECvz5HnUBLf9NJdLpTlBh1ZHKlWu+Wko4gi+QR/hs2wdlW5QaCx0OmeAHx/QUa
c04rXx+utDp+6U0ZIl1SJ+YGKNhe3xW6b7C9Xyzdy4xQOofrUn9XYnu4hwwfaIw1x+MhJDaAj9L3
tuhKanZ0MWR5ZBlwkCsLZcVEUapehi5j+Zz9NWdcoAKwRNCnOuh0qDHinAY4Y8FpzXloGHDD+R+l
cKQsZOy0+2YL6eO9i6D/4yS7FKA1fY+1lP2rK09woOumUk8s4Qr5YtGTB8WH85JcdqDe1XHyoxeF
3/poaKY8kbwc648huUDXLNDmaPOpbK0ITtTjEozbY6UqZWE2oWEiVAdyvPklX80bPukoDoDwfn/9
7QfqTzSw93cV7VfOrlYoffIPRafCSgtng/ZsI0jbvR0AGP6njlrP6rrDz+kHDlxfYnPfz+IaSwcx
YKtcSWyNpliPJc1/Gs8mNzWGYzkMQuC0/fDIN39PWM4P99IS0/wITvXFw6HvGO5YnrbOdxkMXwGS
gjcYQCxD54SVSN+pb3mLYFGBKitwcIsED8BPmjx/ZRN0PahNV3zx7kp+ykpm+Lrta3wEiAHf4i6R
BMke2YbL3bCkUL0Ei/Qy9iX3ImZFVpslEMYPeMnDacDsgcQVXybXjp2eR+DUHPI3rkbRhez1OzCS
LeJv3/HxwJuYSq5Bix6vwyg2AOqOdJv7Uo2ycmTBa7Dk3Qf3sLbR0kkZVXGarNqclC3L9Ng2gtWg
OKRPi/X/XJsTGKOWQlJFPwwEd2n6d7Q5wQofvEaV7y2R+s0am9VCKM13kf9/1hiMrhdtbpcW8AMv
xrxR1U1ERhjL3A3OAN4dq32BDg7pJ5fnVDGW5+A19ZraJBCuJk1J9stVgO0Chvo/u7V1nVnnL/C2
wQse4t5G1jkiBDSuAxwgWCW7AREE3q13BXHne8f7rhn4qcJDOKK9NzdUxD+KpMa3NxwMcqya75yX
aArSJo9HP4FrUDgZbnTnnt5phIo3pFK6yM4buZ1kGAzApngjBj73r9AcPm+MHWzi/m3stNS4Bp2e
r+M0MkDYmQnHpXT0cT5sx2rJkAZuUiRebDyahIu9MU+7/zwK4VyKm/zaHwiSYWVgrTWpc+7aqrTh
LUvH0Ugqwlk+Y87P0v/lgBB6szJUsFMd07CiasEfrVmuQ31YikijEb8irDkOm/GsXcgkt69GsE1v
WX99FniUsrUbFqyQ92AidouhOKk1vMk9Uxy7OalETLy8fU91qG4hkehgbBn2AJHryS7U32cboAaa
VlpF4QfUNUpFsoV44bmuDHu6fjZPZpsAL9B/YUZB6tBe8/VLWizo+F6sEqyt+x7OHyFLZcem6oCK
vuhbmXIBifSgr5QYPSOnIcS1+f0fJfynJ1opABE/wmO6pHnqGqSW4/UskgKl7YAeUR5mnjkxdiKc
W16U6x9XfcQHd7xNICzmFDC2hMriYq/b+h6wUfDjCcdFqPSmWt5DxQDOJa6Zvb06NqZ3H+ovto0c
N5Dn78Rb+0C8jBipxVb6DWWaOrpYzkUvi2l3zPtiSyEgLM3MFhxaLEMeUyM3KnzEDU1mkSiBM5od
w4F6dZycqcxrUmzY+XR5A25XWQvK56aeSLMAN8Yz3Mo5/cl4A3yBC9VuRET5hxfiH0iwZxdRtoMc
0r2BMTotuuworhtqiFODZs02/4nNheUcVQ6lsCUJVdUlAPnTAnA1mz4oV8tvMY6MqM6RXnlFIfad
LMvO3TqkeiPpfmb5x92v2Fh/rFOMw93XJJcSi81y+O0HbMGkqoAKNybbSXFji7qnNuU/BSl9clSc
TaqzvQayEmeDWm/1ShTXoqhDmuuNic8PiSS9NaZJ6FghXO0DX+5UgJknGsw4p9zyI5Zm6st9NIkl
5Q1IZEg4YFj5LFeo/h8+R2Z+m0bxLrnk6hiYe5LQFFeZj4OJszgzuESwg/qV5LdWsVWmHp+78eN4
Kdh8v8uH3uj2t856V7BtYxsDx/fXjeQpqCOIsmaF1aKxVNjQ2pSx9lUy1RsnMsRKQ4CBmjftvZ0U
XExaABrS/8LSV1HPB/15EEAim603YGh+f+PKH9wXl7QRNbSaigyWRp4mxw1n5T3YPw0OWwWzr20y
AZKWbCJpAJez6trryEWrfpMXTGVj/hJkaKfPxDUT0Np8Sg5/fs/KakOzAft5vg++qaTIAc7uvcJw
ZMBzsasxL01BLGuEg666xDgb0KRQa47CjpFqr+GELXIRyzDdIQbURmaNJeo+KsJZ/2kehLEVSu3x
XCcigGA4rn4uYmzmLOenoHNwwCgb7xGsSXX2Wmmsd2+3+VR6PU2tYrapa2Ml8s+TbzaKaix0YIB1
YNJJB0xJ4vEEThter+YqLdRAdOzipsPnZerwaZjy1JDNhHhcuQAwDtM/ZVulHy5KdKw2MWHdH1S3
xZxXXBROgKauV7c52ukBcUDOjPAjyefhJ+JxSrxPFO38Fc1vURpm9hK2RgNj+CP7sZM/SISiQiw6
KiV93erpt77oD4iZ1x23cvr2tPzN6cA1ka4mA2z7JcHFo+ueBIUVL+3M2cJruRODACQefTLePRNY
56LL+zSZILNncUOo1tsn75oJ6uxlTH1FOcb5pv/ks3+ELBSqyLwdYKzn/4UmTINWWVxeUmilqOVt
Xoe7LV3p2vDmg8DOAY+OTA4Gc1Z2AEFIgrUQdFBfweSzjGteImOynXN6audXU2KuDDavNg/VqNbT
Udx0y8jqIzmIQRM72aSJcTnls+aDVFEmkJKxbVYOQZsj2CQSMHxVNQL9gC532Ct/sZLj/78kzLoP
bTHMDYn6GhwQvAnktwnND1znE2Aw4VE0sFb9j4J2MTzWp6SvBDTarbSInPAWVvptzwm5DshEjluL
WNgqELTxo0MEthNx04W1cGmnnucY8CBVdknYYT78e9JFvPcGNjynNbAcwLRw6H/cw19QkfVKBw5A
tJi5xR/qQjgVskxW7eEIeOxRktjsrxznn/LQZv+FS8xLeK038UPL+4Evuuc6Axpuer+0kiOiD7Tl
8WkO678cCqHmbxz2mWRrXC0b6xFNhpF7k9zPRhs6RnwPfTb6T1zyW6GqjEeoqSXBXcKClcvTmnSc
4kupZAzqMRtMsn3VbbOMc3ByjqPNHroTxo6F0QDSUpHOxgQXMupXnWg0BG7BJYu/0Bl1diaZibii
FN6rJTZahqK7ONHaKMGPP3dcH6xkeccJQGe9GKzp4VKqJpGlauBZKZlt6mKQa2uj5Jyl7fldZg/7
4QaxKVRByf89xcb+13IeeBOaHKx5gntIgoxwcs4IXNqByMa1xeAeZ6i7EOKqFFJFMmjCUYcdsFtU
oxhuabccthP14Ou4M2ybUdBrqpHgTiAd9OLofpkcpRudZCeZo8pm+P00n6sqnVC4GY3ytjo6doYY
n0dp5iPROY3DA0GExjKeSQ3UWYYtmH3RVR7taq3NY7RjRQXONZb1VRBANM1cBZ43+C4N/X68NOfx
AM3hc0MO6Xh4AbZO6s2hF766/3DS9guCuWgEsliO2EgkPaibu2e8a4yHg5LuE88DbEyPJb2CORKV
fSwE+/4ClJjOrL3dPOnrSrF4tmfPCbr1nqUavyrjDQATs37Hyr4PkR7HRIFyYA4T98C4guYJX+BS
vQZBT8ycNROO+Iw3rR4BM8Gy+aNlbwvZB/jLpblz5le7iCzvvKVH+sXMiEBRrC3uQx6lKsqd+0qt
NW43slDdqHm3s/MAVs2LqZmPLZN7xK+T0rduyWV4XHmWiBXhrqF3q7iTFdjqx2vFQKdIt/JXpExc
HoLiVS/nvF51NuO421Cee/heiPy5xmlAgHxqfukF4UHOGQ9f0M8RWnr8o2ytt7I1lPBK45P/fxeB
pXuKZp44i6Rz5UtBmSYT5A+1ecgt8o29LyzVdl+fykPZ+vj7+KqFLpWST0d3NIxh0y6w49NuejuN
zex2n+rENuayzAvelBHKj4qSUKdgwZAJ0rHmCWuHk/wkvdFQ9c59Ok8goqTO+fCPOT58/Ma13sWA
hfWt1PD+kvL27iad8ji9eXGEw7v9NNnZK5FETBZNEsk3SjeP21wS8TMk4xEDMBpu8Q2J+3LwRxDX
YsDvjpwsIRIKUbAJQFEJmo1/OplpVm/Y8h3sRKKtinQOlgTPxMt/MhrzxepFmILQ87dVCEz1wk7+
Znchod0K8hx6rfuRMVF0X7fIYissOEU4JuIvk1o6o0D2bXgZG6y8LvVPEt/LK3pamNXaX2+N/0Ua
3so+onGG/TWvof8lofoyBxO0lCB1j9UwHTfAljH6PKpK+R78VpQ1xXgCx3vqOn/Zva/BjerY+w7q
FIMntlTxNAUS+A0EZOfhjuMq8DZN8hRqCPwvM8+SxTmpbSPSOxh+JVLLgBX0UPJvQsWFenvevCuz
D/u+0p+/ombZUOXvyK8WpMVSxg7TDoJH6d2djaZr2GFLcUIC+GVTgETrcAZ59PX1IihAwrLGbdde
sFQ6vOdthmBA6x0Gn1mBmZx/8NnczwQazhXBSTt/cBuqJ7c2DqTN1cOZsWcOy91Dz8gE4CjKiPH5
OLtU/lm4j7GpQaTP80tyPD6rUFmNvWIJs8xy3EnoiW7wjULBPkioTxCPr2F8X+PeVUYEeDzdO7za
IMrbHVE8a7FwjkyR3kWoeP0au+LOYOSaIglhBU9o1xk2TcfcxzVstczNIHrUwc6qDHXsnmZKYNAy
LHsY9ARyILtB37LPBxgStV/sCp9BBrN5kwUwuSvQa78V5YuF+99Nza4UcXqgg5Qt1haoCFEnrcx7
5NvVA1xB9ua9ipzXyCDbz98s9BXDwMrJqVTUGrU85z7WT7trrXCNn0LuNyATVxgMMD8rRu5Crrae
cClXw1cfxg82tT9A3Y80aSRyWkm7psBdbrWR9BCRas8mSxFcEM7a0Edrt3Clpf4wbfL61SkCBqDV
FJ7ddhhq2bedkjJQlYUQwB66/hBIzTr+k7fo6i+FQuVbOyxps74SJHdsRBjI7PbIZ7LqeYuIXjI2
vlKl8/cb4lk9Tg7XlMdt86klpVG3tuyOEYdWd2uYPOFdptMYlNHv+Sd6/POHP/bxHHYLaO37IR0W
lfDK1hduC1zp+qxs+/4yEWLXEZTjNW+J5SVpJlCEcsVGIKniJqPtoL1vwop3Z86csA2urafcuy+6
04Nl01G5PBGaZGgLvWaoR3emdCMTUw/yXJQTwKTWKcPPMJdVsnOCt1JqslI51JpLDm/3cyWYEjuI
9j4AZiANy3HE0clonEhDukZTfxniwslBa1Hc0HKPSoCwA7d0cWmFXSpUdCjG/gU0Kvllsblm8BN3
5HTK14g3W4E5+MW0DKB6Fr2pSwrKzFoUq7vI4ED/9fwqHFdBQ1ZmClk27YWrvLqomsJ+W1IldI1S
xb1jOHUk5dJ3l16hzIcZsgvZP5yqQNqy3rI3CWRzzFyqkK3/wDQDb+hQ5oNmN/YZ7hYRb1likjh4
B+UPcPEC/Qx/IWBt1upUYbqDJ6cZQZeKuuBlciUDUL3YhpIZxvsoQuucnz3PnWWIKV0hDEwbDqgz
bpVL6ytYevTuxbFKgPB4fho8n7CgfBLA878mvN5jfdjo98NSukdosvpCisMVqbjzR7PGevgk3S1c
t4eYlNpeG2kXnSivU1ecDIcYw4/yWkQK4aIXu77s/NotARcqUSFkUehB89SePbvGCwKsgSmV5jJU
ImEuXwPPCeNs3zAHZjzoyD7x9VMUS45yJe/gw1+UldxD5sCCHbUlEhsxvqDM+Y2XTECUCjTPMo3H
yyFNWVD7GpRBkBfW2si6tqgvjI2kd5tm76k9f5QFaV0H3BVIGDnbVN9d0JHJjge1bRcfA1bKtg3d
DRG9eFzJtaW0W2jT3sKVJSvmq4d058Zps55rZnzPW9j+B/a5ws2woCf9v6pxfV9g90nttPlM9MsU
P0KXHnjLyutRYnPsITr0CaCdsUOBX6hrhCHarGJwuKrc199PyMtC34XjqiVflv+i0gZasvQUMPZI
Z1pcDhmGT/G5xEYTuptXlJK4HjBp9gYxuzHR1Heo0I5Roc4XjduwzL8CYWwNv1TA1pYHKHslVTZS
z7vBB0gwbZjCpLSgZe2Co7WGQvnKu2XS3DjAuoLtlszG3/BkQL8aoOusmTH9vxZ7b6Zorlzp+983
WigrxqJ3V+PvYxdH4h545dE+LwDviEQt9+5mAh9h4Wf4lpgSXS3a04h/BXMivDS+ojlQIHr60VdL
LpvEMxUY3syzpOiT8xlPFI9QyiHSiVCPbUFqt0noCYXxXUM1D7bpQPOi8S8l6iKRcoqWhswyToxc
vRtlyH1aan+lMq6uh8dWK90JjScPoCv22id6CtW+bQAKdu+kWbt9P5fFo7HTQg6tLEtrC3o2nQqG
ECltZlihs1HxpABrVPb0E4SC27DSFr6W0QDQCnLaJFWODogHd4d/82vbL+90yaJq3r+qQZ9+sl0d
pHe0YIbKKflyt6481u37+LbqkOTmwqeXhA5yaz6FXTr7k7A+rcUMUCku08AhO0GYWEmmET0aYGpO
c4JuhjwjRaJp7ibg841x6ViWc0Z5uv9NXIx6cWpVupz0pBU+kD3FBaSw9Zd/lsysokR/jSEzm10o
IUhfrHVCrAwCNPs0qrOGjelMFFwQkXwiiqu1xl6GnDqYn+QNVTBbrIAs/8MmrGDNp5khOg/5TJyn
Qi1ukFJE/Nwe/ncfN7qSBtrxSkGPjro3I6QvxSAURfALUFSVDhs57LCytXNDuLEjZNdfFeo8T8hC
Od6KU3w0r83ik0JSgSdP9R/Qh0V+GdBg90HlCWG93psYvXj6xtvNXIQiHzg8PwlJfE88XBDwH10o
61zEpTyz+o9bjnSjb4UeqrL4tlBCpc2Yzamwh36HHdiNJgRxtYItc55Lv89KV4a0tutMUDU4nOOL
VXeB+C6U/HLFsO/AHS2MTsGQLky4dkivr0Gu2e20ENJ20KLUTbDRglX8PfvR4sZPJirNUVSEyn1b
YszNtZmOu8eoR1zKuXkTOX8tDiuJtHMjE4hYLNpM03+qTMgv1MbQ/3KR5A7Hvwdk7CTExpbLWJ6/
R+ZsYKpcCZAoM0nBmlU6uixFBkzEBg5uI5YtDtXh5EAVblVOI9dhVCKN8NSbpYqTYCA6+5LT55hl
+T1PINdMNjltR3r+uhgZuIo9/ENklh94goGoN73Pyvk/agxkga0vAe61XHIJ9+wOuupVHcZMmp7+
be3DrTIaFWoLu8CPJv1TGPBxhmJKKJMAPPrqiygnfKVnNmVX2YeyXOpTshEQiTppgvXBWMee3ACb
OLmwDq8RChihNsms9Ra5p/PUGeWc8FfE7RgiS9XcxBLHi1v1tRz7dhIA9OUJiewKPcTV+LH1enqW
dD8wycmrqHNL21fJUcfA/lB1kaaOfhFYtQ20tcGDVoGCHIwkuk1UTuUwXgL72DE2Pj/OFQ8ctz3w
BGg+s3DxX3f1t6myAucS2j+u8FIOzcW1noKlDo+P2L6+qGBFzgD4zeH60UsLwg/rc+QkgK0Le1Ve
jkk/MEVvwCOZPJD2W2zDi7FF/mEp8KlxmVTd0p5RwlV84UDCY2Se8KtcORLuVjQznpdiOITDcD19
nvBZ3ofCYHtM2bXVOXDJ3+fOI7836vD0se5RFLxrkg1eiCBIpa2zY8hi+Sm/suMo3VhnHRYFoVtk
K6oOJ3BeqzfbyNKw7V/Cc5EvRkOBSY5RET5lKLaxftpI7Ry+VwDfh8qDiK1Bn6kX0sfkaML5t8wy
5CRZBqEkIFPApLsc9uQfpAZ4iN9VXgS2IpDozcrv2eaNpgMzhA7zhOL5Dn3XjYOFco6kiZci5XR5
/jOsfgq6vGkGaA3GXuEu4wiFgNLur8qjdGqjya8oDP5BYqrgiApbq8T/yNj5g5sSan/yc/0lagcF
55oZ0KL3xsVv354y82bFgOG4qROqkWH+6B66wcZ0WnhkXL3wmtuq4+yGyTreGxwkiTp9jRHsWF3P
Qoo8jn5x6TW6O7NmqOhepK/LMCBLa1Rb2ysHGsVXa4gTalmDtGqQl/G5ayXNtHSHM+Pua1CcO5Il
1rX7mCKWf/Pkr7oIe5KJHdRl3TohutE0NFtx2Ud5h4bJLEwP1eLOWLflSQRvjFAqKlRH5BSYWqRy
Z1YROviTF+2Mvmo0NLC9MWxtwylo9s8+YukmufxSab9vIiDdKzoXFizGwz/08gu8JiwgJCDhl3S9
32x0h8Mqi1em8l6Iq82pt2tzdivtdCHo3eVYCE2+e7EmczOYIXTeM2GKzmoKlV5ImGOuRLzOgdNl
rabR8/tdH2tqxUb1j/RYBty8AT6CtEAvujm+jRZkdvYPb1ujQ269WVb7I6FRrkNQ25xnTpXGU7s2
9RhvOXrSvy+4ejqyBxZXWZDKIuFwTvOcdAjiFXVMWlpNnNXbPhjN9u2LkSOGf/ZwK7r35FFHmHXD
ryX1OlP/jDESWDJh9DVFYuTX58t5TjZqXLMI9Tq+G7s3y67qrPGql5sZc1QXflZOe1DUdzwWt+Jt
mPtsb1dNlKMeUOsMgYUxQG/uwPtrcAUwZSuip19Qv6sYwzA9XXE8qZ3sRRMH2MyDUnwBytCtpMsr
rqWgMHCgzHACJ35Dbi5jwMbKIgoFddzv6p4fIu6dzlw+4rbBF8jdlt8zwYJgcx/fLacWSK+XmBMj
6ULiXoCr9gfjRwLn0HCB2m0wi/y2Jl3KKZTvChlMNK/6cjrYIESRvUndoMWRrkUJpfgFsBgggK8W
yORl8ga/SDTJ6uAoYBQSSN2eXX8m/MHCjpnyuTrvkHXHwUVLMjBhCEWAih9JsPycKBqr2STfeQH2
sfRX3F50ikwWQmP2OzUPAkHlJxhaeSIDs8b617P1eJEKPP5AqoW+AgdTCc6wN6U13+42cE7Qh0hS
wqrZikjvadXfXf7sGLKOUzPoBy82QSO4y0/ty3IgwrQW7WljKrEvWusc2dU1FnA3eRfJZ8VzO9Ya
qJnQUUcBaaLrgPJVJOa1NNxdtvJzUuk/nha7gO20j/ZuHLl5wAyfhVCEl0lvIVy4aHAYm/Qg0dcJ
j+ZSIe62dI95k7JaDPklN+iy5Pt/ldbfIZCNo/LYxqFabCo9dvz0ZTsnZ6kVQblq9NeCDIp2tmRJ
+2P1aZWaCow7nhGaMkvEp1g9/cmF9JQhFz41iBxt1fqolvLlQOo1l7GHLFDO213oRedDlN6JcdVr
OS42QrXnwlPfOsB/q1NXQGkJyOa6IU28hkijKx3CX0qYYlC9OOWrha22f5QWVmG2dzaC0fDWjf7j
FrGpGDNOthxtkQ1BIbg58qdS01sPhSsBWkIwvRDvv5f44VoXHiejkqD/9Glh5N8s62ZhHcm5yQwy
q0RhfKw83glttLOEgGdj7/Vp/9ov6GgqbY7zCylOdkwO/G9F4MsIYl6rONm20aZyWx5QzfDvr7GT
Y3U2drLycSAIqQrGuJoTT3wOiguI6oYSEvvtr66hnxzf512GnAoGYY2eLvp3tefsEvg1HBmZFJ+G
rPQO81RfxwGpcfE1BdQoax6RkuwmOd6/4hqF6Mla96u10klgmDfiASzBkYJQ7z2BPHrQMCESH8mV
8xFEX604sdnAwIns1qttPrEkRukrmCTx65C9A0CNttsNnL6XwcjUCZxMG7L01iN6nKyNyzu9Cm2H
kvjeMcu84u01AD41rMuTsqiZiRGFj9bf6HrKeWXp0FXDxJnqGmjjAFAWkVcCVZcYaw6SWHYdDtmN
MITbYkk1bjkdBgWMt+YilIvppvu3oZHu0kjpIKDv57gJvz2ZvFxfO+leyV0rA99E5ttSRtKrMZ/C
oamTDus3NYW5h7ZfV23DC4mmtuqLr9TN+6EBhbhUt1p1nyvZGEfpjJlln3Y1iUXyjSwNX6ZPzyz6
p6sEd3XwA8W9dORzbmOe8bxTZ8BmVTBeELef+P/sECp9uma+6EqL+zudskd02ltorZngC0lhwmmB
6ET3t9WzclBIe1gMDxLN2sQZ8ouz5a+nnwvhZa2I9Y8Zl5TVVkC7ZpuGUtBgX6bw/umn4lU4rLSa
Z5FTBymTYrIDaonWy19eaq79iew2s8uY2Np4CPoh7oMI86baHn7hPY4nHZiuYaZQQmYGnJ012wI3
WjtQHMvGlabJ0Vx7CGkDmI3uNk5h540CzJBRkvXdD3JiifqPKBs/xmQwb5tBOseSe58U9gWVC2Wa
+VYfgPnxqF7UqnnZjTamhAC06FN+6eOvvy9u948w7SjXYfcI6WT3o6W7/xdp2LxEZgX0EI384+dT
ou1vNqkZ4zn7eFCtONdvvLLunVIl71xbyzvQCu5odL1UCL0O8AucGfvi9fTcyfSjGLkTzcvp/HKr
2H26hdystqBWqU3VMBinkTNmuoKzxwocus/8mZX7KAb5za/Tp9PJmWZfqOdgEKblwSdl1iqJpv+s
Jdy+FdOpabbD8VCuT7f1CBTeA51dV/+4x7BWwA4H4ex+Ri+x629UdyKCX+DCvrQl5b7JuqCD7fqH
zBS+0v8tkt8ludmtdoZU1UNwv816HFThqJ9vn8MyQ5+VqRfZCs9FXVjGkspgeivJD9yhvYN+NT5w
0nqoVI51ZK8JK/z8T36/nR1Lv+bZw64hZ9APRmwEg+XQkO8t+jB+D6APNCQ2grbOIYibML34gGm7
AENGhhfYG3bX7g9ZSOaEaAK9dswsl+/+0kWImFM7GzSsi712wvebpxHMhBzhIyS7oC2R1LNrzQav
l8APzumDnmcbLKJl+Jt+Z7nqfGWL2sIWVjZIYrguGKjlC1B50sIrW4Wwkn9Zud+a5I+UjKJeDNvZ
KJ68boxG58d9zJe7Iww38KhOubW+MscHCMplT2FS2i/gWrjzB2FDFqs6g2a17A/ZkBeAoHP+2ptq
/zqBYgpO8SFh7SK0ZekbT1d4uVDqbMLxYXCJ42+jKAD5ntISeKcZXAdUl9UL9DffZ1InhT3HTXDe
ZBEWFT+q+iCrdg54zrbewJP1ij0FkCDfqastwjAbhnvlLziAe5D4ja0ozjzLAZlsAsLGyIokjp+p
ns51LWPt4dQh90nPaaJLuj/2upwehKmd5bPkTdyfxvnIFpQmYwqARnNZf/xzeyu0RwpI6XhVjilV
hdAyIBE/Oz84BHrUGb0Nnd8cEgwRBHC05k4HWbzg1ZFTwlUUZrF44EBNsLsOnXksgilrIm8lhnb3
AYxAF6d3FzddHfP0T1/WTT2nJOAQ5jzSm3QkQ1Z/+mCV2GMEpcK3XAAJ6bdAkBNn9Y93ZwZkXxc6
MWrQ81jimnb/sPl6vgXK0wpX8m7GrVEZQV1OsBuqwgLskltaLbIVYY/5rJr9Vs1MGg7//sq3SRUz
obaWZ2S8ObKB/hMRBU8xzyNj3dabqA7BH1bUcRLXxguhRh6JFaf+9W+YDLD3XnFGNk4wppN0p2Wt
JZxVbikocTndIHaSQmu3miHWDtYzaeOvt5Lm+VifKf6qXWoh5pNOwJ55X5SXNYMp01VoZfp/agd6
as9TUJxdEeAk73O0P+dxKJYB9GYz+zleVb272zN5U4db6mBV+b8uF+nGD2xB6T7UOrNtkPmOalky
hhl8jHhTvOl7T1WaAwNO5+ZmwxZ4fInBZsEsLTYLWo3GQiK7xnIXCXlV8pufTmGd0NV8+Mhk5Mq6
UccpJfLIieEIKH2v4uv9d7YlIesoWjqRIc4ij1EVd5Q3cs+HjKUKYR2ZA5Ir2CftUqn+5Z68W6u0
G866wGipviiHF6DIWizPXlW+/2kERhhZzLuKIBgcKe/p1VEsU0kQvzOmTQfHG5mXx2UsF6TSMrtC
Hh+bD3L2Q61rlVZbDuWR035VElgWRU3fqK47aN4+w9A9XP2wj64EmE2fE1mJrLhYfcMn/GGVA41g
IZPNstztzKxxDsK+onaGcDzBSUmVEfuqr7ieQfmMHeiiVDd0ncdCkXVAlMw2pZhkT+CAg0xPXBRJ
swpolMUpdz9QihbBog3X5navWdWUVMxRWwKlaPqZc3AGzo8LdvkfZic9tFiaSrHSVJEfvtIG7uar
kpV5HiiXfMkG9TTanrEUmmZaRmE/+/zYXvQRa2SG9X69WeAzXB4CaV61LJfTXN6p4olwAkdiCcHS
OHXJwt7xPPWl1vuwQUNX9ZtEC6wTEygGFyyvWTigqrkfkzeLZMfu1NCDQedyo8pwSSFTVYbrF7rv
URuv+gMpjcEkGW9WxEcKubdAaaO61r3utOfFU8M1ItW+o/s3tigdjEbAOQpmcdBC+FHpwKnv2/Q5
zorshxDAuse31XmUx+2UdRy8+sNBkODS9y1xH5kmf0oDDfi/4SeXGpPbo+ehhXB09zVK7V2vNDRL
BpbC5QrTHbW9W7E5jsBb5FNwTQM0ucECWY1iQFA2XNnUoGs7BMyNh7JqecWe525vxxdGM1JBjy9A
/M8ltXK1AbIVMQyO4wf+pOWix7LLQ1ADNTPtJdADAzpBcCHwo9YYT28kWTcCZEWRCc43RlvJG8cT
CIUhGWOxmqyfsPQzH/Dpd1laeUnyGyKuOLv6a4HZbVmt1qem5uEagi0gVuZ9VQIU32UcWzLLcndy
nxn1SYMCVfEDZRm+RmwXFQTbBzqVTCy81CdbAxHNLifkCmi70mtS7AkE60Oh4SBRFtvxbhILR9pG
UzQBh96v8YfLewHT2heuCYjGTfud7uhnAJCMvgjNfk6E1BmgL+DiBtHbgmClMEi71CVdLyYHJGl9
IF9Zhw+7a9Udr2Tj+MU9j06bX9Tgfq8tpdX7M3pUSU8WnWkT8N7Z321P2hB03fFoIyui0nJhiqWr
DulwI729YziHodpAWgVrQUPqU6gecBpU0y1ZeMHv3QxXnaio+U6//svMgQIrTRHUjjaKH/hD3Zsd
kH/y4Y5aGJF6S/+v1wJ1TuTg5Z6n5yY1XFy0i73NJTTOqoEASsd2/FfwK2/ilip/K81fP08JQhhT
e9ipbbP2p9FaTwbFYAOpTp9grlzGOIrNqm2tfl/Z3eclTQbNt1hAIANELdXV442T3/CuT0o3sQ+h
LdFNjucEOKO0xevA+3qL38kB0knVi5yw6T9cBIi+ZewF70/bmE3/mjJXMWahde0jIGn325GWneWF
rxwePPmBoco6xLWLOxsP7dzEF1oHorWYdjiImi3CiH7NMLp29mylDwWFUxx8lZ+WPZd0d0el+/0y
f+9QMkw1DvHA58OMkB1iVh9S+A3p14dxYVdiHoVaPIWrt2T7lhwahrccZZ0uJZL+coVetMOhybJA
dayfaTlfyvwr8UVPM1vBZxfkdRtxEgge0ZFBbUkzCH5dNFoB8NKyKcyPNA2j9Ca6UNTQVOlpHxrH
RNTq3Tnl/2glSKiZz3YwTVMoJIk0No+R5NiPz6DOZDOFKJ7jLZDxJhH5AdsOOYe3Q7UMwY8syY3M
tTl9yYha5sWM1m3fWWhvFjMezqjbkcqHNqKjfhdYTYVeR/E/ZsyJXPNJ8xM5P3UhA/gNsAxHZY25
9wHolFBN3aVPv5LfAyQLMVVFa95OS/QOnrfGKB8ayJchLQNGGYprs7ttgArIBWgRycwO9cMF9i5w
WD4QmTFZJvMwtv0i/51tBz+Q+34fYIFhEnt8cDo2Y7f/gLeWU53MDnQ991302YzvvpzQHOvxWPOu
d4x0Ey0GDJwG0J+Vqx3Ic7Okc7YFn9RVwhCS2E29z228m7EQ/9mFyDa/nJ40oZjaNJ0atM1gKC9n
gZRuuuS3v8SP9kGXl7Ol19B3Qfe4fqoTpcCb/c951+HwnpuwLZWtYwCYhwDJIg50xSjeHcxORXt3
u45OGWBEanE3+XJ4jaqYTESAi1UV+LzVtvB7kEmh8MaLO9MLpd2GVDiLRbX2SmZLlLwm/5EaNTRc
Pq7zq2OQsfUHOaSRiLr9wXr7xdBMEz1UNiBq1pNf92eNnToazuilZ9LWkoMLSX0N2KRygGpkx1no
2Hi4dvGP1zbwvqL04ZpRYdO9GG0U7G3aYj3nQcat4aFQf6fbMqa7+q0zZX6Np2JUNtP3IU5/4+Eg
oM/ulI3p2Jxuv/0hWKMH/2mVCn1uajY79Bcao50zGi2CAAbe0tVAklVUy/Bt1DS6hlkfNno+j7I0
ElhfyKo0VKLDLHzFos+rFSCmY2TYfRBBOoRapP7yRe+1WhGKsXpV6jUZhyFDGQBmoAtfWJAySLr9
0SacBS5ejWRTwPDdtRbYOLoHYb0UEjR96TR+4EDOzz9FBJf8kETrR0/RvhRAoRhAcMt8+W5zg5AT
AMis+gtft3M2JRgorElmPGFE5tO5Hk6oDK9/ux5Cq3HTJgMDfpXW+XM8Q6uYFognkhCfW2J9kd37
toP+paCuzXhTlRZNbgaMnS/d1z3DIk2T0xHmSpC0PpxIg6gHU0pvV37Dy7oqVupIOEyQJis2wxRw
YPx1dEMlsGEkPUu5G9QRewcVDs3eJpSykHTlGQ7vopy3V/HRawD9XaD0dj2t89BLZAGob6m4sRlm
Vh+RZ20vswvOskBuk5zacSIWy0eLoePVOjnbnKkrijK281AcIzWQNGmMi2bO3tWUxPX8WDObPUX4
iAoF9pXm4PaXiT9wDiMBnvyciXyO2z0NHr79lOBJ7yU3lDNfW10SuaBjfrmg+237GynEaeFSVg0o
4b6Kq+Mbxyg24yh6xDxi0ZJwcQOxtuVZZL0ySZpM7At2jKsVevPyIg8Zbhck61Zvb34rjpQBcD8k
HEXQ6ElFuZS7HgRc9jhT1uwDO4fraQktUn2zgKH/JuDKynB37SBz76aB0wgrJngPas25xqApPsf0
CCiKQH+oemGUlZVXQUbhSXnVxH0zBy0v/h8XtHvYn5ngERmXstZqYQjsgqoqUO3vFLjQOt+tb+WS
kuYfyNlad+RNCrvIjYrMiQSQt9UagS92txsFxM8O3UvCFxAxcqAfT18H/hdW8AoabWJYORs9TGry
I/l8DhrnhQo15AWZGhCboyXm06hqz1Thltr9GyU57DuI5FPn+SRRgdXyx/OGdzr9g8/xqaHns0CT
YV5B1oO/txkbs7NLDnrSRwjZxTaRUbKMwwr1kDe3/hUt55fvE92XOko58pWhP8PgHn5yGa1Dn/GN
5OignBYmHa7DSUMcWXL04mXnF9foqNief60E3RMc/v9Af+mwJJjR5riTJCEgK4CWr4FQ7xi/EWUh
SEjO3JCV/XyHlZ67h1expYC5QvUVlYpZAx6UfgPJ9tlFEFjEQDihhShp8KUgk10F2DqIUCiJH1gl
xLxNCtOrNJtpev5phOeeEE40YtAh9N8GX6Zj3d8t9wfKM1JwnOzyGoybCzt41RFfXTNo4Sk6RRt4
/rIIIm0iPBZyopRZCiA6FHcwMAldlEdBNaqlhhd50vF/kWnFyJWJ/2PJsm1rQ7L2U3WBUStheIIT
BmvzQyJCDxDS7RmxTzVrKD1+J5BA+wrnyLWRsz0arHgJaq+hw3GlW6HXNgxCslqM704OBiFJPQFC
9aFM7d0BcFC2HxvmC1DFXPBA7sum+0yrWuQW9AVwW4cfIG5M6rmmIQKpaR+NXWNcZF2agyIWDxoK
15tDk7FSQLTqihbZpQpi1Us8bhXQ8Y3D7mRnPZvsd2Jlu7MnOdqTt0mATLI/yqSa0EwSvBn3ODBZ
RarTDRHTE472TT8NbYEDqViIA7QDm9VTgXj9Xiayu1dd5tUbzJUNDrk2jEO59rYhSS/lP4X+QBP4
4nOH3T+cFPShhDtdsippJZSJnAoTAJhtFV28DhglvCpaeNerMypSxunxf4fEqpJqjEy+PgZ/ZPPi
rDWWCmFJFRIau8ZTxkceAtGdy5RzsacdEMoGfhPsL4oDWgKpPQkWsR4V2g//OxbU6AHJJUREYKt0
jAqYyC2zLO2bZz07IMSDMtXtfCuD09mpQX8/FksQMUzvgtEvUiyK9EGVjlSSasjnNjqfrVHKTFLy
L9QU/YEZaBmqLJYeXIL9JmiRNVVLl9kJyLuaDHAlVcn7VDX4My08jKsPbL0bQEUrSYvGIyxW2IsQ
25b68//PsfcDyLdk2GK9dF1LoQW/qG8Zo6VXIfsnJV4TG9vGuKvZEB7wjwsqWINh5dfOT3G86d6L
+3LvEKqZ22I8ZJdfGjXsQD4+PkH3pLtKrfWncooHxDwoxpHRC5G51KoxC+pdu1mOIsB1wRUg9FYz
WKdzEckvvb+uWLNC3cOY3bfhpdmDdYyfATb6rOKA3aChf6RX6MtMARDTvhCwIZ4bGAD4CWI9riTg
0ttPnvwSAjvyO5+/NR+3J+chljR5NlEueAFuvV+K10pFjvRAl6N0PlvgSHBlMsS2862b8TeFhfj8
fPribh0P9tFct8P72U3xV9zI/fQLWyPCex5lIcQ5M8K/MYT2Rw3GMtR09xsjIoDtT+kPbagp8cD+
jvPjFPHS3WHlrC9kL+n8TJTcqoJOLU2pzBs9Pm4+OFLIQwOz75//Bw7EiCkLE99gFsIIpuQQ+yD5
vNRIXpoUgbSvFlq5pF97dQ6mgi5eCmOQWl/c6yX9NyS15pvvXrD671OP71n02k64Yvwav4EfBwHi
yHG0JDeKb81Su7IMj1UCD2doshXgUDMW0c1//T6UTMlfZhK41tO6Ewalpiz9qrhmppoVJJEoN3rJ
EHAtwXnBpVn0NfFO4ivmcP9HLmUbnAdBxL4wwFxu+sNC+t3BDAksbG8wsNn9KHMenOqN9HrSXFhf
+jFUscaWusmXQujxoCj2jCse6i6HYbkZyU+VzWzuiIBg8Kn+eeF6Ccf71bzVukEVVtsDesyg+Srr
qMP1oAHa3VUqZOTy4AHuy1iyUo60eZsb7CgltBDr0eKA/XkbaTy/Pd/F/Mi2ZulxiiY2GEs2EG46
jGu406FlQ0MHvUiiHYuFi5bldwq3+1ImkOZsfek3pQXSsvoOVUnYSQD59aatTyhmqYXi3Q7+8K5c
vkFOSXa9ILFEhlODgjyi0tGwUAmv9+j0WMJab4R/7MLTWczu7tZ/036CPy5zRgxXE2iijWjjCsc9
KNedK1Cif5+b5d76JXstNAztsECs46lCDXAsuawLtx1QB6SFFifpi65geZSWKWNXyiIMkZDBNWti
nVGo4vZI0tltgFZrQc2ol0QOiBTCRKh6LXsXh6Uq6TZFkx81sgrVnip2UYOLZAlHqePJYPzXHsjB
aEeF7HeC7/lKrZK35tlLNZQioiHQ3wNkyaZm22aqnAJIOsLCvLc2sOariVorQtTGrhcfHnV+VfBP
xPX+1LMekMAEuIodIbTfWEd9tJ7ONP+0SzI6gW/2Xp7ox+wXVaMSyu2qH+Pf/Nu1heJ5XyOm7/CR
wgF9/uiBZdBzwTlTJsHxdTCi9HCX+NWGZu3Ndto9OIJFRAK0/BSsIaV+k0GFirkzEgEn5TVLFwyX
X1L3UikfN4Sl3uBq6z2OWClllJx8N+nDaSa+4lWkqV9qvBwYtbGonnU/1PS+PaWQNkTtGhDv9h9R
VhycRNWsDn95pWURaPKUtXxM8VfcEJeJDDmEqOPniZ4xj2sZP6qtkmbCnJHtAURd1eWyv8kPvRCH
RsPCcGNzchkbbYlnaWQ7GLlRLWfD3LSrWClkRc3KaLX/VYC8JOfSGJkccH8RfmdIjNGZWPPAkkyS
7ztQsCwZHeQlFSLIgWWGObXJPPLi7fNcxUBlpn0a0jXPyB8ti3J3dMvj0CUOVQNz6T93Jqm6N4pZ
xWTGxPXaxrWVmffj0hDhnXwsdO+5Sbdl1vjnVEfCJM/e4K+CFjLHNzG4kkb6jKnKiZc7KmMRhsQD
rRIlzRG8ZX2pucJkzTN73rE9HmSpSRxmNVT5HfZILG2PH7BzcpxQt5tjeNf4ukdbjaNsIqSnsr3/
M+Ex3/3jHUEg0AansEntHdLkeApI7+9zXrbXoJ73uQFjXkpG8yehJHQ0a2D83lq2aWdp8UG97GC0
Wks21wmEBLIUpnOqXL4Mb5kte0t0cMabwtuhOwEljvWJHHYv0+bc6kAJYugnInhfh4qHUKvH5Lct
0xlAMTtYLEf5KYDtomecPw4wvoTz/WGzSRHcp+p3azOjPK6l5B1kGzoGEkq/UsDkTCfYHGttIpn9
TPqU5SO4Xgq612IhU1xSTIL10O1Th5R5VziafAL+o5z+BjVTcu+C5kQJHTezPUfHrvnROjXvQXHk
ifXYuxfZ9k5oYmoDBBCYib7BL9UqSDZvyQstA72lF28nNek2NnB45SfUB1+dCatUoEqNf4/lIKtm
dLHOSvA2g4bl3VnwkoCUOqKeb01isbC5RnBJmFteSND67TiLNFPfTIxw1Y2dq4gTkpv5+H5kzlIU
9AYzj8V+bDmHZz3VLjLyl2THoufL07iVT8gLaJeKRyeXy24hfOUl9LosZtxtPBqDIQv/nIlMKqv/
okdkiitO+0osoPPApJntWgUmEIQxovETJNOfY0Jgfop726CJhaWVQ00GjPz6E51OtGqZ0P/sFd5f
ZXCyJLIosnWW6QD0asbxYAFURqvw1gBa8aGKTyJlU5jTYA9/ykJrjdOMGOAuukvg+V0IJE8Be8Ky
k+ID81xE5oPzh27YEAbpnpuC46VdI4OelLtN18jR31MYUgipH+ELwBk0uuZq7f4JOjAmZTUm7WOA
FUtiTFodT6i5sQ42uG/Z/UJgou9SEffM+AEt146qorBMgGLTxJpbipvX9L3qVE8eFg+mO9IrSYXo
C1woKpviIdH0cLDbkH+UcoaltbpIbF92jPQjNvkpb1o4ZO5YyOTZnka+dSmEqMdO6aKRUK+Cfmo+
vvC5ghFNYeTRm1e7UsZa2k7HVKyrLUq1zsAw12YLCpHQXscHT5gUd9ohxS4n1PBCew73oXCE3H4d
k7Gwk0bdIap7X3BDF+/V1cvWse7V2x2JQK8Whb9IVTk8+T+XN9tI+I01DSSWKfWy1kzXFrfzuOFi
iyGH+RjYkbALMgSzbGj8G3R2dGpxfTPBDeDA8WEWN4wxU1M6DuwT3ZixgKmfgJHQ8o23SqzU6g8W
DM3Dy3L1cngQw57nIaSAC01HJs87z2S4ScMQorjAE5ZLa0SF5rLL4mvbSzilb8A4LziNDJnh49Hh
jbS8ilqcZKoaGfU/vpzgomZvSnhh876G8P92Gp1Hc/A/p8sgFBOfvC5WWe4QK3EAnWMdquaZRGUz
VvzRusVqlYiz5r1obKxrt2KMsQxJ9jcODEHk7/kWDC5Xfqnb0Fl9ZQoyXrrQ7naXrxPdLa5CLtvD
TgSje+DkvNwYtT6ElCEZJT9CLJH2SBMXZL58XIa0gwzIExGGzWQNwfi8cIg60ZuEia7Bs5xOfe6Z
ByGZgf6Kga1OAC/V5lJ3BcWDhjpz0KrRADKzMwF9wH+c3JQ/dvDJc7QWwV4bMXXXT6Eq2L5Wa5ig
DfmM3oIstZtJQgce54kvfmawhYicWDmd+VFXguuRBp7pA0htru/8Mss9lCkEM7rOLwqgH/TB7oEi
qjyGQSiqGtXpcFNqpfewjI8fePeDtTN0d8GQ/4791/etu+pZwXRC9UGCnQW7DeXu3XHerjVYcgye
MB/MXmhIuHuq42HkjKZINESz9PEnzqjg9AgAAwgg8ZOVak1vE/MirhGokdAaiBuqxQt51pgis6OD
OrdYTMGa/30YLT/aojivxgu/IU8OUd1Ah71hBV5DVVDi2Ala2CgFeTaGHA9QIYWQJ+xdUJIqJ6zX
dyhwB0dOQ57dhlZxNfhYzTsxionDYPXSXg7ls9BNfl+z66WBV0AJCJRyHKYRJgrrJY/mAOp7y5HP
CS9efkioqW4vw06PVqaeY+ANBoLVq6O01EPqDqk0qSML8T/pWrKMJBcIWTIoKjFvFTKeSR4Uc3bA
y/86VbEtLAxImsmm8KWuMxPm/iOaWw6C9nPrnsQH4LpuiCSD61Z+FtoEacz2HhmnG62zbJOjQlfZ
NLTyirfBPemuXLWHPewxIQwaxESOSfTHAHHyXH3vnZwLumW57Ve2vuYG+0PDfNUZgtt3VuLw5ZLR
zK4klFxHd0FqM1PIdVQbAR9yLH2XCdoxQfUDOo86qYD9jYbQsEIu38oqp0h778WZ7+okqa5BuVL2
nHFDVaaTMi/UmCLDKzboRM/LJtk0RbkUpOEBrH0InXD1zrngtcyhaGTHZt9fLQ0wBBEEP8R/IivF
lm3uibxlYXO9bjYwbsfTp9aLBcAIjhVGRnf7XSvQchBW3t+h0vT6tyB4o5RpefeT/qrB3keaiE4+
mWbuJo/iKz4yukmR+KdYxFDtc45sq0zGHY00VuqAOidLbum/sbTrstrHIVYk/o1tNrFBEOBYEske
luirMsUf0GQtG+iUr6Sh8d8k0mOaktINSkwcbyaQaEK6n74dc7yKpwUfCUvRPDN4w0GWQN6HSt+2
KMITQzJg4SQaweetf3lIwaeayMH1R6+O2WYn1RL/8hh8ygK5xAluwH2ctWNpQDqYgO3xo5HH/dT1
/fs5Qamy2hB8pirdRI+VoMetbplkq9UGDswzNeshiqFgRht9tWsvhlnFihb9evBuFF626KSI1ot2
fo+6XTXWAV2woMTsdaVZnD27DZiOKhroOdZxqZSiRXXcqR5Z/Zbk+0T5u1iivoh0N1e5k61f+697
afvFgiFvwBMwnC0HzF4qmkVIPIYVVz/7gSQkUFE6PpPxHG37tPIoPY/tte/mjaqvXWC+k5q659CQ
/kvHkQvlJktMHMAsbufoVVWNqmXghuEV4SkzNHaxoKOAdBE6LicMCU2+KoWE/ZXap/vNK1MHFg30
qpGjQuP9PTulpUtNagfDbZyD1VbNW3THqxO54oBR4PF1vuL/Xml8CAUtxqPp96Me8g8fZn2aO2VV
1cgtc1KDyMvSrv/mfok+msBWUgkpavoouEKKXWB9eyqCzbySaGFsVo4pkpRvyQJg0Iq+0pjBsNr5
wjp93eLKihGF+7Yyyxt1nnLBloxqHlFjF7LOwW2wk3o3pEbcuotYiIDMTVRwcOPh0XyxA3iDIBAI
3zTj/Bioyk3z8SCpH8WmfeYQ2iPrNckhel1BjdhwQwASKp8OstWDW3QvG3b0118L2u4Q2YPFvgk0
UpyttwzQAmHbVqUWVMhOIQIIdCkrPdDLWiQsbucmpm8nu55OyYjyQADVbPbh7wPKUCkcj3V/FrBh
ZkThVWwSRTGOXyy0cQugkec3vVnf/j8iTAVN2aXHlw6eAEEM/AJMbuF9V4lI2M5itDwMjX5ukEWb
xPfg8ws1pR+cLXZqkBAz6tH3rqNKMk0wpFcyMU1xS7qPJz3XpfHH2zARfrIBzDIQHHkXldIzXS/o
ngRADjRZPHcKO9D9SHRoN1u7M8XSVxcU6Ta2+S/e2xuUzoVzlp4v9aWrVyAIg5mDdFQJPr63xp1m
5lBMme9lRDBZsOnsmhcB7QrSSWqL1aCN8CvczTPiRLa+JbK8E31Y9LV+ohyGeNyxS71dH0dum4o9
qfx6HxW9SomwOa3jKgzVCmyU1cBCqslX0zNiu8pPdZbnk6ut6+hHliO5wwDiB6xDY54UtYNliZ5n
0ZQa1WBggrxZpQe5FBo3iZxTh8RRA9hLx/W0natJFzb0cXfVJk6AxOQyUC/SnweTNf3lcBmU6yLC
cLV+wgbAsxtNOodoVwH1OycVk2B3Vy/ptd5nDDWvx9O/t9NGfKID0LXc/qlT3f2okKoVXqFdFH4a
kmx009zyzi9phD3MMY+T2N/F2HG4HN9+c0t9lioOu0wQHt0yty5LGBg0FtRNOklFjIY5o0znEdi7
ezwQskVfbDXwYdtNfOas2JCACCrqQ+S2knQYXGwf6+13fEzOdrycVYrD4Am0VREPnwAErNhXUwbT
sUY71I02Mi2P8WhOiEBe9pSB8BHAwecPusG91xftWfh+e0CI1vAnpEbm7U+wWnoohu48RT5H36ho
1c5+PBfO6mpU+4igac9nFFM61nhT2P6IboYUebmo3tPWxWMEFxnfiodjZrTUw7VR4sZHAgf9ir6q
6Yr1OK5lCWD7OuqWQnccOw0pGJejdgHlXW+/m1WCmlcX5imKl+YeiKtLz5qS7QjW2ksMLBao34kX
AnIigFhfqJY87jV6hmL4I9XNySnCYp3O+FuElH9IiDwFqgmNMhvKjAaqlSnkLowtRk2Ou8M3AF3c
oQt6aWc+wY1NGG69n6+7zFZpkEHgGITh3BLR0p/+q3BMe3XeFAg0+fIdT8qcPd6Vdjq//Zvezl5+
MUqqEPZOKjHtkbsXdZ35jiALSM+4brGfAIYYJNIbzzsF1Mwl7sRQxjw0wuG+Js9pUGKvIOFCd19h
TwOq6kcO1BCbeTih+Kf/FplWsO+sL1FxRhg4sufnujWB34K7mpg2Uf6nHzyRt137Awa681nPQfAq
1TlOUTYLH61NJtiPX9vNM6DaHAyZZgfcTYRDzyYQ57ouEMDu4uGJw2uROk+hNC9gb019rX6mkWp+
7Nb6ee3Qt5rUq7ZBiBDuKfaYeuIktOsOCKlK8Qh5h9ZsDkwEdGNybj4fWqa8vvMwJDgmWOhAbpzi
s3ZEk7BvyldKXtxhSpNANt/hNeW50xdpHnvTlnUqPaaCxpS6pRkzDb/djx0d9f3H94ez6B3Rmsua
eInIewxJrAhstnoAv7aeIm4U+H/lq/lw2V/HUYQW6vlKuryqjUtA6mb8vz+kttGMGnLedgdCfZ0m
Ezn1xS9ilnD4fNEbkcD7rDhqb3aW9oEJBtGnBZMKcJdE/ffp+PAWwNvCW3J+x/RMWlkaqPIXVAbq
jBx0HcYpCE3YliKuHb8+OKZKMHo7RHzP4XMr/0ZVloLGyJv9+XvdT07KfCrLq0LmIGtgj6JocYqJ
1/xTk2YT/9WRRWPHU75eL2NfLoRnzZT/uFTY8xEZ3UBlRMKAUN3lkz2CFGqo7+81qtt8LeJbWDZo
RxlcrxslkEB33UuEboCyJA0I/juJTI8x5ooB//4qHMUD7l52Z5kVY6njt8zorpDSBd/jAxUynezW
KJlp0m5TQ6EHLf3levIHdrXQPYdPAIpAeWtH2c5BLBnrb/Le1pS+Bjo9gieqArniNFxt+vH/b4Mw
dcXgjVurUasjtn2v1osNrr9tzeK5OKId19IutWfAIg74R+p16b7h/vW8oYsBBz8/L7OE1M6/jQLN
NGmb8X2lORETrxqxvzDyFsqIbJ+OuOv4JtKiAdYHXfEk/a5NFN2CoZpV1EYyP3/yVB6O8Jvj/Nxi
CGHbbFf2csZ3dMbtlSZfDZ65jBHTvVMHTeTCoLlnnKo4sIBcDg0eUhjFbBV9fhga4HWR2usKTF2a
A1d41/VHdFEXDiAfWRSxjblfjiabYQjxJpUp/ko5xovKLFe/0incQIW/FC0SLGptaSqL7r5TJbpa
iVTjAvfGZuohowoCcQNnyQmpM0Q7s/BLJhGw58Yy/zbhgMqnVFuVGSue0kYWWOUF3KObkKMtH7vK
MDPQ//6GWbyV2DtlhF9c8AmmCChKCesvdEzZJrC63bkRU24lHprF53kzcCe2M/DEtGA9pfhzMJ8w
QwgYg5H3jiVblduXCRgzYxZTIYoKpN+5kJWMRKX43WZwQ5pUZRgtiipthYjLLRl1X4yFWBAZWsOC
VV3q2sPm0QyrgNBSyrGqmS8eWtca/UJbkMRXeLc+zFhsm7EelnjRceJPYwXH0ynIRpuHbR1dV/nF
rbFqgBrr45gsjk82xzB4yFUq+YCiaj5rcQ9m+D6gn4SBoJX5iit0DfYLyDLWqliLhlptXbW9KXMa
nfA/ztYdit7oDsMVgnxEiFhhlGZUVEBa4bvJfcdrIbuYu0147j9A/h6rLLO+ZqCBF5IsZiXSw+l1
kf1tT3ZRk/v8rX2QAxWhEaxkAfyp5lEAZ/ApGLoovWgRcDuc4O8zUzsZh4QJmv/l9OUslS+8AJ8A
lqN0LdIZq2IgU2oRLeNgKMnCxBn/wbdoKmBhdhPAi2vO5oCTenpnPTxstKkaPlR3xgN+3305TipJ
TEhQI6Q9lt2MuO17yD0SLvP9lfVZ2qqOMuOvR/tPWq0SgsaJMp1M8HjqrB/soLftcW7hrrHztmZT
PL8wAvUTx8g95kKa/T3e0q0zpbS/cTwr84FUjcM+ZEDqOshdR1WN73hfvSEr0XuYCIs72ISuRsXI
vG6kRJP2FpYc+Hr5bXdpXxNHoJlwK93+jVVmgGtkPn5xwRpICgHtSAUSgsyC5rWPvJKunCEYe+r4
eG36YGhCsMrPKZXSml3kjk0TSUFx6eywxIoR3QjEWm6Kq8xnQEgu1PbEQMWfujRoOwWNwdYHlIDx
q7tvLrXqIUzyFiYg3xveJsPfH6yo8HyGU5IauqNmc8dHf8HYu1BZBBGfz1gK0PizF2o+P0SBr6xb
+TH9Bcz0zWfy9AfaN5fzUps/mG5bc1KOhg5XI/00MVKX7bCuPnExswj2gdSku4LoelhoQuZA5DP6
8pt8AFIdple7Pavjyyi/SsxRV0A3KkUNKWgRdhPrq8H8Iyhfi0wMkaLI6jzfRNjUnzi4p8fvE/tm
LSyp5cT+6q7N9b/qwMGe9FbLiONGeL8ZZ84UGZrICe8l79rtITZZQFjVfYIXk32Uh0YqfB8OCGrB
uhGyvX647pFPrgIn06A7uargMCQtmH3BUKnDCTb+XXqvJMTQGVIWISQwsP61bN2lGE8bM1MdaQik
3tL9AAuLLI/xBIFgRQ3U519zPoDNK8KEAFUDURL8ku0uj/8+ThHz9wBs1fNxqPtU8pHFGCx2IWxt
Ragzh2e/GFNNZnANce4JbdooMBV/E/Iqf2ovxw260auIZ7v3bOBHDlvATpGNqdjq0YDWGNBuMcVL
Dv3ZEH3R0AsYQ+b2IjQEBORCfVobO2MnU4K6Su0N1nh+LRzjiZnxAQGVEzZC9bahLt0YOXt02iYT
uvG/KXCB8seOYWQxTqlsef5Xaudty4dsVnlAExWSzy1Njdn8+cGvN9HX9oilXYQ+GbjgmbeCHc4u
/o9xrXy8FJO8xZt0rEJavV+OS6uCrW/npvgL8S+W1O5Vz0pAFliuiG9liL1r6ZOfrSf30X/ef9K2
8+AyVWk9kyEKfwveauB59fr2rxV58PmJGJOmUGIC3CPdrUbPTXa14R2JduLiaRT+6Y1NUhan6rLu
ti6plPBrHPwYdVKVbmk6sE91nBsNa23gjhIK8OvTZlvHv4x7vEBQDURtsScJsGtps41lIJd7lldS
G6i3G8ObXTE0M5JyLgZlEwthY2xyQ+UfXpkhtu8JFBgodu0AGHV1ez82Lm8s8vNSwMSQxOTB1nrF
SX0Ni9wRCTVs1dwvsQs7TvzMHoMgLL2ulhEFn0McibXUa40oZkQcHlad7uhpdpWzvpd1zuXQTMYH
h6mkGyHEKnbpd5J+N/FRV2cPw+LtMECgKEzKItrZOq+kQfhJiowZJmUuM8QT1Vopsx5hm4H6BhC8
o9T/NtoD+HjTomnX9ASNjjOfOluqrsE9Oun5EAgOrsLN9giRGY38Wc1gjNojlo7yOmRRC/N7rzZ0
8hQ7d+3PlfMTx4+MmMhnYjtWqCtaJPUedw2NdrcHBQiC5EESVM6ayPwVyYpZkVlBZcxT7Vxu4nZG
I1Motlp62m1/STfjNGzkoe+0C3ez0rTz1Slo8Xg1JOzHskA/7s2kjJXhsSrYPP4Nd83mHxQRLo49
351L0vxrByOLsUKdzb7PPiPuXdPyExe9XbANK4jyKek33TsHndkAr5vCL5uNCtIkEbvDGVEsMPSr
IVmUsg6ZtxaMDGxH6nTeZIWdbfbE/k6hH8xf5zz1XNgtszlip7YNpcYmf/i2sWD0WNYkLcHdewbs
6VsjPFcppbw+Q4vQVgvG7pVMlTs3fbCehCO7/7cYRlE5WtV41S42lXpXaAFoFmOlGEneL4NIUKX7
BWQN+dWtWQmWisRXacr+gEqdzBl83xQrPTMJ9/KIh/Tw5AovoqDI7mfgc6wUOQ76CtViyYDuaySR
GMsAnmE3wlT6CsyEqyZGGXQ6Np8egT0Grcoy79GMrLRUwnc3jF2uQFT4NezjyeCU+U9nw32DTBbi
S75+LP6ZD3+jLaCWrJ/+kR4ab4qhsknrcFKeSFaiF5g2ay4ds461BmmhBxO/0HyChmIcEZnLWXOd
EtpSRwMYfJs3D9AKYQsDQ/t4+la02u4eNBGI6iMVzQbCJ15eeNSuy/GRNMKywnK+vTtCiXc7emjs
nsDKtFp/O06VYLHSnXOQ4HCBVnz1bUNTJDAIYK92pK59Ue1nuemVJXHmhouGUXHekZbMBEhAkvFv
u2SSSq66Pv2LgVuMw0TvUKY1aG11+c4dASMvN8EbzU9GpmWu8AD0JFMTJdQVzBYmUFrm1v7zA1/x
9F2ZllT3WLqEXgMYgAMXygIiLUGiUbAEZstAuEI8/v0TLkXQ1irNm+46OOUefypaN4BKro+7RWCd
QBUJ3uu9nDzh2eSLtYplaG8U4tm3PjHgtLTXnJ0Atb7JDg/rilnQKacRWyA7L2gPgoul3SYN2EjR
wPhFxKR0o4+cb7fq6CXzYwY+baBy0Ytch7UVR3/FMGLpRw+JO77z6VmBOYX24GOzpItXlo/iTk5a
Ni6OnCowcJtOubwL1be7ho5kwm+qNgkRlCEwk4PPez4F/+VIzdCwWVjl6lCWofHNn6NUyyZvas95
X7Nb/bKezHsYHCb/HWRXITpjnm4IPF1W2kVyPDhbJ3o7r+bvIG8sMdjiX4oyRWQcdTLWCxG4lgCm
mbfAdGOeN/DxdjqjI5ofvbiS6SSF98AHI6ju2L02xoqgCLEajAdDuLOph96of8Wd4y3xwDJjpJwr
Mybh0D7SMflp2Lz3jLwnbydlbnkPh3lD4GcY4Qe8RMeUM16q4IIjBvmE5I8jCJ7kF34iusCZdM5Y
52rJsK6rAqO1nX0RXm24igx4L4Y9xv2RxLzNHV8luInBGwXSocvavfteR6yBmv+cjSULE642rBBk
ixpysO8Et4ZfZj2tHVleojjJmSmtKLzBg5QVEPuHn0TP0RR8CYmH7pyhqQJfWuEDtmEN9ABckpIV
Gq0aWwlAfvAzyqhVLP7YtsHcPWhZVcMBIlrVf5M2LaRL/SvpQ2NFittmDH4la0SHCcuMOPMfXQxY
QoTur9HECEniiVpQbXWiR8ZmHxp86LuAqMUdhcTaPncV1OXB3S73yFpUQ5vp264KYZIsiarAPCz7
1kOyLHNz7mOgekB3WR6Tk0xZ16vKm+52y+8FT8sYk1//SvHxzylPl2mLz3A6yy+Kis0tFi0fRqhx
ns/Nn5r0t1403PqpNllq305X4qjCUVwC/0tA8QWgqUfcD4kEn/B/DBu0E9+XWP+EGr41SPMr0EqB
RSspFxTfDbwINz5/05j3AMZ/kVU3Vk/wrSSOhPzx0FHbqlS17scP1EMCB/ZP8rAlIwkAexIDxzrL
1kfjJ4NF9Q4aYk4Kgvu9E5eyWbD25xzaeYjaIAySmTyZUVZirfnhCLNuVZPN+RmD7EvhYnou6jth
IKiw2zTrQy8S1vtZNVdTRMV0w2AahxCjfHbjgT3vaAJoJjkxNZIipD7inJ8WjQcFhEEX0TL0z1eE
QBLx++Hhy7s+2eZfGHB3bF2Z7iwtf7XL4mccD9k1ZaiGaI7F5TQon619476rWSVykV7LQW7UJ+Wk
+wS8QuxvzrKeXuaD6mhr8B48hIjdnx2DS0Vf+1EUwYfoQnlls9gj9V+KpHnzmTdji3EuVNEgOaAD
OsIN2UoQrKOj38r/lH/UOrdkS90EfMkailpMsTGMcq+gotcTA0+wqaruRR/HEZA/pYQUJLb/OviO
htA5Ni2MoelX0NQlJvtPjVU0sFUhtw1c93Sw9cuQn2pYCB6c4e4uv3RzK0WTtO/1xcE9xJ64nd6u
fZTUYQB5AUQ7QqkYyqWZMy9dLxiR80eEtsNUAy/VzMBSEDQO/DEjjFBbj8K4cebN6jKzF7UJbAh7
Kz/tXiGz2ymaKVN/CjQ8LbO4RnyGuQ2/GVxnghptN9qn2TH390Er8TdlUDC59JwWI6ni086zheKu
BRTk1lCMLkoZv8hQwk/l2im9y101H8MDYZdP2KYUlZs+1UJGXuFixInCKA4VtsLOUcyexJLifBp9
3vj9MqYQCyXbrNe/028zw8MYxgfix8VM9T5PVUHzIWEEvzjvUvn860kE11sLF6T140jPnBN8X6Sc
eKUX+CpH8+cSZn0PGHUChq8R+gnPtVdwjiLzrJZ0GzZRpXISODY7L8/+9NtofE5x+D4/Z6Meq0On
HC2KXYJ2UzMtQk/RBw2vfbR13uZNbrWhBTCXWZ5qMVJhr2TBZwJLrZVUjDCTUtqhw+0ELXbRSU7S
MG4AX30gKHgl9eymdL1udPGG9w1r7aOdl2+644/gvwK4uh2Ddizg14Q2eCqaoAXRWJ3y//WbOoOY
dyXItLheQTdG1mvB0IVhPbjWZmyEdnr12g2APR8YIZRFxnyzP4DPKsfaw83ZrqSVmIl2nDwZJy8m
+bPUgOoeJR0KpJZ9gvBhvmlyP/BsIkSQ4inPhR99ZkkE08IPvU435dzGg3HWPml4/mYa4aXGtPSi
3EvqNA9wB5QtxJ3G1owjLGL5Hht25k06yi3wKmWGGJsoM6aZNunHtSyMoaSiyV/QdYMZDJoqDCTH
lXpDkI3EZ3GzAwNuKrehJ/ygXASM8SjFAWg1vl/eAlfOTHq26L1qop9Q1Mr+6DRqg/650bXD+EzL
ZWkF42YKClzL3vi0bBPVUpJyspHY2Ol7NhIBGOI7tmQzWb51NVa6g682DWiwqIxLGB1SY9Hum+7R
maATHvvXrpJOKOSFDnlxj14xl7TgJnfpmBFt5/gUVkWNHypQXSrDSMzyy3KHRi2AunHjDyumiCpt
6UcoQU41JV7xY5cNn7lDhArCtUtidRE5sWdlI3K4rfhecIMwH4Miv6Po0JTkWc6XUYU87Swc13PC
1gf4lPEq7LnOfflcyvmjCxX/BCyXxbMU1YqjeSzt8nrSNltCqhoxAZxw4LF4Gve1RQ0TIaj2AT8+
4PGMELXbao6v7zrY4qlEPSiM7KbvmatK2X9z+G8utTlt91OikhOOCI/Xanf+yffP8Rwv7Tfi955P
12ALm24IbZuECngTqM1C1bx85Jv7X87eMBofW53nXruezR0l9LND9cboM1UORF4kYbpBVQwtXyGD
zC9FvBT2C8B79frK6e61DTr24PJZeH7AZqtaLFebzVBBK01L9pXD2TudyrvS/Q9EnNecJB7a+CZT
loKS5epxdhAAgaM/nLfByJ27extxVZPXL270TyKAwhglrcUr42Ho6Kmi3U0VDHoDqC+v/GdeMrpr
C6fbgPT20itInjw74XbVlngd3wbauOwR5NUp2h+EcolVebiTboQRIX+zO2QtnZex946FLT5E6TCr
my8Xi9+hO8Ps5bIj3fuREgjcJiVhEg3WLmxfNPivOhCvfJo6qpdaX9IzULpWve72nvt+OHEIIcxH
d6rgQP/BeIAlady87Nu1PuJ+mvTkGqfxPXnKTkH/5HsuC9wdegmTX4StfoW7q3pd/ATV1ZO3Jzl0
B7gf16ecs9Ow8mAlUAGnpImQQGx1cxPN+gV7Mti9UYAmPTDdLHDKr8amhLzrvrMi9YtJOd2A/SbU
J9m9yQofZZMJLmwbzELXq3HXMohTloZh3gJBfHWli+vcki/PhHlPj1smpOV/mVgdZxYRMWQulYmO
Vctyq24RCE5P9YCtmE/NqLPl50m5DX3XwJCysMf+/JR47kPXtIBYGAmsO27Oif7THrs5/zlEWHur
HrljVkVxf1CccIYQNNkqXlDE0ReCFOgJP4VWiLuV7RyvUPN97ulNQzu4rqP+EVFNFZzgoaAksQVq
PRvmGURuVhiAHJ7SHMuCxK6Q57E/gav8GeAumqn8Vle7KJwAtUY6vUJmZpr91qpP2vbeGJfh67q/
RKg3eLwCFm2dSXuxUCuNOYNWC3jlneRB0hQbDQ53riKX8Av8WsriY12p2TAQWRYDQuXBmHnNTwnB
z0qizxP5kBJw7LV9RD9uQgyH1oYErweaOkgtDn9tX3o6s1vfRD3vYy586ZoVQBksGxa6zWyqnWS/
TKhGufcN/hM2GzCeexKtWAQ9DG7ihkRAuqyEWbxSGNlfIBvduch6dIFhh06jfaCXoSJwZWb3pnO2
0dKhLtmqYmRqdCNfMVVZekHxWV9BlBNQ7rAJDK2XT7+iXgcKDdfVLx3U6f6NAz7Y8FKveZSM6Vmj
aPGyBNdft1WkI+hSrryPivnMwQxuzpFM/taSbBcCknI9ueM8mOC9QqeUPK8gkSJ1QpSvE7E7/2QJ
39nLXwJsuA814n8WlHf+9CCpsuGOTO0kytswVMrOMpnkHpTVVlcNEaTiTkPg3L9rd30yDHYsVved
W9B+sM2I0I8cVDxEg4Yywxl7aqiOIA1g2UCFiyFDj4jb0q7mc8cjiyrUbPdPqtX8toEe/gjt1XAP
mFE9MQpwWZd8elrKlC2gRkGUenBVQGUAId+UVquXow85r4RjKp4zwsFRitmS8yuwvukGS7FJQtwA
Zjc7qfJRNUdBVHzkbsq2rPA5cCiLaOr0zy1u4/6DW22xqDhfHRNuvMi1WVSNJLcxsIaUFKdLtdT0
hNhDFVvK45uO73EutERxEGVAdSwHC62jU0JPdTpYRfGWMjsaWg1rWtiDQUXOrwWIS8a7tKUQ+xga
tDBIXQDWqybXEjXTK+3amLP+R96YzjmiXAAM5xeqKObsNS32/7Ewj6OblfwJf1mdIrQGgWcf8GTS
kAnwFaDPyt86Gg/JSloR+wv3DOJY8pZYm5ks2vSrM8VKI9nasGq1gWZeK7Y4Lcp08GDlOZ51DcgK
tg5lMoPzze4DjYyLY8YiEXF3vmNVa8qhoj6LExvIJMyHiLJTRxZMv4SOayQh7Y3rt7FglnuaP89B
DRfuFTm7uWwTE032cTouPBs5tYbOvcZpD1AXU65ZZiZIWY3beSVZIc5Zk3T48lj+j5sFxTyzfRU7
wtkAwpBxUwWrZtmDFb3IAkYqlv/JUzCOhKlV1/R7zBTmSITcRLMHDt1rD7MRFPh5496ircacjdVr
MOIipv81pZI0errvRxNxWxsRV00nuqDFW/TyO0dsAZ5FsBcX1wKdhgnny6zr01TtuVvObBZhfGrz
AuInHRM0fcKOH8EuqAnD1BrG7Z+dcAuZTFY2A8PaJe28hj9nHz+7aeq4tE4bNbnu7l+lDN48uK6L
LZw6kaTUy1oYn6EoOMcD4+VfNahhB0EEB1COw0Vd+qpHH+bntNqcuaZG3HzBEgd51bb+R7tX2Zo9
9wae6rTzbccfaUtqHyG8WGetV1h5mbKllhgQxny84FVAgMtqhVlbHEgDl6SCdja8M++fZDFC+j2F
tp8Ibw0jLCOKd/g58FUauEPhhlNB5BJvu2ZEzXtaR8rC8m88ENSYZwMLeV1/jbHsedD8k+gTHNYh
P2zheqCEj3rqa9+d0Q23a04zOOhP3PqJXxQGBpmjM2qwzKaOlRja8RFsnYygJUFyTHcAApesF2wv
gyKudP+TVA/CsbdxcQTAU9OLM3ijZOjkhMaAx6/1aLjekGXlAw323olZwJ+LIhiH67R0JA9zea/u
V/MM5dCQyCK35LldE8lxVQ9iIEWSOPJBHoT7pvD0Mca8XwhqAPpfro+eXYFK7eTIdqRYK8e/VlBz
xT0DkLFpMDRYK1QWFLAtLPbV83mjyHFDSQvLZOCyexg02zyPVhjRT8KjRkIN5m6o1/r6MfCUvasM
i2W9pOgI6TMGy9uS5kWbA7s/uqFXpMxCX0leC/vqoII1K5GkfHp3uKGgdw7/y6RJTZJ9IM+oSZ6C
KoVsPwhZvz4URhPn+pOuJQIUay0HDEtF5TAfbdBcWh9sbae/RPdPOMsAtjsC6MogLen7J9ry9RDI
D5OhvNSFqfeoHCs13bob+HypWDxheexfQ9gDtx65ThuwniRRkYoqgVL/AvUz3Wwv3mdLmqS8tB5f
gHXBKU+FjWRdOng9bOXykAN0Rdl0KoTNgiM299lxA1oXwr0pGxAygrefIHg63RBCw+Ke0vxX6pHt
N3gyx9uXgBF2K4DD7B6IUviXzM1+whB/w5/WcM3wb+Z0cfgxG0QztGKMsuGPHD2MfZ9Z8J2pAy8d
uIdbqIE72KENHRPh1jYRX/hiShX9tuTxJCwxpE4aLbYzYaq0F71lnY72ahd8KHbYfchthT8gwwmF
9AwfetGYbJHOPhpG5j9KZj69gp9EYHSgP2FY4WFgqOOnUMnLvRdUcRnIpAu69AP6l+OfOB1JSm/p
Fe8EIRkg4zB3tM5RovJYijXSpgVNq+d2o8UEwgciHKer+umxPHR0xauC3hxLrx5XtPyDB721GmJ8
WThsG2E1Q0ha7KclwwtBtxYsp7yiDu0paiQh9copYpPgNGXcLleb8QkW+JHawWS728eIQMMVOck/
ci5eBW2H3AcLmDapzqDqsWbzp3Rm1BlyW5W/AKqr4d4VQx7eWkBjlt/78YWvUEeG44KhVerMOxzt
Oc0nnGOVDYkXVoysurOVvElECje0xAPME6HC2Zr2HmmtMJyLXGdLlKcx0uYW0nQyrtydQy4MSfVR
6aKLyqgtsHhxpxm2q7oOMSnV+1HonGFggQzYl4/sPm6LOnwAHjOqOZUtjH9eGktwllhiPBjsNiqc
dI8KXdeMsiPQGbTozBpJigJ3Ps3IidxOS+wZeAINsjYE+hvagmvOv1MW6thDqMoDFTZ6PaxXPgg6
BBDhajjgiTQilIBqKrl9LO91C+iVEmzhB1oT+KGuin3f9VjrBfQxF0TElBUmB7hd3THQ0+AMTJkd
+0CyNJ5p6JZ6UhmdwJSYRpfmGzaxLMM3IsN/E3fLoNMoRfG3oP5xi4g0WFKlQjdmCB2n21p4azXC
exswR/F1pV0K47o/8Aq+ve8NQgDYiEDccGDYySuoKGO0giFtvC7qE7AUWKmly/RqieuB+GBF55vm
QMitlmrEx8Gd1MbMYKxdebsfr4zoKVWcy9wiwN908nfYfzvEJOdgQ4+p1j8i2DcPUyJaFh5rER0X
IHWowEIhLuIKUbALWd5fScxGdUuouXpjfNITAHsy155M5dl1nR8u9LsvYcRMga0EZ/n21kxdBiz5
wPW1Kcuqzrjj47UDHyD257xqZb4VePeX71GSuPQ4llncUza3POy4dO3FvKlQ0RlIKXOrScoTNRh5
fGSKrodjweosF8zI37WnaAe75QODzwssVoyjtPXdTsxRzTK/224VXhUjAqfPcTNE9/ITa5/E79yC
cXUCM8a5g7tomDSLRoqWiYeD6G6YptJ8J+4mw1IadR4lQDcXHV7JrJPFH83/MucomXBQUydLsQEA
21iJB+QkhRZe1L4MATbzwInRPbiC7dRreMOGiBRQFsbrEENfZAbFNDjQb2nPo1uYsrLrh1aTUqPk
oUszhxZynIsSy8s1DbqYLCk0Eu9yWFgM6lCpEH5vijw2+l0V2da78WCEw1oVFMW9quIMjdONNaZJ
qfdJDVGeB4ktvQpvyIsQOftoxc9Cxpnc8+aO7gUcIA0LRJ7lR+3tU4NOyb7boh0DagT0WWdMKgag
E1pa56tbuUK2nwwACo2MqWubHX1SzM9zwBATa9T9XUJIcnUyo6XoQ0mSJUSeV5V56+vea+75mUHo
OyMbkI7m4XJBmUQdejDzboLeQIIDsX/RdmVWvf5tm0phiQc0huBGH7FaQic821ToCHizz+VM/LS3
xDqId7xPW2/5XYwLVbw6GKPiafbpVPd+to7+XW4LS/INEIj1QXSWpLp1rValVt0bBV82r9IuxOdg
8Q6SXtS4fwJFjRAGnPfuAUSLRNJtavJuADXv2jTjsR+j5eEqU4qILp6VO7Sf+Zxm28dPgXck+S1D
Ekec4IQgkb6ZKnDWYEDGMjPf/HHxcoOU4Yx5cBdCb1BMDe/anA5VMMTthxbYWJSXdVYQQAi9MH5m
Q14fCxuLaZv+36VJdKDWu2jzQA5ynSP8l7fd3lPOITanTLh6Ky+ALWazrrdPBMowA6apfVAjdoIW
wULH+S729m6T7FgK4HUsygyalsoS6vY3VG8gHDfaGtqdzyPbhguKsCFcXw55gwkaCM8rZK6ZmSOf
9TZ/0S7IzYf9v/2Em9jmqmRjsQU034xpThaGy9L8YE4+kPBUjUcjRfWd27d8OsNclq8oQM8gWe1r
6+/RdO+Qiz5/a5le+xd35QIE/RkaFtMgtxpSlBbLOH4S3cKVv+b1Rdg6xWkCv9LP37/KilZJVZoQ
74A2dXH2fr1/aqLeYqlRw01LDJgcniCyDB+HP7C608alzf7M0x3WGvLShYS6g4TVbXtUWKSv1F3+
stTARzP5dLmSawwxA3NXe4U7Q2oR4U5ZrgCBBVNONTEdDYk6C6WaDcPf9qOQlZtrhDX6g9EEdTO3
SpodOnq3olIPkEi/8RwbqF44ojlK7iyWd3QORAbDl78JAoVuUc8bQhseRupmNrPjaUKDw01tJwoT
skXV5o0wab9ha1GFY5RwCD3AO5oDUN8TpMxEQV/9iO7F5qrh+Nfw/cCYDkMl7puzERiCBUlrydtn
XFr4VBWDbyKD2e4W58/3zZGlVPY/Qu2EYL7HDlVNnziW9Lh2C75G3Kl1hjovRo6BIZlw9xP3xyBR
KbelKkQ3QmYji1ito+vzcSk8CW6erm5Jic/SKxI2LCH8Gc/FjsGrxRtwJMQfpgyLRUYpnoQPcESa
xzITrbYO1NdXmCMcMxJmbctTWe8ghDjS57li1QFMH+JaQReVCL48hBdKooTUZDBVhOhIFF6y0SSe
E0KQCP5A+eVxOqfGiz8jK9PTyp9AwtR45pRIL36PrPLYRAiJjK6PeSGWPD/02/ZHnm0PHHMIPyPV
CBq0rgBonuNX5FnRvq/6Xgw/X/gqsKd+X9S2yQuy42s7L0MzBWEVUg+a5wNLBPUJvl3WPspdfjWz
3hLTrOpeWcpKj6aa3ho59ehnW7F+U5c8iJzHiH5sYPxJpSiu1VYQ5eNTM1DNb36bN5Wqs7kts59B
LNEudupJoRNKD0FqBrEioZAXpMeOpgKdOR/vdFHhM6EnHoz3OzQAxpLmff4NdrBB6ypL69wbbs+P
KIj+91DxHc2OQOC0UzSFAsrw6nRZqA+kJ+Jnpprn9ZFOGekOqh7dh5cglH9YIWiG2RebUTpNisAp
QXJ7dmxKtfNSu4fDWQOOVzE+jNdpB6IELFSxIRNIHOpuDBYSXWS0WjPWkIwCupK0pver47AWtCRz
fVTs8WNUSFUm3b8wuK9iNjxX5kIntAyDXUgRLZUSvOtq3oyBi5USHddINGVnDRLnkcIf2Vf0hqtd
LgyhptXALMTEL2c+OIWpeXLIN51OpbHQNd1Wzpcn8GTOOjUsYaF2TipL+mfVxn/tbTh2pIEQ68j0
3cEKn84VKxm1ND3mhSXolXUxFrn5YEa1IEJ9t0pKAHdF4C80tOLdwuBiXdNLyHE3UGIMWp7w6kfj
sFZLCuqeU8AnCGBRajVTrCXW3y6hLR7+7aSEwAfWxLltk8e0vBuCubh7LDUD0bH4rnXGp5yKV2jj
An5Ox0ujaAMbSFYDKIXzxHBoW81yQ/hHh34dZW4WyTFere6sWrfC4nS1giv2C/ynr7Mi2/B9gO77
2qMV0Q0wUE3SwPWBPinqzUQxqGrns0Vj8rT5N5hVPA1GCNAfQKpY3MwmHZX5esljQ3BXwP+68n1Y
5TnP2rZGLbB1zuEXynsTeEgKsEnTMlOmFEaCCnbYkqtMz8ybSk3YLpfSOoqabhFK8g5BgrmeMsUi
RSJZ2oEyr4XwIzanIGAoFyRfExT7vZWrHtqK6JLHNSHJyjnQCMz4vOXiUpryMhwxSfUudGeqZPyW
1O7d+d5mSHcVRTDe3BOOJrRWirTzJ5PYrMt0uTvzg0xC7UTGL+Vmtdult50cgc2X+UagrvywgBRo
meRhANvyq2pLXndaOYb/RAd41m78zu9dpSztX5OWqlUdtHVQVTi/cnLamYpzRlixhqcb6B6W15i3
BDglCcPEYR6tBHCDS7mmetAYLMGBUPhrfdA8PGRqfKoS4A+egvvWrVmjFhuV06PVMi4+oUFDQFRb
NhWjuxaT4mVNSlTKLCcOY4fqqaXEr2ZXK+LO/epmLCKbl4WnX87WVTt1CLDg9MEMNa9W3TLr87SW
vhRxVTygwhx+X8Ww1jP+4h9KyRWJWLtbPjTxJFIgAAmOSqQkHP2XU3R0k4WC1vjFW62SHasP5D8W
d7aoBo0AfvJVjDhYVFYbWNk9bX8UXChiyBosTraFdRU485+1UBrNmpjya0fAeZeY90kJUW1NU4bW
ox4nmRVC/ptWxceZU+m9/jV+f5Q+TUHetHFk/msrKSS6km6+8gD0WXSkfcysw10ilirX0J4C7Udj
T0Xi+e/WNRAaHuAzo/dvp6IUC+mkeNM7fc0bZNnKvVY8tTCKCIbSCVFQKP/3hj0eZ6SV+fuAdOkF
rOuPWfwv8YnIPl4VmSpMc5aVWrdZahDzUYX2tIeKJT4cE/hSBo2Ao9u9OmpO+5/jZsLU0WRd8F8s
YQ5FCgTrjXk9Hn3jHFAc5K2syL0vImS6QPZRib8il8qqeIy0QZrxCQKEZvF/gLn77m71HnjW3JAQ
IPWLK13gfZcd98LyNO7jeFakmsgnHD2kQntuJlmcsC0b6rZQNZI4XQ1UQ+md9SSMLEuhZwZFjVBx
jgBwByXvtHIqlTcLQEvUFedUHXE0nu9LSIDFMsbMyy0+u+4REoKdXYum/88mn9D+y2CF5B23Cvve
gbM7EQlGvE0BvsEZgCTAHEgQx9pSo/HGwwnLAv6n6tra7XUbj4dO/BoUs6l61hP8/h5N+HF+5gYL
fvBJJfDaw6xLeVNzrcg0Dp6165fVLJ6KHDbZgM2zi1Q1Ne29fp2vcvI+KLXiVgT4YiEtnhb1L8EY
6Pg89aE9XTKSHX7SvQu/Ps3YeqeVeznOxikQ6M9mwaX+BpxFIWXNLwgBzkat7UUgrvhwJhCr1SEn
mEJ0HkOEOUEGXWSHEDQye/VL2g4grt+pCIWEK92cPa4HeTEhO5bcGDEF2wEHF71xIQUQhwcncKJy
eoPltKURH7FGOpNU2yZ8ULO35fvCk5evcASha48o7ADmIC/FIYIXqs1yada5yQLY6F1ivsLRcVHs
i/KgfdXgn4rvIIVVQBLsI9pHi26rRzx7HrWs+499pNYoI1DrHPz85/+NqKR7iFlA4k89cB9Plpu+
pFgIVnTGftHA1zh+WVa0itBjpo0DOlUZxlDjOQM45gSIiozHif5tTFjTZ47gV2Ut9+y/wCNQJcBW
XEcp2e7dRlJ4heWI02mvLXa89C+yE74HNx1Xnqv0dCUElgmoWpgE5k+B2BCZggcib0HN4c1s0Nqa
I8Z/WA2Fh6OQQivuix91RPTm6czYQtA1M3iDHXRu6h038vl0+0B9ajQOfM1do4s/H5fCQoy2Np0f
/wZF3XBwRYTikBY2P9kUm9xRyBr3t9TjuRAv8DMmvxpiausQsQBZ9UOSBy3qNhbFck5LiYwJee1h
ltS7XZc68yaDgnZ9LASHWiYMRIkmFjipId2zxpCYiFZL+myA9+ay3UggN/LyDauVPj4HE5GbQyXl
/AXV5qNok5aRFi7NU+V5xm1S6Sq03hYAYbGUR16RUU9tsZ7Y8DsJvcopN97oMwstyjeT12Dnw76g
koz7mIFn2Pp5cVBuSTMV1lxEGTv8GjNLrKxvyCYYfXbFzHTrIsgWyHrnOr3pnmYJPeBe7zngXU+z
+PMAnRoq/c+2zl1c6qbcB25yNuDZHLBn56sXLEPJ5HLCEgPswwdjL6RgW2ywYBd5TDD1y6QgPuuE
9TXnxFWFZpg+oUulLwKX2hXOCPJyNqPQmNsA6daGBiSw6q64gGl8g2xEQUrdw+3B4ku8AsJq/AnT
2PrsZvIMytVgI5D7fJ0TGCJx+xE8AZXCu1pFrjZ6wJxPC/3h9QuO2O5Uc8Am+TukwCEv6SkjstBm
l2rURClDYWRfVHgxzoNLLDJcTbvJR8RAvdPCkNWav8cnhXdmD9Y1qKViitsubwpj9DS/4lPt93m4
JoRh1UuixahsG6kJy2kc5rXJQZbBcGihSz6GFzA5XnFnbJ8VbJ+M1T/EsDCOEdQrI4rfhgcqiwRT
eb+xUcJ+g79iWblZCmRRQb0yp7WN/2AETqH+Xo8JUKbjutH6fVwtRSoQ9JBjQQ8YPYVwjJdZtu/C
wdPSmwCEJRv7bae0LNSZCW+feQXQTIctfn4RMO0GIjL3vtslIqOSWEpWvoTJ3EYm1w7O26MQxG6a
ltX3EI52YZPoi2NTQFvgP4+krzuwS2QnOxSzDtWQ7pEJ+PI5xzUcYvqXj3lMxF9Wk1fNHipqaSGv
ctspgajcr11Q/Ll/EPg9/g9BpAFrRS8KMW1TIdSyKIOXCVA8lQkp/CDhZ+hpwDSdbMiOgXJFNNfB
Uk4IcLAVRYk0pqkx77PRjIlQNWktKTeCkuINWZjudZaUPHIk7D7urSoBMSF00n2sI0R7BE06QtxS
MeYs+Pl1uSRtkX7awLv/a6EVDv2zAvCtKJhBYb1kqk6BgFHgh2e1dcrLW3vD+MIpU1ippmUw1dR8
PYKTiVCsHGALrkm8fFDW6ZEwa9J+A3qcvfbLvCl/mASlNgPp3YBm5mUQwOJNFnulAhIy3lLMuQfh
cTEDRA4L8NRCuEbq8LF+yTw2On91K4xSSRGGxk55IQ2mJe42fYGl5p2+k3wMLmkbt7pJPlXxzJoN
wZSWtx+r1awR2Dp4iFyMWSQWXOwSrW6v70VUFTPon5NdU1/eRQeK/chCiybnKDq0Gu+ob0tAF8EA
PF4fJrTqpGGz3u7EZNht0w/rZmbopPfLNVMB+rR9BHwBBBhCJIrqv60b7YX13D6y62TMVj+sKlqC
r6aOBrxW1Y0Xub3affJqJ5gxMcPt68f5blCv/kvTmqcC5DrvcKCiJMIj5HHg17OgiYahDUaDJdo/
qwEwWxbVSqM4wXtSmD7of8KI9eD6wtHPi0401Ngv+qFEHuT1rHLFte4hI7VUDplVdFPZcb2kUtpK
peWtXlg0abkj1AtMeV/UdEalzPRoLfgChp6GlujqFKcSctaPm+8DKiSUJ9xEUDA1GTNDIIKBANaw
fgwViDYU/77fCtYE/nSeDTB2ZMggAY0vJWpIDmHbxPn7/fFkaGJUOA11tUU0eRZj2Rmk/uYAVtox
dQUD3LhVsh3LQyBn9axjWWZ1ai+SdCC498uh8wP4TyC2+bpTz3UciEwqulyoGmT6vsXaCzQT9+g2
z2t6icQ45Lo2HV9G5BKv6oxoJaP6j33ZmGhuW7f4Gk5bOaciHR9FHm2/22HGx4oYUIq+TO/43mfI
ozbR0NWOsO0EYbMYLMGdbHYUtRfRWQhYyVWs9Mlj8cEXs1pcQ8vpefmN6kSu8dS7XJ0FEnqxFgp2
QvgGnzfppw2IgPZb1w08hudKupZh31EgRStuFeIcrPkuXQRGyIvMAif4QBx+m/GEgM7b5KSDXKzE
+j7Tl0pUiXnZNHC447RaUZOhweaUsDdsmBer6zH7F6rQNOyQz1xz0rYkaPo+Bpfy1rUlHLyze7SZ
CO8GlJJhv98HN3RO/6VKofS0peZBo4eQOmHeMzgZ6LxkJxPbMqdFnOI+/hZAEAbi/+9Esb/mKEZ4
HwwIhdSgkwMGAmD4AaA28z2zXO6SQGDwKzSTuKCgnNGVssBx7iQ+zVDqhUE8S5fc4IP2nSiaZ3Xk
MhmL/aK2qtFdjndPJrXqcMNdjVYzfCNYXbAasK/Z3JWGBDG5C7qaSzW+ZIJkFJatTrsXCI7KFJhL
V+CIVdTIzPySmgpmoEV+Q18TgAbj8NCZR2i4invIbe2jMMMqvpxbGWgluvxKTlCikmfYCKHxQk5Q
MYuoPgOKjO2rtg6/M2eB8urrb2pXd7wQ4BfxGq8zPAmvpzADXJBHWo7z1XIHF+9tXyQ9T9RsZlpX
L0nCKCUKog2KkIXGnnswhKwqO01daEmTLzKuYuuweQWuwLdKVF1pGltPIEiNGxrqBxS2irmuj0NA
RJXx8nDjdfPdvzzGzy6BlGyZ0TlGKC0vIllHQSO4kwtYV+dCohPPhTEn4Q3X6bxsmtwkK2T+8l+D
AiAkz1flOHoKxV9s9nMjj3fCBMOLFZwcsuSCMc9CH6/CtM+KUcpM902uEROg98W6aV6MiN/GWE6j
v5eYqnr++rsMEDEw4vwaZai8nyUdVprT8LB44iBKP71TrIw5+iL86FTTbJXYeSMncn3MQDnPDxut
vp9T3WxWLQD//YZx1hAXGcyaTU9LsvydmtyoVzyUx+tEGsZQiTZFgBG5knm+Uk+L3ZVJV5QtruDP
sdrJZ3Qs42fRSHplbzSDCQCUmCorwRn1YoFnqCL8HuXIp9g8IXq8xSUYFiXHvHWp/Cb0sVafHnJJ
RDWpKi9098VJG5l1d/5k6GXh5QK69y4J2d4xC/dJaNY125YX2dQevwLzLFrI5q+/+mjSSCUFofob
U0KgOrWBdSYwn2CP6EFw7V2QqooFwomEB+Tvpjayaph6n72DGSC5+TPIchUrtaSJOtefefjHIoUg
sjda0GTZbSTRNN62gX5xhg6IWz2fbFDpJlBcAdDUP2xpq+hEyDx1GdRyyhl8GPTiIreYLkwClJ2M
ojtgoPKpXz/MP4DhlNJgMkv7D6L7o+6aV8j/JF1tY08BWMuqxGh/6d2+gT7kYzLS8KPHQJ6kgoRJ
w8JG3LERBJWOhh0NAZFK7xnVBxYfmnbY9AicxJdVklcJ7UKWcT1t9QRg1IoEI4ED9vJKWf1PGery
YqlDyuxOok0fR2o8h6Mh7VQfHcpKnR+aQopMTknmiHfM8M+FNwp+WABOBR28cuCjMXnyYbC8lWWd
367YSfzvt/tpcstNmuRhn5PHMZH9SriLAlOiG2STgvz8ab1UkNPwXOOYKWbdTWaxiFu8OfHnS2dU
C3Td1h8TzYR59daRiJtj83zVWIUkljge/icgitKpceAWq6HNQ1pjqGUYfRsWyomv2PJJlJwvvn4M
GXIeEzPKmgp/ZrbUXsfb0Nmh3/Xs6ND8GYJiakn/rxXbW+Yfhqirj14GbdGFE7vyo8/V4iueX/3P
m+ivi436oUB52Mnm6J3B/Zy+g86rhA5ZgaM2s6RRv47JzBqkw1aG+7quD5rKVPoInzP8UYhCGA6Q
F2YosKTjAovc7euEvCa8cooNOt+E/q5PWZFJME16KZnI7ZEdptIN8qFmmozsnrz2Mhu4g4s9gRIw
xALScshFMbkQnqkHGHjNBmYYZTWityBvd6fOOf8B3ea3Sn4bz7EW/sN0MsZ13uZDV1qu24PtDiza
Nd+hkKRximH3G9IloTOL3LwAx6pIMeNwNlaE1ifc+P48zGl5XwXZavyM1lI/mPd0yFKG3nFF0rOd
8QfH0zQQwEKBrO7YXpTB0gzM/kZMk8lfIkqp22DSv5S/fghWmN3PMa+7AWXENYB/XYnh7lcWLFwu
fTRlBr7bARvB8JqHSknwflCfUj13BbIwQ5ejvVqu1wKa+1DuYs1LFtUIn06rQ5VVi7FDCfUnmsNl
e+8Z61N+U32pnJeRBLFZSB/l7O9VU32/miKWZ+TEUjVFPYzdJu/z+1PZgTGogkxSakVEfdwtcV3F
Pzbm/flAyewbunGRF4YB6WYkR2Em9llRuKHXbQiRSDyJB89Z3dt+J2+Fg9MmBlOYVM85gwNiftM+
3GsLaP8SHi3MlmnNWAtmJgu29W1oRT6jsRkdc+NX8+V/LWWZyABF7lR7J4DlgVZP28ev/A+k8Txk
C4lmT5kiwLycqcR2bLu4387Wjmk+8yihflTEa2+2ok3567dNhcNqA+k20hQCeLyn52kXs2VZyWAK
otZsvq1pSWOeO9aZCMBdU71M4p2aeaTpoI7rsYWvlV/mvwu9hwzDPb9xomyLjt7YJbCmx0Wfuqm0
pP66GnzymnstG0MkQcshp4u3g2hG1vR4o1ajvL7UgTn7bhiZKLMCACkZ2KxBQXx+Dm0/UDaWS8Zz
h+t/oz+dBfbqqk2DUA5DXRfEFZ0Tp+jsrQutetJuio3HJOa6SHEV6jL6jDcbLiYZuoJu75ITs1/Q
/U4Eui5VH8eFUAvbtD4UeRkeAe4Go7W+T4ucqUkXlcyqZ4rJRon9e1smwphyoM9yJbPmLuZoiS0x
iqToYLDNW5TLx+FQEpBROf2mnK40gEaOwlevoZYMJ1Kwed691fd5jzopFTZ/NiDaa4eGC4KHVdeY
T9R5vLfkZWoPVVfCT5jRp5cpQK1brO+jes8t8mhTePbMLWBiJ64YlRCzNC5Dq/Zqm+Qqc/CUBKke
CHz0HvMb93m0zeWJ8+EPql74m+g3SGd5AE7SgV/HHFskQdCaqGs7GANK/Mby13oAISlviI0J5y2d
gTuzTmY9OjSi6H4AbM5viuUeIXcjNOXcgHOCCGlRg8cltCuJnePEq+J3HdXzRj5HV99MdwjLMxKu
EKq8fsxhAsnT1qeFIhu+EZGmnmRBESNmNs9nBHJa4VOYV/UCZrQ9Bs6iFtsqbpvvxr9/uzSnUtHO
jRTe1jCsEDoFhA40pnTs0aOIjFjOX+wEPDq52Z+aVvPMDpFw3hoSvz5tCqFnz1bxc3WgkaSSWLO1
8lX1Ntt+++SdP8OFjBYRW2hqz6eVbFF42HcEgz4vXlYDVcoNKHAguSkwB/wWkE2iugSyJ8JcZMlm
AgatW66462NgHDHxtLcyY+yGY0kTwH0OgyplVhcNzctOf19O5kZ2IpOZWq6MOX4ZrqiPAk6sMObH
ahu3etQZmwqgdDzcWyezuHWMfb6A63lptH6FqyNVI1wVtl5ADKNGhFvNgR/DrlYv6Gvz9oqa4Vwm
e/ZtVir/4OCmZDi27QkE7AkMze8cNhaJspcxrE9U6G1FWiYg140ZyDW+hoZ0x8A7O66aILYXwoRG
yaL/l4eObYejX3Pf8LitYdYR9nAsN0JyU+e0Is9xSmISFlxUQSdz38gYjhxG7AruUp3ONkyLEbVn
K3tqtwF8JKux2TUsg0DDUXcbOz9rvtN0M355cLqyBAhA8zq2S526S7/FZZEWxESngb1magAPLKKF
B2lwZ6L1hDs6p74rf+lYsAOek/bp2sIWhmGOod1CPOTwYOvw2DugLKezVdv5tJRZI9Vfd9uRqL4g
10UlgWO0O9kumF49/AZWeAw55ghkSnV9tj0IMbIEe3zbehonQ+HX7+8V6Ws1hyn631b+E461n68d
zl1nBVbvjYqBy0YSvrp6ZHfQWonFWHLzqZKB1au782NAqANKyVGhHqefyuzZoAiR8yaEjba11HDz
/+qLK3pO7IBd4dILtRe756+31bPhlukM8LEUt9eMhQ7EfizusxEJUPYO/vIsoPf7lcBemAyPVqpN
jNzEbb8g+9qrSPQ6orIzjGLx23rPl6x6MLkq6huEeo1QVNzTf0p6Zq0/j/0T9DKU9ZOx+KfXhJBn
96w1x94ALKd9JZosJseZ4ILmk+zrDD+8SF67PUzHpM4wwDT16p8DZCw79ypHshEwu1g255agyyHx
w03g+tnW2p6HU69cDyhpV2MqvNa7s2c07pBq1SzaG8YJvUWu3Bzi8XYEfbjN/w2C8EQ31L+8lsem
uM3MBph/xA+U37Xy11tgSC8e3ZB0HodzdCH7M37R+wtTPT/Oc0ThfZhPrAiGHJXMIIrvsCFUv7tM
pY6hYIwRIeW1AKCcOyKnyeqmHfV4NIOhOgZ91xIpE0UM5GV8XkWe/5hcZvx/M7l/STkj9IMvTCLe
hT1khI4+oeO2ZgXTKVCgNy12alNKrCG92mn5MoNJC23wAoKhqFMCs264dK9Bv6QxH8WkM7JJ0Xtw
FkqxrAAmPYbdMMCh96hyY0IJhgXkVEZyPML04pz3BDuGXzzmwYNVrrl57zR7SnPFVR8bkvGn3Wyq
c5E7mmmKdaco383TWaMtLsve4kpA8NhjVgTASuiNcKn+8jyxfxy2O9KOMYhAKvVJNnGuevSrwdVa
Jrm/NP2ie6soGIf7NmKDAkphjgkUI/iw+QgwX8tBDK+RVIyZFjgUILU2GuZNji180vgJZGiYWgWR
pSzKfjrdsuCbAcIxN4Zt/Pq3YpyOQs89yvApHs29pGYCxhkYNUqc0YtRrRnpRMOMtJA4F6MozCa1
+Mz51Z4nVr31rrSMUDk8KeEyuGchU6mv53t5pXIqJaPpZ9EzWAg+oobvbqmUQjyADqpBSP455fst
ZbDzJHLrKYD9P3zj05TaqDLQc0OTpKOeCiFO1XEYG+ONzuuM048r7F6ND8lj5x/1+ndZv7vKm6bg
V6MWywubvbabnsZBgR1wboyu5wDBwnIlak2Nwyo+tyOS1tL5yEwldrGuL3qNFkfApBZQggS1xllK
cNeUM2btPhVkiLeMVq9CH4YSpuY7+NALYIVZHAmtgWYRImCd2JpupsBkuIxTq8ENXPpq+kn+RYpS
9JrBaMFJuJ4/yi9Q0a0J9VtnBnryGEaAKu7kgTPcRYPvo6dn86jw8eGMiizTMYUqPkbwMgXXyOXH
l6WNGmCfHt7E+LNRMX1DA/PYLB7aq94CIqAPHgTgWw88i0i1WnFbeFmSIMa+vQXIYxNnTYlyfXFh
vvXt/biloBWXYfgR+9KTaD6U/BFHnaREJ+O3aNaRdlJyq6mV+w7/4KdD95gPgo4hsohhQPEDexJC
stYnR5GrPJqxW3mxQwVRxgl1WzPWd3iguq70eBinDQJpSbP5+isGfzwSHdWb9PrPe/DxQ+wd+y2p
4Ic26iDfuiREA6Cnmfh43n/BfFMAvuceWWmhqR9lBnMYSmV71c70qXePN27VzDryReX1/dgQpwWU
9Y3rTiLAnQP4ZoW7+8j0r+FsZfoay41H6LvqAuxioSgDxsU0NG8835/3lliKPklbP1NR68bd1+BG
0ahnneVzJyx67F4RdeZvxq4VgnXv/jKhxHLlPjARyRTPc0/F6Rh2WbW4TiQfVFMVakOKzeBZEvBG
KvejX3M23Pq9mn44uPBq5kIwpMQ0auVrfA0ciLL3I4Vlv9LQLPzcp9+yKMhzMi0QcoEZJG53ITQe
oGNoXSBejAidxYjzK4u+ACV5+HiBt9JELPXrP4IhgvSdrzCMo6Mm8in3dr3JVdYrKYjOr7Yk6C2M
Hn3pvzUI2rweEiqsEcIq4krsp7lxW/FImG3hogR89rrVqzLy86R8SN8HRg+sX2US/2Fiom24B+K+
PeMJwKrIQU/bi1RWHD0uWKwMv3/73KLhr/QbRVjlyDbTMDV2/brqDGEQ9VwsK9yW9oCyovE3YT8o
rBe8jXCTNqpf85w6+KWWqsCHAVxKXf9MWpzllVn9sJ8IH9Dh8Xsuxy7Kp87Mb93h8VUvI5jZLh9N
D4kMnrlfZOWqreWVoVEXomU8yN/6d/EC3O5JmQC734ht+AbfXxehQTuKdsNygi3Mn6V1xGg8Ps08
42jEd5QBeFkoxchkApcOSdaNEzCmTTQpYVSf1JpR93cVWwvzhqYdHuCWgdR3m1KQEqP5CCfl3qkC
wQW5JZLKaUuGwrBEsA6Mu0oy2kMYpYqJVtvcQ6ng7iuZsKbMfya+vY+r7IChmFoeSz3yPMMtf3gT
3Rc73t3GGwj2sR7yPKBQk+DNFvrMx9Z+7wknrb2Mu3AC7nYFOBYNsgBJ+74aYlZ0zvE6oSsy5iDJ
G6ODr5weP+26y66ddqCIxUfXK/T1fL7dVU6TLNgslgRlsq2L12S0jFB1xxXLbHxpasKPtmZQvVdt
ual1zm+DKVUes0VbxzJTozuiq2sNhp6vmCKLN23UjZuqAMig2jzU2EXulr6Gm+fSfYhjwHLjFKdo
s/6AgEMMUGe/uA/kkwye8CK/oGJBTsfUs8OBOYGyXhB96rqVhYTYt1BMKBB8MbsGSZn/iUQ5KJUW
Xm3VSg6DtJagFpZ0Rf/j4dTGVDJ3FFzEZZLrlAJveo4Pa/3sP71lObhm6lorqv6VnUbmCETdu8ml
yZYOvQZSlmtGzzwvHg5ddN92lsDfEmqiPZvsbhSVpbhrPiGU2hPKn1vO24BPU0Mk4bW8IPKzZFRz
Iy9t+lkZcyrWuDchtQGeBJJUVo04vyk+kCHvs8o/nd6pNoiMFSM1OM6L3m3ws6vylcTcHgJ7jUf/
Uge06+qPTl8CuOb2oMTvPc5UsceKumkKcv73Xq/U83AA6Da8Rbnk2X7tn5QsST+TeSg09D0zRtAO
XNuEF+daKPL1dQhRXRak38fNTMGZE9WLOAKpd3RHttC32M/iABOisKx65wzDG7SrC8ifV46U9rwb
U6qCCOFkTvVOinaV35OPdxktiVD4iQFgczMkZZraQIEw+hBCiK2ce2cZrCheUR/rQSNtWlIVEN2R
BZmZaqwLIohA7UNM5EAmkJiVRUQikojjk4tx3leEunkRbuRd80m3A5umI2daQ+C3pJNfvS7D5BXi
H30uLk053C7zpeJ/DanWOsBKUQJZQkETTNipmTYPpOTCfpvcUKeZYChI+z5GG2C3wktlQKRPcpPd
Wa3ZtalgrE4kV6QeRKLsrBCfjXPXW5zOZ463K1lT40dLM4eNpM1e2jkCbNajvA5Wq2v48LFuGxjU
LArtuZtqiDDF7MzhLYYhY4yX2C7e6Du4GGpchKHlD11W7665BpNQdUGipozaBgaL2HtGDRU68GCH
A/S4T+y6IvLMOXHA8v6AGXqWbfBL8kt3TucJ6rPeIUTaFAicvNvcrFv7Fbux75S7WVxjYJP/xBff
eglkKA5DegphZOW5/UzDyLv4qbBZpBT9MdhkLvqZg3Nc76Xuq3BKD0mj/rbnvFXta9cOMmaegeZR
wsJ1EzOwHhgXeacLrmAaSS/2Lr3weXCq1BWeAdYhkdiLX5/Q/e7Kl/K2zpciwtVxy64BUJFqmt6L
unI2v2AGwMult03u1d0Fz6OVEfihcWAG3MfYYU3f82McBI9y4QpZpuhrF3q0yAX3tBHOOus/XQ9g
GmHZ1K6uf7XEiOoLrBwN2zw7w8cbhyAhNuYbiWVBZ8oLLV56cQhbjPPo4cswEqM7e7GMQLDys8Nq
WvcrWDlLC0wdz8A07fJ8dQObMmyM6SaghEgSei6O2zMQUlJB9BSfH6xQ7Gd6Ge4oUdgd2E6RnC9v
o/jCcqwo2UyDVczWMHemhX/2mJmy45qnb3aFS8/N0pEvt6dSqOo5e0vr1gbQjOR2QVbUZ8AqjjSl
OOWHKjljQbfaa5GCgI9foHsQatl10Ph2+Jt0uV0WlL9SjQmVOLH+P5mWYqmtGh4N4XoINF08drS2
RXCxrS6FdEt5M65YB1hC7Usg714aTqhug+z4VIM9YKiewGupsNjwj4x6pEqcwIQM1Cqm2CxNrHza
32FoiV6sBXRmkaGgAlyFj1vX7yLsnlJ/mZmafaViruZmM+RPtgdWr00guuzdmuC7tnLiOONOo/UI
p1Qe59kU4XJcvroBplncrKnXQdf6PzvU2+8xa0c2o4X9lQhl6GMK1Nb9l7SJU/+KY3yb5g86avjq
aK+RUI3CKD0G5Pn99PuT21Br+MixHMI3ZAPmKARRdu+KWvNUoPVCJJiwhEcDIraulY0QAe6r6AuG
GzApSVvneNTXZgQJKw0PBMozIegj4Q6NXvj4q3Adx/m2mkBdGsleZOC8bfQ+InT3RdWq0mV3Zvve
Yz6Rhk7KELSrfjyObWIYnYCZK3MHBoakx1NwAjgFzJuen7Tptaj2y75ZJo6CcBaSi21qRQ0bSJF8
z6SrXYowRjoKBz+vHI/8ZcK4xl/SN3i9PECdJt6M7nm16hJXxLBHL1wq1AG58fLEYItBz08uDTrf
gt7lo9HdGSxRwLGg1RO7A7jPiX8Z/n79G+dQAqK63yRwTzeT552nI8zLUeNhS0rlfIM1z1fxblLI
oFkwAMONyjQtIgvOFGOeZqSN0npYqIG2C4Z+STcWYZeTY7I9ld4MpWWOJelS2M09aOWghUzKOOvE
5QlH8DvkxJ+YVqT3mBsYbB6w+VJRx3ISKcbaw53XUN2LuFWGbE29FmHNqgev1/DmTh9YF5n1i3lH
aIipve1yW3BAOk3/8GRyx42Wtbi3kmQwcI2jP7BoCAOXxSTwqOGif+pMvDa3RX4qC6702qYmdL4W
7IVZWr8j+B325pRSnAbgOtcuJoXRgzKil2dT9jA6m0cQe30JOFv5kWRWUvkWmNXBEjPuXRqhx8Nn
NnJDSUdKbdIH93XADhdjOlP4SieaGIJLggEXp8ZPil3snw3JNoj1CwTzX0Sj0n3/or9Mj3eybO0Z
cl8IQVTGoHxY+ALzBB4M8zwTmTuZLzh2s4ZO5VtkOQHFVP/hCRsv8EVcZ+xZxXwkYwRetXresOFG
WX39DZMo2FPq0VKmHtR7wT32ENT2uognfpvw4poUCTbgpaJ1wWPdxBcuJa/cVPTOUaXy7QjVGgr2
kF+qOgDDBG6wIQVk4HQ0kLzlZ2L39olgIPMt6KvFGLS5DHFsw5TuV6NgabhWP3J8kpBXoAZagiTj
IZ5PRZC4/PXL9r8TNFLcWpgoNFaRSkzEPl6vSAdGlvzBzkeHwChra8z7MGwcq8vwzrlS3yrCRI3w
uLVTKRSF/FTMB0+TD3tYy3KEkCwB3E+winDEwEC9HEArCKlKwy0JK6VTmDFcPQiKdQbKQUx/tQZz
vzhJIx2WLLOPaIa4mpfwv/Cp+BJoXLA9TjS6PSE/5tMOdRH5id/t5NHMIMRrnnRrrgesEKUWhhuJ
ow9fpSVFAUq3KtL01DLjXlq+ln+3G9dN6qKpdQmrEI8hpm2WOtUIN9XqnD4bLWvRaN153LgqHjh5
XrVeUqFTjCX0FM+5T57vdQL+0GhG0Vpkk78UsLJkdFSwx1YudacDgohGL2PQjpqGyGTS9DpySksj
GOWga0RgMOaQR8xSfe+GVWDEwqvxEyOXiKeasYO7B9lwjsdvdFUMgkuJ/ypFHMpI3mg+7e5+P4Oq
4wUlRlVHEy7pjaimWLA3dSinxrXdzoJrX6FdV4f5L4+bQTrDA1wVNjBTYHHhtkhXrlV3OpSuV22H
DQSZ5mCp42VVJ6hmNNDVOxkswUV/1R5MsI9sIdo4SQnlTWtTwEVqKekZqKU5gWjsEdWU8KBwfc85
yPc9BDONH7KMz6UyN43IBj4Ou462K5V/Wwwa+2pE5gdbXA52Fft9BG+0zUQflf0t8Mp3L8J1/9gU
W5fK96cvkbQRg66i4dE8M/PMz8AZcmXRbs63s6sgl+hMPRrJ5JbZ51oMzN6baJdw6kcuDB1M3bCl
0f7zOl5OHJVj5GQdGre8VpW6XtJO4o4xiYpTfRtMYIs5+tbRkk1VlQmXXN6N2dC9SyTgADJlfglr
5TYmeMm7LgMwQRwvPBR7S5IZ5Oskt9BHeoz9wjj4MsezRi9S6L4d/w5uot2Iczq2XHj7YzrK3t7K
x/OWNb0BajBQto89B/WcvJY9ReZKI+Z3xuvk7Ucu2lewEcJf7JvcumrhytEN5J7saDvWzvosXCQx
DisvbJEKRIBS9gwa8Bk6bxd08Gh6YGLGhcoUM5GjxwcvKnS1B6Ibw0Z0dlB+T69fldBdVt7Ip1mB
2bF4634ar2W4wrhRNz5Jl/pfA1T23ZhKSvNCPfReqtpSYnViNnRfGunbpuMtKTRJzPJiM0jRL3CT
/KhB4NFqP6BAmkc40YRC/jB4amQ3QTlG8thpbbWs0Smp3KWOEGnVFdew2s55rCMpl8ZaetUfIFMt
3HGRvbxERjrrj8hY7heCNxD6VmdvC2jkFSHagzCAu0r3CrPDoO/XekahVgcSwO+fmwtU2+woz2Z6
bXnZMqo9bQFg8mrKq9lGIAMER4g2s69hjyKpwQfX4NldxfXWFBzR5gLP7QitscYXOA0bgiOiZR0Y
rctxqxoHusJOxt4kDwpTxoX6UIvgbYVwVra9tCKISOmojD2XzkSMUTN+GJ0o2Vx/AemeGnrLn5wO
0iCODoOkv3aQR5M2K4v9GAUI5p9vtv1FUzmx9kRTKk6dyCmCCcwe0E75AfKbyx2oEbAVTwbVkEsc
QSppPyTVfCReFl/fBD7+dT3CN4i5gz+rdrCU5SwVuG64LP44gTHYiW5LjNzSFgCLBvi/LDwJYMHq
JpuqsfciLJASfn1HqzBR1CGLdAtLJ/H9B7Wnv5H+J5QO8l6HRDq1DrunEQZQrtcbXRz6dCN7mp6y
RvkNIIVg/7v31alyDwkEfxBjqJZcOeeij7X1H3wGR79c7v0KlUiXssp4vqlk5W7SL0B0QbLN6E5X
0GaJUqF8G7/nMoZ3NnFJCBu4ZnuETtKH9ltmMU9w3zUUHnh1tfCz+cR4UbdFxI0aS3zy1ZKjjpfu
85hfdZ7kMYmfussfin+WolRQ0xmp9AZHHH9FFAfzquuLnDb0YSScha8nRb5MFJnZzw5yvi3k+U61
FeoHbyekpNVQVpMKeUXw2Gg0nfFYwmtqvAGNdyC4TUs9qA22B9IadYQEdzSyOQg9E6mlAmYQKXpe
k56tHbvx4HwUvM0EoGSnXa/XhcC+jE+F1Y4f/FkkSlcl0pwwoQyW6QWuEaNZy4eksCSvPhd/zHuU
Sc1C9nDLmeTUVq0AVTwsO71rVDl518GTgj4iGAhEUpHELpQrobbpHZXAFlctSWhyMtoBK9CG/WMc
gevfT81/k6qEtyy8uCREXos0VZyvIkigUp0HaDSmjHi6HV5tDUT+jxHtk7d/ZGSj3zAbesrrDOa1
09r1X+5Io1g/fo8RjOotzuCfmktIZCGV97UGdVfP6XbH+evOLyz8vSLugM8peyRN5a7eRmcYSFjG
sTAJagMCdWDirMZi27MpgckVQzGxj/rMQDHHbSsIWTStg569JfM0Z0DXe26/LsjLLF+6vO1wUuNa
tFkyK9nSiLLpW8wFy3HjFjN293gsyzF9nLFzJfRp19q8wYa6JZDlW47CZnONSMYPrNi+PYHDGCNv
aEH5jlDxeYr5YXPNQg2SwW3RSrQca27EPHphXtsN+Asjf9sUlggIXiq2Mt4jkwNYsbGLj2JIord4
i9juOVfUMciW1Y8ZLoFYQqN5MtI9la7o9q++2HXHmHu+5hFSqX5D4dcLcaNzJwpo5yW08x0aEVE0
Uimr1T0vZAJZ0TjBfOzZ6p25MQnCkoWT6p1u9x5veONcpHB1vnAdPiPSAW95zVX8Atn5ystONmWc
1bExxX+emLD3wZ7IQ+z+4h5ol7QVdzAOijHKcyPwj2THi1Y54ICRhlXPvEpoclzEDb7+KD9grgll
wonmxPq5Owv17V+kEMCDrUPOE8r9QZrhGkjQvmkLYi+NnAOZN6Mw/UR09/3WKiAjr/OyCKhbvbu+
UCSoXl+ydu8GZSpc4KeDczslnjmPjAOeYBDchoRq0ghoSDXvGXE+qJ8Bzrs21gYpNnSDSUwcmAid
FSBln90nuobow45ZohXrKlcUiEOlANHRFgWYr5u0ZsJHyiQOLjUamjdsmrs+zzGgHY4aS5DWmhYF
eBrGt6I25EcIMfCtDYRTvVFcSonrgVdaLVgSd9mMJkNE10YIoJNqyXn9AFqr71araeiLAEc+aDgG
WEwofy+CxAWknEqzjsaXIU3Hucj4qlI2ctxvvTHhajwCwAQXl/AG82Fqr8fusgi6J/ZLTcrFpkyA
Qwj/D4vi4jyr9DBrKPkyPQRuYWA/39zWG2w853dXFLrZ9K+iM8G2fWeraO17odJjWTthzLMJ9exC
mzDUiPtTAbVV93di3fgvDtmi3qgbxmnSpns21/bf4eqZMgq9QZXrIcrFKilQHv6RS0dbb+O7COy3
bQCI/i6EuwVq3EhsO4IdehfJ9H9Vox76Q+1smJ5MHCL3Tkx73Z9MQWNRr21GtpPfiZ+znEINpUqt
UYQ63SaNjHDFWBaWIQFv+eyUjidgV7aVoDJ+DUrZBASkvvtDpeV2msrz0aJTLvxwn5J5vqOuoEPp
Nnq5yfGH1epk4ZnbrmXUOAgxsEaOnLNRkzhTNEm0jJuWTuvENX9kjeFz6MSISuRYJNiot1IlxbWn
Ssf95IsSNjHtDrk5AjIKqDpvQH2kwfA7XhqzD6Jy8eGyrAOiHUQgZQcKjecHi5f3Gjnq3kSxfgKi
c3WIlYDAkDeutvTZxeB/yjU3nDEuzhiEGuJNBDB1RKqibMbD0kiqgxNWQODvyTr1RwAyZsO4X7cH
/kHa/WUuLdH+VJhPcGJGJmKU3Iuif7Mgf/lEq4MaIGE9epOcAr/S8li8wnEo08dcWRyts2rnTL8S
sFatCAS+2nKrac7oI9o6hn+EMjrpaDYVthJbesSdSPSAaJ6JMnxI2ySzwtl3D4gLRyKL0cBTmSUc
5ZcaL5KF7sZykePfad3/Jj1EgkpoMWdYVAYrKlZ/7LP2jkRlFuMRi+XFHEaXsM87zrZC63kUimF3
R3dIn1LCx5Ksjk8JN2fz7+kfh68k1wopf7yUV/a1ZIqtkKqnAsOt8BGxMav+OahFGADrd0fc7Kz3
vW9Y9n0MMlael9YO2SwSlQUh0yWVAaXARtWpmHuybc79Bg9D/RkVtkAHfar3CuLQ7wdtHzNImIDu
1fw/NAmk1E4azxr0Lj2UuaEgnbaXAAgeLzgXrP72iPrL/r2glAXLatlX6265zHUe2bXX2GTAtxI8
E/0Mj3jT1CbZq3CtNKFpd38rBGXvUAieb2dlnaQOXmtmBtUV85Ltjj8+n5xMYLuDhwjpSUEp3Lx/
qaNExmq0yYCklKNY2wWFhu/UmxcSsCRUWtdiALQQmDB8dUmnwOiOi/JPcHLJupwYXL/MR0olj1jP
37u9o9bZHzBI+7WzvBqhOmunA5BhemygrMPrzqt4IqgU/IICn2QTHxKL2yiOjxepiATrt3c3N+m3
1aKwaFrX1LJs9hYXxDWCs7wZpfTkK3uV2ABwsyWU49pkutu10y4+1WXq77DOrZbNh1Ky7GPQKUov
K0KOG1b3E6RoUbOC0Hpg3++8n99BCwXBTb4B+MZpekxi3QzdCnsv0T+RcBrPj3Upnb61bwc0Edmj
5MQxHFKhN3dmavn9K8JwsSeacgylaO0Mk3tEPu9Wd09bGSL9B/luHL20XaHM1ROWJmYZZKBfusaA
02DOWNInxO9n9P6QITmQJ2NoInE7gBeiIniLkhh77zzX2OfY3Ps+lzRjVRIKnmFznlKhvupT+hfb
gfbxo9J0/MH2wl5jSVGW/VvU0kYogIkIrWpJ8L54Z2OsNEwaksc/k8oFlNlRSv7ryanB8ul+7Q1r
LR2wMV5SfTAQzZHOPop6IvTikR66sFJP1JCl/RpK9LJpQ7gnYq+Th9Gy+jyneh43RmtsyEMdh+TC
/hTupqM8goWLKk6w3lMxk9Ur/iCCZyA3qZ3+z/5JOlpOBz+pR1u8g0n8J7AB0vwwbNj499B/hRTQ
sxejmoOgZrR+emE8pEw8E6yBo689iGN2j4yB7fzGUkpwtZqV+9YIOa4wpdeq5Chrj759GBoi882r
oBCNDTX3dhgEMPBaUAW9+mB32l380uKUkrtVLr+cWaSMg/5MpxqLUSFveL8DYO1bpikWmLue28yb
13CTRY9fVglqXPwAxx3k7Ybxq/YUq26oRuIMTZ+/EXQV0p/ZYNGJ8Do7qsM/HBqX+Ho0DknNmymK
Co/XuxCRaUx3Z5RYx+uH0LS6imF2WYyu+cDGgOxN6lKrMxfJOzq2Ox9horhEbDStN6HrsS0VymKt
WBZdFa30BEwaCw5YkAE06TZZnErOaRmqmiitnauzpEuTbbt0PetiKpWZlk+jMT57KcoqEsCOTMqM
xFvjgJ40St4aEfpymqw2mXKJhOT4Z0Pg9UPpgzVIQWqnIbOx9RG8+7adQfdjvxxDE2lCK2CAwUa9
ickKW2VEhZ1HeQSYPvblnXbhAfRbZDOrWsl+ITu1aDjFFucFLr1UQLfNytY/G9x1sOVjcBSfGyVC
0K1ShRGCYdgpmWviC//wccksK5d463V58N1/mADndS/CQ7B/ZxxmaqOc3QjALjpaF8h+5V+9Yfiu
W3OtBLTb6dfuhTFWOpbc5jnnb2UqUKr/ysjgjz9yuIG92lFDrYbTxcIc8ufIt3RtK846UduO3yb4
gQswdRttUQFtP2pJLmqWp4COfCXHv0LKD1mfFr8UGjk7n+QsKGZs3/isFyO6GpcM9YgNuliKPgyf
WvwYx7wBI6d6YUiyFSE1jwd1jlg9VDvaqQQCNI1gvoJitrD36iHEpJISjJdhf3aTaPusoF3/VbIK
V8uVyzmmk9yFhr/nJK+/qvY4FbLLWLqfnGuBSMwy9OaVZOn6KvuLlvtKzQVug0e/8+Og2W/29INj
aiqtzLbSAnbN8sPUghXwuZtU0AIL+nsFZs1orzRJRyDbgOA0jyTreGlOYA8i0rXynzzaZXeWqeHu
OjFjPM3MsYz4hhBwgbwYSBri6eYECWYKDmUioSoh0tdSW6A0jt621XgBOicEiTYAGbeQvillgM7S
Tju/GkPDWJTYta6iIXI+pHoP3VDdtmDNEi/8MVbzZpD+NsMvcQZT//arOPK0cjAINQmi7X8Yhb4I
eiq78p1gzCPlZfZMxDOR14t8DSUf6fPgr2QUs4fV9I0SCPlwL0OovAgYHvTza2VBIDkJMj7Ytmps
LUtF0tskmGRIRqmN0dzL2fGrSvA7kagYr9P0KDR4lgU2t9Tn/ELcNWyGmi5cPtj+RVulKrYWejDr
Y7q7zIRE8rIic2qSd+Zy1vMT2KYSppo/pNeFu+W7+YJDUnIMzkT9/wVJHh/CAy9zZO4aDyEKNMg9
VGEZWqK7AASxIfabZD4fof6++tEUQ4A57fkY4iBRD+iRbtdLXoTEEX/E0zt/h1q8iTYW/vmantzR
37IghOPOKj+oEaXKSFU9p8v1nVv8t2p6thB2tSDL/PmIOZ+LiyCuIXjnEOcuUu0GkPogWq+Rsho4
hrQbSDHo/ZKvQ9iYk/ErsjeH4FHgnsyeQv2RlFLTq9l7OoJp+QAKR/O5koi2Nu0gttiKS5r95Dez
XOeUhe3xbGUn+3JiBcDjiBAqHqnv/h8zEkTyNMqXqEiTPg5dKzwEAcSe+0dGLW642tiaBXjXHfrO
6l0+4cJfgqdb4WjgdXs5XXZtfc/INfxfc3/4CaTzAA+gmjMyUhwRnqqMgWhoWTyi5aWdYc0jeF+B
3XppHdNP9WQZap85fzmr3m+X4yGcRVfAYX7kGKtCXLA0KwvOS//eVQ3+vr5V/HvS3ItUK1AVTp0X
9FG4I7M17TlQ/7e+/Jjjm2TgSz+YVZNYgPVe6zSvxqDB60SYAxaQAbxJRBCKMvV/9L0rGzDSJ8Kx
+eCwWW8l+AqWlOIwfbd1u1xJ53cckX5Z7F+7XsK+kaBk2F8gtTDaCPiL9BrP8tg4ofo27ODOi+NY
nVAnxIySbUdEoeRQBlZ5uUscGruXx0RPOZZXfN1hgClho0UH1nn33+ygnPFoou/Zg3Pk/5jcEBMQ
kmYKbWnGXUK5OyFtoAT4prQnr9jT9/9AaBNsU3FzZD7HvsIxaF+LlY4Nk3yaRVq1dxUiCc1sFYxM
GxPZXYKO0jf/DmMMIy8sS8ByvHPxffmLLREiQ0rlJtx8veFZvzyYK7DLkc7W+CSskOwHkvMeRvCN
i7u47kEwLsmmMvlbWnTblHdd/xkQsqqpsWwYgJ8b23DstsRrxRqKvBGIwxQ1L7/rjqZ3+FHV2k1E
IayRT1trQrNQ+fUUGfiRsGY0Kjfg8GwNlF7C+RweFb80B5FmBKSaEPvpKAXXJikfSRo0d41wqNIN
keHE4mW59SWlr142+jitmPEw7+uBVLn/y3leyVT7W26QiomAH32juEXF0TN800yQedMIz+GtGh0K
KDjMg90ezRZ2XuS88fcmOpqtes4JyeZrwiEJygAfrgT2crGZMre/XG8m21u36dWVWcbW7i/gGIs9
q7dhyA8H4Swu0G9vBmk/MO9aoEw7dAbWhjLDCN3oLTXgtOKVevG7EM/4yLqTbXSyy9UWWQ7z3f9a
C5xLcKyTMlJF/W9bdI5yvxJFF+moYmEUaW4rzod+sppdvyet56fpxAuN5QGQiSsVdoifCfGMK8iM
TnBqNbXc4G4IGE33Tt3zTyIcBk+TjjtJcQWRSGHtG3AJgA8n/jpA1OAkN10Xr+yyHl7deJY4HcId
nPX3ym5rLA49vCz4rOhiawLW3FYRyLEZnHtevjEvMHyZrloGG45BVxjo7MzSSLk7W+/xKRsBOyEb
TPzKlloNHvaQuCjyzhwmmeEZS4JY8aHrbrV9vtGZqPWPq0bUcN7vk6w2XMaeLOeZGy+aasjorW0S
0JPWHctqWY21v5yRelnZAYFtpGgZzubckqiM9E8af3jh4lMkYAcH4JFExKs486UU6Rr+bu7wdUjh
+Ydc5e/XHVTcrE8dyeb3TxRCU2t1tTJFwkCjLv3BQhYfCAzF/mhme3xbZRZinGB0HXdZtIj97/it
s/Hj69nfpqFR+tJdIpv4BwMAS6hBfMOvocec2Z5LfRnNpqs4yQvdwGONcRYXGZKIFd7LS2pI+de+
3omsY4ISy7wPxPsbSsRFOQluwzY6Uf/KWmKjABs1lgOHvVkFseEzzeRF5e/6HfzqMslW2LncxC4I
0Fsn90NTVcy1oj4X8Du+RNLWRSnmttPL0jAGqsZ0S/ZnZI2qolAjgZBcNZLSF7E/+JnEaW22DUHi
9PX3jBUVvMZtk61DugnbmYLZZ0/gixOdqEsprks9OeZsevAaaK3L/pDqLFNioRVxONF0LylKt27G
I/x8osl+eUKTy/EvSW3pjvJwRW24A/3PkxpDM/jYRqdIDI+34WY9LabLeFyN/nId+WkOd2/oPPDz
pvEE8lR8060LidEUuDSxJpPZ3uFoanrJ0DjwR6dJXWAlnoj7sZgaDMNro6juZSWMyYhmp7cR8zZR
PeIjQnmhOjTuo+N1jpWGGPN6hBPfE/uY95xXAUX6Knrwbw0MWOJiGFQaEb8qYPXSSHYaQo6HZC0v
ZXem2wmwI5kCQ0PL46+insdcdoBpSMYT/jLydgRSiRs3PsN2cInRNcf9rDGXCsKOH1dJA81P2BUa
NyUBOqlmHSugyzv6xTffxYkMfTKNbXSrQdg1IzQS8n6T0V/tuedc1df8lT6zDW07dBl7h3lFaiTr
PIWPBNGVOK4BDjF/8pQ/zUA7Tb9QmZXSUHnw1FXLueaYp2/Co7Xgy/YUo/axRnL2AFviHrdjFoEf
cqJfLgpg6aE1MLU/tgwpcF612B5Dby0iPJjPkX+17K3CEhjqNZjGAILT1REOgUqGLYSPEjHcV3pr
fq29/tBgeLjv2yzAnoWeFaTLke8HTX2FVV40g9nmJ0UJEdxTdhpNkpVCQEVV8ojOJbPZBNbGfwTE
CC/dMeMD853EPk+8GIOrWCuTj7VdeermTR1BvtT/HD2g8qJVEvYY9fXm/7CKLO3USSRhbnUAbxw8
ldvz7tLIxXlE7MDbDHql7/gkZGETywOtVpZ6pEoEmmuEdbnYtNdZ3iidchqH4vFrIJ7hIjAgUnPD
UEnuGSVDA6ugxjCKxFVHcQ7M3B+9kkJoepLvh/NYGJnIPcw7WRx5sEVX84EZOVA3Gb+kYWh83BmW
MqFmGiQE9kaZHLlwGZ2X8Eejik92htBh1xsl93viGM3XAGXx4fQBv5i6sDdCV9D+5DAF3E8Enj7P
oFDuWgYdlhGUX4j8zYc9Hd1IEI7D3mImv9IAA7I/CGGrJ+t8XNK3wHgg93J43qlCdKSPjFySJLfY
HOH5S9BF1R5+387vcmv9kr0iujosAQREjFhy9P605bBQKf4ESs4U4fJzVq3Q13foJ7VcUnwvc9zq
I8lzNkoORx76rfwcrRv+2ZDVuTzHE3Qv9biF+A4T8j71AfTklTFmJtJAFPRf1q+ZjMGpLUm2c+BZ
aiHeERx0uEHnvddxEdlybu0MWvG0avZherZqtDf0dYOv6yd8ZWf8cQ9TAStM191VkveTjck04trK
P13+5mZj8UcgqxHc1udSWehzltRa/R4omGU4z47TaPPNvclLNhueZGm4qBIZiTC6RV3sax+CfJxH
hsYuPF8h/lKS3LeN7ELIWnFM93k+dGqNaErSPz+0RD8Hg+fyUAhKa8Iyv1aGtrRhoBW2t9fkS+QN
rawi4Na2MkNVKWjqLjma2ztWTRCGfiUGBekYDX8xSotj1dRuQ4Gjir7lXZ1TUtjARKVM6OF0W1u+
nBBx0SJH1+MwTi/gFryaPg5UK+AS3HfLlg2T7L3HZ0ehVf2ADC8jbQa4x3NGxI0D7EkE7eEYPETD
0PUY6/dYCuMn59p8Hni7FYhEH+h89MX6RFrwJluIsRCk8UbJDP0UcPuArmAfRoleONIPsKuGemo3
TYBt+QW3qDyop/CDBWESYJiidSRFsDGeOdBWCwQXwT4mrJ3C8vqJjAakU3sJJwFlU1VctUnPsnr3
O16tRyzDm+2VKEKI2U4Y3SKzVRFa6FIy84ERbbtzb8Uw0LXlYhqI0Fc2bFSjoivaX7HMdJZ7GHsI
S3ImIYXXoN4bA+5r8dbD0AnMg44w6niy8t6UIYDnLksFQShBCkROm/utg1iKui7mFpA426Ilyz4J
rFNH+8kVS+CbOWbHx0yCZHKUbEPTWUYQDQ40dgnvrH6XhVV6s9Sjz7eMRmMxGupwhPpFEBta/Rml
Y0VAQ3+RQJ4AqecH8xvhVdOAudSd8HhKQyf3z4+/mu2yZTuKY1hn4mT/Hg4U7QXESvmBxPdZwLWY
jGmLQayCSvpa6C4tnORVTI960FW0RnkjRL1RtZB98kIU7d4fPUxCunQXERvkZ9q4NUjtghb48XO6
LdUNGMX5emYb8nV/8jlPIZpm6smGqtrqbPc9Wpyz9lG9H+QXFfgBX1Pz07419VlfObXzscRTHUmd
gI1lWVePfnZmWyVXfDyuy0K8x5p/3Sw9UiysAFjMNk8PfzEmkdwdrkkPe9rKUN5OFGj83IsPJd7p
ojMv6ZotB576jr68VwI9yuN10hlfVnLdOzaca2CQDMl0jvMA6ZHoeOi7y0End9k3jAKuxo3bxJ9T
wYxg3/8UYPOV32f//KZV+wTKaM9UUIYx+h1o4G3l+iiIJynr8534T2s/4j08v9rDNP3PtBt7Wnyg
hdxcEXkwHf2jk40fAvQwjaKA1wmQjww8V8dQcBuYalnxJ+Bl03sbzSoecuZ5++Verfgy4EKdTmLo
ZOSQciTli/04GA4Ie/nre1n6+gAQYkk4FsUFbGC4I83ZATM/VLAuh3rsweFRzYnIBwg53SDNWI6V
a+C0OnO7GIfBVm4lfmWrXfVd81V/BYrer4OXoWxatDOKSLvjB+IzURK19CsSyPZLXE37259UzN+y
BQga9LWF1NOkOEGlbZLVQ8mbqyYSil7Wha9AHZJHqlkBaK2vGd9FF/16v6omBwmWunvvL7fnC18B
qR8gI5W4Q7cG5JcuX4/M4026odXvUmxIU9iTaRN/mlzuMxi++LNimA15Af1L9F7j1opJuWqTJys2
j48NuuvJmqmQQZud5TUD/P3+J+pCBkxGFEVDrQoEiLSgyKAYBOafJ+KDj8kXLUSehvyW4AtiZzR+
zZDP3N67Ad8CNyb9eeKQY6jcg6v7C4+3niJzP8gmaBJkgmLblrRF027D49GcWjOwn+BVQwr/51+7
5v2OzvHD8Cws5w5MByOy9AzYHQs0caV9UF6MI3pkr+gpG2eYPwHQudns++KH2PcAtlbA64Egp5lC
f28T83RvaEFy0Xvw/+KQxhPaVCn7Bk+RsigIpIt/hGqbbAqkSAjkBnB+2etAnNaJr7qU9UlKIzeL
LU8UcQAL7JxNor/S9dT0enOudDU7zAE67Dizf7+ByvBy8y4nQZGr7xhuMQSCVmm6VW0kxx8ugVA9
85ru5l7EQAJe4+Qox1KJDlu2FHUN+ZHL5/tuyvhRlGDUeYSPOAOIwwCycacpWmI0dAbKZTeDsMhT
T1kLjpwubGkaSx4UDqY+5UUfGWPmK+eNSumiIO3VlhHtKC0UOPwSmhcRoiG1pkWLZ8vHhjTg3Bce
rZtvD0GOvktTNLnd4fWPQD1P1eWnin2tzajZLlD2orQI+pyjWEDtWV3d0Uajm5GoUUAWtGEEUuuG
9z63G8SVjdb0FX1ykDGqcdLJbb3sG1Q1YlM2ghL5bM2GhzTnl0rirmPmcHsW+GQeXUZ/e4jLUitE
IezitWSbpYDRrVihoKb/Fsj+UNeT9gBTbvD2XuwPd9NiXgweZwRFOX1U897CoxoyEiWxmJWHxV3L
RwPhMoNBH2lNP6uZF0ABncpHJ4SrMKOogiM1v5958DfQtqFetGdQcB2/0cx6SLdFG6jBkJ6ZWcID
DCWiVDHVdlFZXpH+bm7cZg0bUv2QJBCHZheYRTMZcBuBsUUwGVuPy5z1mPfyYTEG188WK5hPQlVM
3ZaxBB6wk00kYBQOQaaekuEvLg7z74gtNaaJqJgSKv6BgvZY169bXr1rX/zkaZwg8OAk2HEjBZXJ
tm3EslJ9+b1B+oPdf4ChxNOtFxOzd16LQzTonv595iM4Uwvr8SbcrB9TGdsUgB3ke6JKQth4rcsd
bLms+T6AjZubm00nIaaFv1kw4xLVzLrjQSAFM8pD3ZwohE1zuC/a0zjKZhMUvt7y6CqFF6+F5Lt3
9R9pJhP0PJPu1BQp+XTtuXipJfakBq/eLquzFUYuixqLIxWMTHSwYaCUSSh/s6UXChozjjnGpb0X
7bdMdhT5VU1pPs3/XatVMPKt0hb0jcMiZjapaCI4ljwd3jftJtSyYe1UVrR5pHbKr+ujDsyb3YNZ
aacuDdBYIGy+s9+3G2aT4LOlfGfcIRKt9936368+JldAIl2t02ne0YOjgeGZgTywj+P5r95+PFGx
1GSszHspMkeq4Yv2BeP03F3BvF5IEV92MGjE88aeyDZEqx9TZdHFzyvRBGFT5HdcAz7xWRGWO36n
WhiR0yBiOQj/UKoPAs71k4ogb1neGnUaZnuez9sN1SafjQQgop+eKFu/ZNN2JKBkJF6BtTUtjjHm
RhfUeMilDlNejRJFjkzUHnk1kWcU6MSRaBy24WU4BpHW4mTz4Sv644hKhphKFF8FEcaxU7Ss0NKq
+pOTXXlz9j9Q6lwVI49XWDav545WC9vulB94C1pfQVVIVyZs8aQvoR8MIWl7ASi/GM31twEyo5fB
P+siIihk7QdIyoeJw7IHB+cRi7GaDHUKNNCsrIekf0/dyjhq4XOg1GiGCSlSCr9hU3pRNHDTtbFW
3EkR7/QPIuUX6Z1YnvimYOVESFnAaHtitWuOs8HSgs7QjZEZ00PPGbT8DGW/OAAes6dKeiq6zH3X
Uah0dheozmq4be0os17rB6Sm33JaHEERFsljVqDHNPn4L1sFf335E5iNYLYJQ6KaWuanZ3r9dwVN
d1ZIyoDhaDu1PzqW/vIwR8Teo/xjv0GiMTYgYdoYhy2pfYfgtxSW4g//KwYUMFsKye+4lLgKFmOV
vi0eU1ERWpD5ByZ33sUp+MQp3XbFaWalk/MIzEaShYUIyEUPQibBBkv9tgevmcnYHMCBF3wU52su
NEm1LH3eD+sExOtTtOn2rd+pq4R4Fovk+oveyLwQE9U/XaFqcniSz/pHzyCZ0aTE7+ocGr9PDrz/
p1CAbrcsaEun4CROwImsPGl8SRP5Alq9n85z7teZM2plMeEuAlv856QKL8UZEcHOw35zkYdIldwp
D9/cen0Ctx2qRzFe1xNLZdsEPTEpWMj32IsiUz54bC9vPm3MMo12pVLzQd1GfiLDhf7UhdxInsFD
ku7dBm3B+g9nNQVp/CY61rLhCpL+9C30/RCWxzE/nFYnVyhyD7B4r7xGTkySBYuCotGGOFtVbDAC
a8f6+5Yh10LCcZ5y8U/mTNFvHB9Sgn74AW1Q7fJzfvOv0E+2bZ3JcI8fz3Oz+0XuW8xJVz+4fqTs
elRVYX4TYdrtaw+tzm2M1zmeufByXusjyq7LjlKZAKgWZwG/Gwutp9OThLeQLmubkyIwq+rx/hGi
tzv5uax7yYwyqbrzNrUBeMQ7wO/tWwPPrlfZJzAQj6+N2xLGI6EzzgoijcrDLookfpDGG66y10KU
kb7f1kkVePL1MJ7nZAM82ckUhiISlacNZ8XrHtmZQZDuKj4RA3sPJhsTdi47kd1sqc2oUn+TlnDe
RtTEmmv/swMO2ehJ8PxBwiaL6e3svnma7/KROLE+oukeP+gLJG5Tlw2ONLAu2JO9bY3bAPENXY12
MKt12H5rVPiyhu+wifANT8mwgDOkgrhicWSd6R6wKIQuOk4C+3LNrrPFU6PKWDXMXxGnWJtQ0WMB
VMLsnj6lhjBsCDD33GkmXTUC3TM3icrKStSsA/4WM/wm9sJA5OIONkRqPeg9xs35F8NyfcLZEDNC
SkC44foK2/bF1JlZlLR6lMqim4HTlSDsk2SN7WXHr3KogN8YBSPg7nEhyjUYGrjUkOtwayCEgXWd
aPyB1b3HG8v83mKX/FMuzVR77074HTq0td0sK/8V7WmcZtssBV2uwtuzjDBNwOBxPUDhNLlzvNjf
/TXy1R0lMoipFIVMrPgTpp/E3w/GPDi4Clkb67TAdDK4BnsbCwgP5oCVViJzKpzhmBC8p1bxy6Zb
8yZqC/tRpcAMRFaDOXvBAi+q5KTJjeaYy5z+FdgBHIil2v0aWjH0pTb960LrwXoothtUqpQ96ysI
3TsWXwXcIHs+obKfTVQW8uwhMBeETOtuef1ayUtiIaZjWRUF+Op581JpShkh+IqJO/i7vVH7jq/R
iSS3PmGYvXJTGtESizSF52H2x3TSNoxxBI6mTWokXwNxuUixJE6bh5PzxSY/m5lU70d1GJJOpNAW
sKCVwMi6fX0LmXCFvPdi24zsajGri728ndsCy8WiNFQD1BwHQ2ClfO7P2QqmhDljRW+Fa2JEGD6f
Wk3b+knZgUoHt7OD+gNFFMdKzumTJ7Z/htD7nBierImw/sUqT4UAldWno5Rm7iGs56xHh6oWR9Cd
fHDPkireWXlTq12532Y80eNEy4/0eSv9ndmr1btwxPgyzQ4xfTgO5hrEb94rGp/k/xQNAH8sNmt7
L/3lMAKu7ffTILYVOw4ZtiQQn1ZscXS93wbjCVvzsFJEKf2zQVnnQGvuMjnC8K9BuAC7RqjT9vX8
QndDcuTa2/j53pudmVLnTDVnIzYaUrZm0/ZaVuQObB8oMPb5U2Wse1w7pKeST2m0a1L9zVL3AbNJ
27Yvcy5qHTtN3ZU4m7l1F17F/RUttFPK2qgTf8nUZ/SO+ppDL2oTHNb/oICb98jjnc17oKzboKPF
QufxrIxnPs5odMgc20mEjGJAdaXOkx388Xvi4iC51r6sA5LeKFVuUW9XNh6eUxntgjQgpF4xtvQg
QUE/qEi0JUC0wrB+ByxOyoTMqY8tWWsRNVSDiewHt+TdF4zBV2moinqXOMs9zFW3ZB1m2x3qfOe8
fFiTWnMqExB2V7xu/ox/aAbW5dHf4UgktD+PV1XmY+NbOuK4uEZk4B83FdIeTSt1VB0/An1wYLQA
eSzZ+5kQf3hj8Py3W8oGF4Oc832TROOfGJSLeiYbNHKavE43aREcqJ0DWOMo1cIkVyUJCvINw/X6
ZSGRXqxOXDYfE6yMhUc2QY330hwztdro1h3cOzyiV56D/r4RIsxmn6IhrNqc150kr2z04qCG0nX0
hOAxZgehnHa3zX7v8bTdiXNdndBXQF2YlLu4RMv8X+KuB4e91ETIMCB/Itp5uM8DEOp8x36fJrPt
CH6NxiRnasjdQaUj9CJh0mDLFjliQtYI+XA4IbyI4eJxZAxRHjVJCWuO49pd1r8ZJk+Xr6fcFdRf
lVFJj1SCaTKR80srQ9SeqeZ/S9s8ORMrSkCe7bpKKA0BI/waFdDn5IZN0SR/iZi9hviza2hITZNx
zW6RhS6GgwhHeOY+VCsCedNTDacdE1S0PLeNCvHZtQIK18+n9NLcTloE07A8TZO43BLzdyIB6iu7
W8I5GnDmSA+O9P7+UFjL+MeDeDscASDdCpBkG03/6YKAMAiUypNogizXt6e4C0qgw2AnNG9wYV73
BmmECRnqNbySoAum3s1iJKj++xFIiv9jOmCJT8H2SX2HJVC8AQ2YaRhJl08jAUjJtKy4DtKLden0
hnnPlL27fnLJ+IaqQhDDYxas5OeA1cfi0CNBqTb+ke9gmjuLsy8AnRRAuxbFAcZ+8eg4GTBL1MGd
pO2UtUaDC1p4HhlEBV/GSs1Aa39nPFa+LSZfWYbvE6rAM4lbo2wnu6D/+pdFiifWz9kO0i2RMmV5
lnuoY18SLow/uGaAVBh6BjkqqKjP29PgxdzZoYQi8AgU8rWdqXJp7d7AT28cq0z+1EpH/PZ3qO++
aOVeA00UiOQ9w+2rupOsx9BryTRzcfe1oHCynSM6063q9VlMIfcj7aBtdjTMRgJHFFNSznhK2dxc
Fp6ObVcPqE4LU5k1kZ+BYAYsQFVdL8OuGefUDnby3LUgnwfjAy8SEbpk4Ewb+2aNsHN20uOS3T5v
b0BtwZkQbMTA96gA6mGFpmjF4zHkRiXUS8GtnKkU8YgxTB8CnUw+oqSRNtWR9TlboLzAkoFCY17L
wDYSBO9rCE5PoCWJIUQde9DoQa8rPa8PgQebsGw8iAjJ7yyfhANRFwl6rQArws34CUQYxbhIAXs6
7H2gMy5Kl9cOnAMrVOCbwTqRttsDLpfmULLxGfLcBaSl5vxLNElproHf3koKmbSVTgnlZFPwpegn
IxIqMh6LgwG/EQ8VTooRxjZbvGYhK3C4xUFL0lZK3tUdsW+bn5HpYT9WufwEGjoD4VYTdKBBFI/Y
Pa6c1f4pCnz2zxtiJGrWwbsiS3ApqfreuMavcTYBTbvAMNvnWBU4AhS6lxnQQ3S2FBYO6IW2vnGE
O4bv72/Sc4ohjWVEsvn5b6FBbyl5ozQoBkoe5RbY41oGsAxd5r32vPkxNdU2h/GB0gGpp2y9PRuF
6gUASzn5bFBhhoSJQnswumoy9LlWK1kniLjnx++C0R5KbxayZfAWbdx6XOO1TEpH68a3Xerq3aIE
seeKmMiVaO/7kHDsLxP3u5UbJcNSsCRBXuwhtNwWHTRFF4sgzU2HnzuVvXbzPvuxqzhtaqUhhgBy
z0gi2y0zV5zx+0BcDs50EP6Yt2Gdou86njkFuv3E/F7OOnF/5tbArkYJ1x8hawghDFOSNOAsXo3R
Hl6shBvgMjm/jZgyJFDnTztqv0cw4+95VQXxngzw2LQjUpOLEIX/+TzmKKsYItbfYjtZWd0vq89w
aH5uHwwPnoY65AJ4SQ1vt4Cj2WY2zVI8tNExrnCovBQ5R4N/F65JnIn0UavV+7LjLg6AAfDyhzUQ
wm1VvbCq+/no+CdYYMuj5j4AnDwiSOLKa7on30B5ALvCDNqm7/LFvTIsCqedbKDutulWqbNbwusQ
pIb+WEB4ZaVeCf2nhvHz8xZ7PUlW5CYtwSA5TRCA4brG1X3Xcxm4Mh86wlsgUwxqOmAyqQbnmMe+
DMFqJCfSBJ4XmuGbV3GkefZDAAu0tKE1hVvBTgDQqnBaLmbT/MudsQtQ0eSMM6YwJ7yJEAZhYCdk
KfEqc1rEDg3JIf869LNKJv4LGKrfKlfjWApt08lAGDk5PxJvdti0dDJ1Fbnm4rTixYdpEyC1eUkC
vQRzuNh8vhirwOUhjsj8kJki2WN89SCECQH+aPybt9A6hLesGNZ0qoCAGsvZg5yKzfQ+MBuUuCqo
u/QQ51FN9eAkizC5tel+WQ8CkSjSVUVNfwb5o7Cq39ySvl2qWUSXd2gADlLm2mur68W4+L3yB/cA
9tHMWedyK3fA2cJtgPpBoL+9rAZS+Le9C9I+hVW47ErOWQ4WH9q+HzCVbteBlnaN/44wDdJnERAi
v3RB8eyxqY2W8g7oQHygw90e1Rl1NHF7YnZWuC4cQa6WSlolFP98byX3iqv+daamIv4j8Pm7wKuY
jog/z2AR4jy8t7iMctv1uzMXkmtCQEhTia+Tdf8EVnJfcPIOPEQJd9ENvKyfFR8BFxrn324yE6hm
ADgxSnh/ujD+nyAij7YyW4M6n21x+TPi2Stn5ufZ+8RJ5xG1AIoD4FUvnqto/mmu1UBi5kR1tIYT
UftGP6QzteXIEh7n/UMQGW9dx8lKcuwx5VwDdc0v3Spr/bRw+HHCuiI9HK4jc0UEfrFCcQbfmIi7
D+ggttcjtvjOlZR8EwPXK/6ZI6czumXDNHCRw26NBjoiRWChSbYoTslLXp6G4N9w6W1IvIKqeuPz
XETMt9BQJRp/goKlsccWEKo21qVVogBxKCFvMMv5bkOdejqRdpp72TD9pNBKSB/Z94S6VS6Oz6Dz
r0MRM1cqpT+KaXLqaU6edTZ37HNxS5S7wiwjCf/IyaMltOsd9CMDYHrp4ENxNvKKSOJ4pBo+nWyi
0mfIDd55VWdCm/qerIz/o26aifOpOANillWY0lrHnOpVkXdO/G5Aowi0NHbDsf4FSlFEdT/un6q3
SRTOFq0Mo37c4HVin0/+GMSIxBDqKnGcKJkvIWMkUPD+UClRToAi6r+jYRC3GdWJS0/XINlpDYYw
cnQpVHBIPEgDK1bRc86Oocx5GOKLtgzOaQBfkBR9l9Y08SWnYBsLQ6D/mTkfXR/dXcZFmF6N+vaj
LNYo4B32C3R3xHG+rbpeNA7WLDinH5pZOsfcMIKqKJKiRRR6PRXYqutN/C4ytwu72hHrvCEi9B6A
/hsxGrbUMr5O+gkAaswxBDSggPmdo5tB8cwtZ1agu1rryISptqJ21HMIwyAckC93uIAEh4D58mob
JEwKzLpdbXWbdZV/YmO2DmfA7RDVvp0IVWWHkYxbtMJ1rVq23U0HlqYnxzqrMD7d3mORtWCEtvlV
GaF3q5Kxj1YLz5Gwi2x8MYFEQBl6W8YDMjrEw7ljE+eh8KwzQWsPdVFlgYOquj3akdA++vjr0CoL
u3iNkIdINrIz7R5B76wxByhTfrp65Ql+G4xMssddm59RFjWQQQd8WjCLgWmMjHT+u2+L6KG5PAVm
aFajoemHV8+YA+BGyv7B0p6VX2fnD2haQkc13Ps9PHzSqJpgmIAim0XEtPhdZfG45KehkinX0JuF
Ng73lJLXZKmy+qZxqcraMXcJf5XcqSb2QrCNvmB2gJX6U92NON3hVpud9/Sy/37I4we4seSENZE3
CfxrnsL11tbYXJPF/GU2xFHhORFIzgOymPhcmgsADTD6X7DhJrwa4PKiD0X+mhNg9PTfCDNGbaHe
2iCU54fcPF+gT06vzLdGB006OZgrvNujeWKuz3O0wJlqGFfEqvk8uF1iB3WNEUvdqqmMEUoum7mb
Jy9GK1kZSSVjVaGr8nhHds7V6hjszz7oyLKWahMSaI90F9K4qmt7R/vFytnSaGpBkGi1wDP8bkYL
D8Eky1yrtMcTrf6CCOn1mXzrEuzCgPVGQP08Zyy64VCZPM3VHyNn9iG9QrEK5n1oARVZ85zQkGj4
IuIsbsYGfag9W1X+MMqO4pfrO5Dw67c0LTZrHbNuk18gcVLzlpOQtjfUQlKSPIdonmA1e09FBwEi
Xyrhsl+2gIuf1J02PPSvMn+D3G7F2IYbVzaGcfyrkQ142WovF1N2MVeOSr+JDig613KxRIHlUi0f
0K9DIlQ/I8cTCbUPzHdv0MHdFJ5s8749kapJ6MFlWI9hycQt0hyNISO+A380CXLP552qAPQt3xma
//8js09H0kdNJhl+sqONSLllOU+fDwaqagF7PikZPHiv5bv6D6WMQ0bHzjNsWkA1fkMiVySAe1rw
+y9Jamucn8OYFJzvTo/qkAAAzyfNfvMbIRE3ss5rI3Hoiq7zBDbUVFZT1uLoP6AQUVfE4UoX+T1o
M5YSGHv2fCoY5C4tHaBoSEQWB07gOru2ulMe9o2J1mxz/yjuXq+DTn5xLb+81RFMbed40vfU2vK4
ANy23VCe+vbQQ9QLF5UP6duYCltyIpV4zd42us+vbdbBpT6UZ2bsX2peKG2B1tM8VG/3RDKomyMN
W8Jf/f6OJsMdeGMbb9fiDlwT4KH9aaoM2fNbBd6dszATBd8Qb9mc4jhfiSzOiYFG1zyONJw6VO/9
SPH8910wlWAksJcRlxaZrfn1YX0lV+YULfEDph7wRMybBZLLUqbGPqkU/xm+LNN+gXiY8D8Mb42f
tdHkjYIKgmpjoY1WbnSaCU0O9mfq0gZ/IOrnNkZeFfw18dHj67iS+jPfoUvSTu34E1MfNtj9HYHy
1clsJJdH37sPwjyomR+yyjw8ase0nyIRI8jOkuKdszB13euP+3CK2Gfgb6JXBuafr1w53aZ6huHw
mrrwc3rXSB8XwXiKG8el55M7sPsZkH0OkECfTt8XKyA+sNnvY9ZiSh4mk/5r0Rb1UxhZjUuVaez5
PMCLjji32cLo0Vn+/WAhTxWN+sQ2D8+lmU7kXvamp1RcX45jql7UAunE4h42IFucREiDo8dHjFgR
2EPC/CKjwBSHQiY/eMeBkayMVbSWjhIKgdNfS08G73CKUxNOreisbmF4Xi56YPNNp8MvrceWHMbl
EAnz2M+g/WeMBAMr41rIp3SQv8e+uwXtCsCq/qcxxv2H9JFlizRGZl12oS3dcCSAX7j36ji1QVFM
zVlgsEwtcplHNVKSP4FFkJlwUeCEAI6jVSHYTLtBP/EfYVv2ixcLn9tXsR5D6lUgAJ5u6Zlk8kZq
GXLiChaUy2UDX3nGTEXgCB78u5pNjpyM5DWQ684a78x143QV+llY3S4BVfPxbN4qcyHj5qw1dZIb
JTlZTryepG67f2l0u4bhrFZ2+hH9PbA3nLNvxIe0ZpiRbluT515zsozJtkgPvJ+Badm7cFmvWcR+
VWtdlNOXGYUqQd389BWdCRXASstWohpBRSs9GQdOKO0HyYxlPraLw7mAtPJQhDL1oUzGRYUkPYFV
7d/n6YqEG59fWt4gHqyIHeO2LLLF+ZN17AcnOFrQlejHvyGzJxncL3ig6NgG03rVOKB4uz/UB2Na
jVQuRVebHN2zX7s7U2dZBCCS6HIDL6gDYWha6qKyaFyI7z6O91FnkvdAp9V/+Z78LAyqxITPqbSG
74zg4BgRY5/it478iQQz7SaA3PXy9Z8Xoi+v+v7//U2UqMNkcNX1hGKIiMAMFvRla6VPcEAsI119
jJwdTNn2xEgxQUbn3S0hteDczjdnkVr4wvDzNcHwIbJHuFW3a/+ASrKjE2FNZ63JNVqCUP2RFyxU
1ghgDGCB983qgo5a7NiYKUrJk+dK5MDO4lnreGYJLnuV671pqkQJrIFa1GAz5sIMF+EsQJO6Aojo
2T43zeVLHJwwoJjdnI7XtNGMoI5w8VkCwSqvsxamsNQ066RTG81PTYk0zZobkL/6d0J1YVpAs20x
uNAOPA4M+x01M/2duJKmPLNhXF3JPIttKkkrCvlGIcUmRhqUyIZbV+H/g8RwyZaEexj1QpadW9Kh
dQ8cJ+Zxr7kQ0oSzmCwzNd7m3JFEM5QySLGObzCroaMybt4wqcvOGEvk7w2ZUUrXKMzu9rKOf+gu
WjuJ83GuV2fu1lZ+/D6JlRWkGX4y9Ib08VMXa02UByXEq08URCest/DUn/ANY/zcdR0LmsKE/rmo
7lBmL0gefhOVQR/yRjyGk/h1J2IepQkqzizHU5Wnp0i4hIBRC9yRMejAR9lIFQqS2BgcOi5mn0d6
OPANYD2R+l7XWVua85go69lYB/mIxwbzh2LenLyMxQ676pvwvkzZzW1cgw4rpNpNXT+gk1og/Bi/
WqU0TPqUbd+uh34AsqqRBhhjGP4qkcGel0FdXR/uzA0daMZt8g2aTGM2e5PAZwvMq3+g6hA2EAk9
hwUSz2rkFF9eYv83QnevXDKS5in9LCgNbPqeXqcBCh5hR+qMcUKsJG0YFfMhT8jd3H7xZf/Sfkkc
xsl0NcRskhjVtJfHKckLCM4rBbuO8UjN6PffWEPFYSvkstV7QUu2h1uzLbXdidptm6dUJu9I4uFm
yzqRufwkE92v1cEDuvOe0hUJKNTJRZujI+r7nni9uVWoFPKpehIE5bhTaZHYgFGNduWSSK2Y1Ffp
kdu0xVd/X+dZifew6ifvRjz4HBsbbx2vpE2xf72fDntfWXzQlHNb5QsmOK7xLq+SFbwXvG/Dp6hN
uuCMrjMznUwSGCf74DFnLtOQmxTylFdwGpq6YjIVTEwvg/idH4TV0g4Gg3o4BfHYw5NCEf5WwGPP
JkMyRVV5VzLCIG0vek8gJYt3rruW2I/OFtQieo8X+oe8hND6xKvbQYMaLEG637Ahj3J1Gq/0Cjkv
d6uotQUhXuYtljXrF8Y0HhCzNzVonTpcfuHwBWSMCUqNIib+NFxEGIHoa6aS/XIa7QSXPBIizmYP
s/vqOpsHVPd4PA9iucWxRbaYGDAaFzbnb1ZTLOlCXJEvmplWsmLnT2kW4odFSes2y4GHqvMFsEOV
Gwlc1k3oNZiI6C9WimLL7tIMcsBbzPCvSVSkrDFnzOy3okyHTkGcVdNlUpXS5Kvg9FQ9rDd/FDU3
5UmPFE6ZdfGHOc6p+Vdhupq3fgQA+FtqgVBondH4jF5bzvbgHveIoLIe6v2/c5EWt1gHAa+JrRe8
W5DSpLxdWWm9coD7Wza8MtYmrrL7JxGuZFV/2ZsbAGtgEiJu0w+50v9wa76TXaJCHQ+XvyhEdH3z
XiH3R3VSXukF1YVdq56ZV95djDQHg2sdGWuGcV5cZBsc83Mnfu71/BkFFTTp/KFzxtc0GY6KWJzu
2p19NQ2684CLlVUl2f/kI9ZFIhbBJYh0FsqcKFYxf04T1CdAHbP831Rteac0DKiX0ZP0HwMsErLC
wopExMIxiO94xB5rJ+rLev/0uAMw2fK7ORN9jz+5uuphUHjTIZJkJHtgPRMMadsDo20Sc7mdW0Iq
vpkU6McjurRh9se8TudQJI6Cy4kR8lXkAnyoB/wJXBJsq2uAa1fQbJEwXX+p6AxOSFcmzA6yWj44
o5PFmgA82zxedziu11oOED+VR+0C8AORr2EzD/0GW3JNQTztOYJTdjkhG2tVFv+nglZy0eShZRGW
Ds09hIZtX7SlQPj5c2MFy+51VZ9GwBPCszcuAHhz0F1v3E8FhIYwX/GBjlHrkW4T/RtWyQ1WYgpe
wO7GsmH6p9buMAl0mtkC+wjPIzvWVOVP0i7mxxCQ+kGvKGrN0Vq7QfxPfe7ss6KgHIg6vmgx0cq3
uCWtEjNB54MNmKgn45SEGVd78stzt/S8P2K3xfW0VuJbMMB/P4TnWkJyyuBEBCdj0ztl88Cl8q//
tt7D/JSw+a+G5szB+H8yG9X2yuapEiGLsKGPEeRNwq6d4Q+YEvK9q1Al7IPfNaS/6HTXbYCd5vPb
5TdBTvqbg/zOtNJr4l+1J5L/6IE0pu4eASjbww8Vb/YTz6xMNKF+pEb1Vu4HQ5BMb2Dk17/7DwJs
J4N4YRRYefIdxX1RsglNV8fJpAtSlyINYwr7RTdvjlpP6ztBleMA+lkusUNzhcgLBd4+KPSaqLtw
UuXVV5yPt9ezzyl1CQP0IU/xepCuNfByBztuwrqjkdTWrKbNCayinpuAlWK2nvI9HiaylxUPO3Ue
ph3/WTtHsuQYkfQFrWEuDdY6pApxg/fc+JINRi6mrR9UE7EKdYvO1x8i3LX/x4kCGyF4JuT25D4t
R/S3SG17aUV052/X+ZDpWOFNCGE3T7pYTrz96mOGOLZhv0fAa5WP5PPeFqFHAxgRoKqRVxaTqh71
30SW4OgJVh1PK+CSWdhpqAfWqkb8CEpd4lW4k9XQBi4zcneBtHimK0BjMq8VJJDp4nkWTsbiSiby
foHy/mOjEL59A5WyVo0Qc04bydg2DMoVrIW3we+XHBxcniIx8Xjzs4CwM4NHelCdsdj2dOof/65A
RcuK9r/hLyQ6T63w5/gLb3YktFML6V1MRE7F4o1E5N4Qllqg5araom3wfhJu6LDcrDYnFyuEgEG4
F70ZHIA8cFs1ApOan67TawaeumxJSis/n0g58+1vsFNbCzkHSYeG2UZR1rZT5sqHwURvFmNOFUyN
sFs+rsdnMw2yjJO3G3DTvmajBxTjWectiq+XUxH03/pX/bqGF0NUk0MzYp4TCLcs8OS/BYxCHbl0
hQUV5npipkR5fa70UOU3jEpabRVu9THxa2g9PgxcT60n6N12+Uir0RNqaM2fDLNGREEAEkASFZl4
SkXHPn2OfpN4lkbbfDbDMoLmr2DkscN38ibYvTRpikD7G11OR1Vt5H4KyAZSeXqqqKFRev2nEopd
/StNg7W8oK2cq8+t320T/QZf0OIAIG1OkBnQezx7mrTLQQrgeYP9S8Y8wJsKAlOZLDTtEda9THhQ
rOhgRUC4vVD61Th23rcVILosdvypvQjAmAWj+CpRh1J1NOF4jTbvET2bIE5YA/LD14GDn7fIlGlK
yP3ZMlfHqhdqxtexZBRh6Dvh05HEkv010WUeOCfXBgxZauzsmMqcBebTFl2uteXsUFkDxobbtslI
rgAdnhUn3Q1ieW/kIMmz3fbB5HdG55xRabNDn3qJdDuZeWinz4Ckbdg7KXpHOlMBN4SXLDIRRktq
ueT1vCR2lLrGLdePNmqVTzX0JWFMCPjA/Ar26aHjO36Clv06nTmaX+WFBAnfkaPeACCwwoEQPR4c
H9yYRHfrfk3NRsI1q8loj55NKzS+tAYl43SrnRruujb8ixUxUzdZlsE2POG/IgVPfaJSJeSejAds
rXZi44Id78VHJTadbmDy7gYwgEcnJ220ma+Tpl63Pr+YY/6HnhmqQieevJKbnuFF1zyFErYv6qJy
z69sOzoYKtl++8Im7QpaUaP9Jey+uhXzsb8PHz4Mv6sdxyWWaqDDuMgwfeVPy0izFNhFHxl4NWg9
nuz6i+dTRp8IOrY5EdP7vX+sb9i22h6rwWKbCYZIdIp/aHPKtWj2/FPLxhOl+sGqVdD5iOhF7BI8
PdIniXgba6kfwxuuqBkGf1U7spiw5hKAm134gpQH0RTDdUImfBK2vsK+7cEKkQ1J+C28YdI72BAD
33xrKxwOLXg/h7bpMNoLxFYBkS3JG6uteQbKDVRS9ndqbypuUn+H67QeFL6sezWRgD3DqEtftdGh
PtD2sv5NuFZFQ5NnF6WuWe8JUjVPRcWHH1izWQHc+hwMfCl4CQp/4j7IrBVHNddB/Gz5oYytKyDE
mFh8lgtQrmYuY+WuMrlavarGOYfG5Ei/EqgUVo2rfZJo2xoSz+LAul6wW/vBRky0US77MprDJfjJ
mna5S7kDYYfSssBGCa2yEp7qdYOgRfybWC96FfCXJBGiy3B7VXAt4YsjE0vNML9l9E7vGN1dKOJU
oZH/NJu03KpBjRryB3qUHlxPbXpcYYO4VNPmjl+S7B76mpnKV/LV+OS2/qB5/m6oki0/3tS8M05J
0H7sALqGj+P5gWE86sWUEf43SC/y6kvtmttLRhsBGDvJ6CEjuh7mUvchbQq5s6YSc1+/NutyPyK5
xZ8LuxK0NCZuXpGtJkkhRqf7xMaiEMFmV+fQIDSK/+AzY/uhbDGsLRFs6xkjI6TUsSuEQf/OdSwX
x3Qn4pI+UxlJDI/lEaFSxZ9nmfN4VWJDvKToiPW0+9b+Xb9q1ZLCDPBu+3OtS4CBmbx2ppXTJI1X
OoEXk4FOIOb6KhnpKLvRaAmAGanddEvxRVYxT7QMKUJsfdvWxY08poPdlxPSgfD0AgSHLxLMup7y
mxSD/uzZtyjyZbJcC+ZXx6khzNG1xGrv6O1BomBM99gX66LFS8ZqYch9CeNR44DxkNnSZmAgkaaY
v5ypgbN63cRk4IpfZXWnqqT1w6Ey6NWSmzyZo4g3qSCfC6edm3foe471ck/mPrXingddv0AEmdhA
riOm1Oe4BCRJsEFGqbulYBa45BV2eYNCcPYx1c6LpDa6jhqxAshw4IAXdMdS0KNi+r5S2rbPWikr
uoa0Sy4nlyqsZ1OK+G5RmaEZhH0980DmQfFeLBfq4SBNEUlxUOrfKvHyTjmfNqY65fmMYVdwN2+W
L7zSM2+XuOyFCDUHDR7sFis2PcELZvq5oI3V83r/6dCSi/BP+eYuqu27YPZv/iAvNr4mFfjgoIGW
/ItTtImLnZXPvyoaCCGrVBTJxMYHcRY+BGJ2r0TWTZm8p2GhnMxhYb1APKF/tVvwLpiF+U3K4u3O
IsyPzTO/zOvjVOHDqFR1lSmjnVb9HO2xK6Jl66ns4vkuaH3VzL4Ed7HUjGArfs7K1/zVLHmZsLud
4y0ghOjL9a8EzsykE9RqJl01cOyjD0vdW4lHIXCB780C5vdWXFxKxKPdMCLPT10ehDhtr9CYPJqM
uhWaOrbParBMi17C/5hHhsmSmMD1XtbBoQPFZ0LzL4QkgvEe5L+GdO4UCGgwCwNQp5/tc00oMRgk
LfmGVPII/5PiOcomSOa6dEWvzqJwX7OrrV3ZQBheEmqEUVJlkLbF2TCVENN42Gdru5pfMeQb00e7
e1cnPczCt5J4xUevBAiwwdti8OM3kWOTxzOGfRr/bcXwdnT8FKHpeE+9AZVe7OIWE1RwRDpRRa1z
8E7bYLTeaz2hmQ4TzBJODnfNRpMiLJG3/14Pc9eI/aLhYRYiKoyhYCJ4i3Legp9woOV7XD3Rh4SQ
pw8RRPeBielu4OS3VRasEEQvYxXie9g6BeZV+VhB7Z4vlPiS62pF7t6LLXEHivzOoAP5vThA+kcK
KM+WHLximdl5fvnEQqOjAJYiDa6/H2mIqp/JwAbCMD5aEu+4EERzT6p463M8ilcu5WaSFx2q8fG2
iKHZT0RJiOJDxTDpxasgASK04KCv+l7Q/TSH0cC7vcOdaQImfSefoKiQwkqFEWsrIGkos6wp27a7
uIGnQX3LRFhMlS4+CyaPnE1wgWiz/nLJ7Uj+iZzVJ8Ofd4X08L4a9pieRKl+hNfzWweAzwUayjci
5kRivxDfC5/fTKSHTFjrGyLfgREiXKynw+RbDzusItuuKcQLHfl28FdOaHA6L0NaRvf3xYoy8nkv
QoWjvrTr5BSdc8Aw2ifb9IFqjFBUg250A9+ENkO+tabkPzjEmQD9q2u9gnRUWG7aTkze8pSUTAqA
eW/PoxO+e0/E0DyOsKQ1g0MYeXOSq3yXIIQkh6ZhsJKlcAhrTVzAr4tqXFUFybXG0NWsaYdhASTf
rsHOYB/iENGquPH5yE0kz9PcPcsCOkkMXfboD0hsl6my4zcL8fbhhFhM7Dn4/rdgFeeOJhIlnYNY
fnzTSsDVKfoz5YXzU5SG6Y+JCokvd+8Bq/yp5kS9RLCJlEFfwsUftGMX2BuwCUA8Hojh9dP4JVrh
DZXc4sdcolY5RgSw52OayA1Z4k0guQUW5QFTlKb4DT0RfSNGob/4j7r7o5uWk0iZBx9vE3O2I/tA
Vqz/prpIE/14pFrweOt5t33Hrw4oDi9j3hTDsi66UfnS1+vmepwDIOUbBsKyJV3E1bxyJIHNOmL2
WovVHrhjfRNXjmN787kXG/U+EPaDL+TGbDyhJJn1deWPOLj8ML42xTHocftt2lVYSSRFi+TyYn/K
75+Kxi+grbDga8rPIYrEkDWILGmFGPJoBAhtxyZpQdXHebuo4b859FEJjDPvdO0/4JDs0cGhqtZX
h974k7anJHnkxVa78sNX+Q0hPRF5Vfg43p3UcOQtqLCw71sT5QonxwA59FMEHAjoxiWZw0UDt15T
3551ggKIZ2EoGs9sjFUyb8MMObtSEK8/Y8zwaBa31C3OS4iuyvgKxn7xm9w7lXZojVl036eIpMCv
zggeNI0qHqcpQgsWPzAbKWJFGC3Lu44nKtNcG44Fn5pMaIVoDYNojjAmHCQKn55b1Iz3D6CfywWl
G9i1rvJAfVZyLkGRE9ZQuOmjQxgvBb4TPqqNknBm0YjWYlwl/QvIPBjCj4ze+Pe3u6FiA70T/eYu
dWB03b9uV3yq4CEl8v1OQgqwmjj0gcvzQkYGnY7FHqfXVYt8/kPlpIyNNY+TwBPqJZbXGby1fF3n
IwgLlfbJJcCk9IPlvA+AzsjnYd1a4dpiaHBOEmChbCE0HigrjxW1OIZG7bYr3ZbMmbZ79poEyxyh
BVTetAzFwHh4mpJkEQrMydwhKeA4CiYMCqb3gJbrIGst8tD0ONpTJ+dKpbDRJLbdD73VpIdRYXTQ
JJWKaiKMKzNsrfZzc3rPDUXzQYKoeB6M6GUnSuQHK0rxlErO9GbOXJhdgdwASN3SiP3qEtiZj3pa
WPUmMkQaGDxfhZ6Ly8QzB0+vyDnN2YLR/tercYPb1NWgGvAF8JIDAb/nUzbJFPCiOYFxR/tNaNFn
WmDjDE3nS0L+P2l2jzPD2TF5AKZdyy4O734wTMURWZxnvKd8LysepA4kMICRkTareRjjoc0jQAwX
KrUpAraOWhR+JYr7uFJwi6TbY080Ti8wojrnhrDrqEy9luoi8CfzcPxi4MfbV5I2S2lQ8Hplp0DG
fdyqlL+5AjsmdLQoo/T/Nkx1E8id/IgJU3tgTBIO4EJTgXqbDjx5Ea+5YlXo+LEQrSD44nKKI8JI
y54CobznhMabzvacV2StQE0vUsspQpvrYlCfWmzHXcp+9d7X/ykqIP0GvMzwZdMs1jUWUEsTmNTU
e9OQURFnlsTVBI0DyCDeFNf+SWnuqWOinMrEzs2MF7rE/+aaMSkdX/ksag74x+FKkCj1p4Cwg4Pd
/OFFEWBaO+9dEH4xRBQfYj1l5VHHJlihfRFEdqRWlylpSxzQqMY3je2Un+LWhAghad8XfdOSY7nU
P1SfSDzJs8Pmdki6GztF80z3Pt+QT2+WcbNe41zDxRuJboCqs8RNhigoiCh9ye/O2UGdQsmoNkn2
j+Ut82fcpHTxItKlvRVAySf6oItSAe+TaZ2iEq/qyUkFbjdQUno30Sm+eF8/SYMg6femXpSZ3ctI
Y/38NcMMKRTczkObS8ebp97Qu69cBkx7iv1PlBRVkX8JXgrVTq/ZJnJqG8zOisuXpiDg6EmuiyEb
Z5WmrPvGrI+ZQoDkLkPX3FQmW3YNVT64ablD4Z1xrdWbCsggUOb/jE8q0IPpIAfLSHhc8KG0vT/w
mbD3AOazOxUo2L+iHxqRWAVQNJFmhibzmpeN6nqYDmcyNCn9lqtRYxtmb0vDzXPKyP5AXl7uyLya
H+T6r0AuqH6db0Ah4BjwWRnrq7S9PI5g4ZqyPBMmjdL4T/9peAUyCmCCTVWl775Vz4Bhjp5jHI5s
1ETZjbIN7B30ASzi2M++ue3VQ83IFHr+MKBPmfqLAd3PcKcfKhy+8W5ySZznPMJBlQV8P4MynsY6
iXOj9/XsDEsKBvMtqtRzoH0mpjAeZZ2gdWj6F+8NwMB8IlFe/F7J0WLtrVwUF96RT4+2Wjt8O/WZ
UijmpZuzkCvOWnNACr5IsSB6613/KZ0A88sspt0/POHmqE8/IDBAPRdim4qv6y/1hhJ8zSTOXeMI
/wPOb3BglzCqbXBoy3qZMCf3DzOnkCLOqsFYq5qnoldc0rcS94EDs0GgosLNKBEQTWi6eV9YbPoG
ILN56sGXm0u2w31P/P7oOmsJXhn5DDebTi+b76iVxtNgXmlXxzWAKNBZOd9eTPN5eVKH/PWFSViN
aUMAVo8RsrRftRJoA+6w+oiO71q+7d0heJSiTl35Y37afdgXWpUqPGLyECpIpR7YNW5lCoOGxAo8
MD3bLvoq3uWpdQjNid6b5CQzmjcQ0Gwpv3mZRs9dekuXBD27uKY7EIfaiIpfL3vRVuABYPm0RQ4O
DfX5V3BAS+RgouOb6Vedb4ROdhtbSzkRvUTxUuI7phqjja/QzVGroVMHNpqKX+ppU9OFTGxGN61I
BJTTSzMTKntiJZDVBPn60usddU0nGUWhkZIoJc4bo2J9WI7DcleeNjmZIXf1Y03+stFVdZXzUUKM
IqBdGbMsljXSuGe+Czik2zzLTsBxxYc1fGOdoIHV17liEZ7eUFGNBsospbwwbJ0DAPt9k6FzLhO4
nEnNwxh7IjAksttJegm5DMDfXOwufRShGr9QkrOvbkj+JOzoNRnhzyTBtrFXRdXARDJ9K2BlHAYL
Byrz5rIcBmJG9d4y98twW90HPlmFOCJckIa8xNFAoODUE2YNXqU39CJ8nJZMnkJO0MnfNiN+eYtD
VpbmQU/+K9myimpDLZnlf68enwiDQL5ajoBhNU97t9xfUIDymPxyHJQvwsPvIaDFoq3n+IaJog6i
2Nv2zmiMCVO8MI3nsPClvdmHkEFcvHPQvTEHdjT6gsIA/Pl15I3z3AfuVThxwOKjfdrlUB/990Bl
uox0mte/YSFC6cCgP7xtffZxF1M6Q9VcZjMXIt4nI6CKAKz3NmDHwAVjDZOifNc6k/znxvXZCjL3
qqEMbmCSIlqdp2Sj2ZijxXgAo3B9bRcRqWO5Ce06orPEo2SFeFK5EvUP+9+hWWT8bud9EfmwiPRa
Yma2BRMLOfKTpO3xe0+xUR/A4sTtphal60vDtS++CATMzKg8AhYmz/pHPKkxKc5b0QjTGDgJzqWI
69J64LJg2PnXiTe1fcix6pyl1t0dswLYRjtJ3IKzdFMT65lVbY/8XI8c81dITHCQcvAKS2oZsLTa
7UJKEegC+lft5l3WIftO+QdAjOXYE1ZAYUxM4K43Wve+W4BnFpE6k2L4Uv8wNn7SY/Ih1fnSfBd2
J/jHWbVOeeDA5/Ptp6ihLByiWV22X1df3lDFWeurpYUb+/Kva4T0DV9gjxPWYFKcPkpkpmSbgARI
72zuY6pd4/0UkXSjHbY6sR6Tuw6KZCUYLOWraX4YjWWwtS1KyuXXQxXGrvQaDqyodQAA1rnAZEr/
0incXtzdqzzpG80f+xt/5mP/MSUg83f2+dDQdVaePXOzb3oLDPleA1hxvtTqtgMhQSYmZm3Yymbx
xl252nP/L+u6CdKcK3eFNP+N3neKa1GPuCwRLygalObV5XL7L35z50lzGEFb8N1h6k0ntSnKvcjc
axP8qQlhx7cSaJFeJo7b4P9BITYoiHS9E2ICVwasl+sgtiQhEsQMG7/sN9EhmsXLnX5O7NGnRQq2
xr44E/1VndckNddxddAxStJF04v+SbdtKSrjKDhHY4noCqBbPaV7qXBf+h9uG0FL6q5dh/kn69v2
3gHhMDJyQ3MQ/bNuolIp+yHNvzzqmlnpf29FuIMMlDwEpqycIg1KGzAbkefcPXk+rQ14wPWShV20
4w+B2Sn53eVxXGoDvJOykoKdIGAul6CbfulvdJBZQLWrXLcfRSl4LB142KDtB6Zkuct64+Qu0gE1
gmBaaTwjy8UPCfQRsg+dNgzCEtY5m5vabeian5smVzmPiW5A2iqeZn4C5pc35fCOPUELC7/rWxiR
AvwBjpT442q7Io2zHrN+Eadx5FFEnmoH19YacxkAJqMjoeZSwAm7c9eIpEv4RI/LR6UfZ7VR8EJS
HNfsFAwWF/vg6Fd7vLnhugf6S6lbc9S0cDdwQTee5WbZ+i65gdmfJKLMRR7XOdPrthqtu2uu4Hin
bF5B8mLwBMNqJ7+AKvjLzPuOtpHOSyMqF6HgZqiQxO2djdIFDgat1xiI0+geZRFj1sKGKJ83kkDH
/mgIIWuELfSzBkQzjoYmiSlQQz7ngu6IjEcdJtaZGR6dEqKqA20ThViiUlgiO4qDfHyQiuWNVhw+
KFKKCknprfUYe3A+63zegALbQL1p7L3LwJIAG2+tggtw2dWQnPhwfgcloLats0yVeICKanbHrcc4
X6lM+XF4sWyELi8iWa5EMn7tWrp8YcsHx9LALPVOFvIjRY3XfTEWOsYxjmqJUhv07ghJ3TGCisir
rQodpHxGayyw/p3878Zirob/ALvCRBKj2S+Q4dosXk3fnm//n4NDtbT+V9tu8SIslwfOSAphDSB9
QcTVT1QLOFDZ1HMrEWBMeEqfddElbwgnpPTOXxRJXmpIPxc1WYViN1Q5kqVTVw03nVSmdlFDNxtk
2SZRrrnwDLqdblj5b3Vs5i3EjSwq+E2E2ZFgJLFKPRylFtLI+mbkYUe2ZoTksP78d76hGO6bVA6c
ATWuwhGz/olRaducr+j5EFv1fptcwZR5e1g82ZQI3uqrgB8VBty927KYtPOlRAVT9RrnghX9tpKh
gvyw9ghyZ72p8+LhCgRK4JcWT+iTgIz+YA7lXXzYYIV0n/t6N5uFbRuqOoG7vojAXIAR5Vvatn12
2B7iHBsMmNzEYbKKKBi3U0TSDMKdA+9M6VxPnSm16IYz3Gvx41Q3ZFdn5xXQ8AcKtT5cSNNkJxEz
3rcnyBSrZA1enRKUwcQgruGiKYQ9xOT7+gMU2JDKfmEHxLHOqUF9nV/FVQA5nuwrhFC1Zg0o8p2m
+t6rHl9RwpWI1aHd1mktqnbLW8JYy5cw9QHOzMB35yUNz8ogP2Dp6DWjoG3lQO7fgYxudDe0KrsG
l05vVbe+Pf4M0xptHnPp24yGg9+R259SBPK4jGkll8s4gn2oJXroySgKiDgd/JXI2Je/sxBj1RB2
rMmH/SstLJIwheQSdPsJX4VNVMN9oBrzqbjr+5US64W6+AoVDD6tuSww4Mh/tZJ4MIv+Hqs8MVW4
fXFMyyvTMQCaW+NUQV2p57lfVnrD211U5oKrQB3IwuIDK3k2iWsAwLk/8IP4hU5FX1+6WYSUbyTE
IlKqvtZY+JAoD9p/YpfMGrePUUs6NKfN7TQC8t1ZEO7O3BSovHEG0XtZkILg2cQ3kxaHN18K78c0
rBNmKO1mspLpInEKLqMTqx1xGlEQPZTeUJ4qjt91pSBM2QN8m/qk5n6lLuH3H3ofhdB2lkGvrJsn
0OxXxk7BQgDGWCNDGdhspDf495dqRSglhCJJYgfc6NXEQ/JdG4XqhIPYK+KHgRpsRNwqz8LCBxDl
n4if6JsrkuIUhy0epLDbUW859HFJQ1+r8UjD7LQmSQBkYGseSWjIXEnICV6GNy+1K60vH1CCGY3n
h4hoYvsIbQPmFxsmoxqvozl+4fQBBzxirAEMKncTYmR+5z0exhijumQr7IUb2U55LqfLxavqu3jq
veuVTsAUmWeZsOMX6+Z0qCVB0LMPn6DEr4hhig1AMGHKJGwdAwowzLbSovSjK9fjaW9K+NbiClFx
6z0szkv0Yukt2fIlx5gfi5JJNo3c/ppQCR2n/hfSEOjJDkYBzMoDMQvBXysEtazEBkZzNYL9wGbW
0B9rpRFuWjRy9US8JqGWDNSO81jawk0lLVqgVUrd7rFqGjGelrmSSLIgGzi826HsfK06HBZ1vvnq
2vkfHzq+D0hTKnmb6kBJ8yjZnXjlzetfELxmQtYvoL5vlf7088Lsejyz6yX7qa8xeLnwElr2Tuth
vCt0iy+JqqeHtgJsSCUAe9meXSrSd/SVkQUHYC/f0d3u8FSvdN87S+YxT2FwXGX4GK89XIVHK3Zj
kfn5brajg89NjBa12M9mptPbQqJ3rf5DJhvWGGeFRCEq6+je8tnrogI0Wi85umq+4o6ubWFv8C/r
mOnjB7XYhlVuaezCZTfsZle+GC9UOHbmWP4MltbNdnsN0EROv49lzGx36KnZ0uQCvh2UkddJJPdH
I+qihh1xfLBmKif7lyeJdWFS98LAwdtjDeIY46nbKUYPWDJEI6Es5OQEwHzRUzINfk7aRjJTamrq
yMxrtEeK7Fv87pMg17Z9kC+83lZ/eMtgWIrOoBt3U7Ivs6uCf2XYzhPmkBuVntsFX4BmptsDCVmu
zasybmVCAYIjOLn1MjLT+FklhEtNwx/OA5vcJPBx1qxEdS6J+XHn2RnbBEsLsinu6SdEpg4Bz6DU
mBf8TXbkddJc9TQO3cEjo9YiGdxfm9Ho7/gz23+ob7nhQzwz0IfyetxBgc9Iy+a72BfM4VlxMDaG
+ChtqPqMYdeIxqS/I10A9F983cjIyn2TYHkejhN81rD8r8MWmL9KvjFoAV/AILWgTolYKnX/pihd
1iCpKT86YBzlRD9rE557yen5SMb6SmrlsRA5T6EgTZZ4MIigUCWl7QUEi4siE8WB8LgSkiR/57Y7
VeH/lESc4IZ2Z9dH7+BK27LnUKzwNqLjQh5ZeS4gV5DxPPej8FtFHU7XbFYtEVbJwkKiipGKWV4e
W/4s0Df7hkgjFMfxzJCAoRbh9E05f0f7rVTRETKA4ULvVAQGf7SLm9UJF8cr0Dx29UYLqV3dX07J
CDlKln9RjkIGuX2kQVyodfx/XmdsAZay03TcN3v/QL3tcNf3d25nsw8nVWATUwd1B/FqEBO2XNbF
pvy29UcRSL2+cR430UqSt9V3TxwPq01WwCdzCKBK4DkS0Fc9OfvS3mRyd6Ynm37wwIGjdfhirLnV
vcmD74oYeEWu51QZ1jMdqChdi3mRgAkW2+9iLer5+MAdS6GZMrpLXuUDp8Q4fw+f3rHzr6ClnjJY
FlUbxQe47iFl9nbO9IQPNMrRmeytlGqPKhmuf6qVv37MtZ6tlowl6XxT8emopqnxUmEpZRXyMnTY
JcChKg+AYbTBE4dGvcKKhtfF+0mDo2UXXY15N4nXKQOrRwo4Zwr1Z+ZyXP5qTozluI/S1No+M3dM
t1nIjyA2pDFTQirqkgok2MMXh7t7iA9nMo9G5bU5TaI+sEEl35B70TYJRO+ur0xGqJu3OZ7FCgKa
Lweu6AMCGr5wAxj/6rLOIBdGUDP27WKj7bqi61nq46nGeGUNtlZbUio8YIrnjpkCF4xaWBQg8uV0
XxiVr2jydL9tdgjBiFFPc1R72Qvq995umgsfa6WQfQMLjSHEh0s+rs/Htvttq1xTHikSc95ILrYj
3WpDhb+fl+DY+nkK9jLspz2ZFusyU3R1ree5tyCoQd5sPHY18IPMfOvIHB4mYZjd/BGJHupyhRvX
OMSs7Da55pTPwT3M/Cw76+4d8ep9/HBpb1EMUZKy8cXN6u/ocyS6WilyEEJRdW81aCc4ElswMkww
5ERlgCodJr9zzhSz8CCowDMEJyvNP9H958SzaXnHVaVc8UZf/jAaS/uiSdNTWtOBwSHWDvJ7zt6h
PBN1D1/zjnxhCUDzxU1PD2b0UBm7sIdk3B2/NjLg4o/Sg9DSRwPfiyaQyxn8/t2f9eNnRWB/LQVU
NsebMlaeywchOOa4KWUlPfVetbt2Ab7X/TWPMjLjvoTY3Siapmocj2sfNDTs4UYFoyWo2rHHew7m
pz1k+7hiimDXC6/kK2jCV/632CKzFSa2qBI3Ob6IJhoBCbBW2TgLfcYhNpbxyZvOTEa7Et80bzIi
mPIz4czlsIT6bH9XceV636FTwxWqZT7ZBhiVpl/fTDT0yh7qYxl8CcMjWhNWnVYqLMYdNDq7dIrK
EoosDOw07Lr2rBNXzN8DJlE25sphNTRJJMzCufX3pKchBNmLeYlPKpkgvD0QC40X2f+sk6KjeO3C
SA53430ZbYEXKn9i5B35d4ldqiEbC4jWWO4Lqgx04tPry885hXKiDdFTwX4PQsgSbFfGJAli7B/q
yMBTrvpAnCop94lWaq3ONmIgEd57+ZUmz5ysa5s6QNEd10VbR4GQYTaNKNTWuwWSQRRcpKEflPdV
iXwJGrZPZuR2yCVtgEGN5PzDqnVDmPL0G7Td67pROhAM8ShIQHL+lSVpQ1QInNgPGngx6cfuuWxb
5pDt8npGOu/n6/laWakErbczVDZOaEzSiFh0JFh9y7io07H9kyPrWRjBeKORFRkzwVKlKOH/fbNA
lz32kw/ZEfg0K6uVUOSxlXYqLRlo53Le2ANt0qMsqrRcLWYEWyGHvUR2Fgr/ZkA40Oa+ei/DT2OB
zkKca1UI6UblaRLWntOXdRm9EebF1rpN71kGHbKPzC8587E+NKUBiMuPP4MqfcBbtSICxfWPZVjS
rDL2PuvuWXcWTVTmODLig843w97KZDkNihStTp2HwvOO608z6vGUb/IoyhatdLvhiZ8ir5AUbWff
L83owDieeUp7sZZc7ZL1WGTu3u/2d3n5Ml+zolktj8uAhzeMYguY5fNAEMxFgcWSEsjt+OrImwM+
644MPl1VdHAf/8ykieCr5akxxQlUVehGZ13hKdLP3kNHW7c/DLAY/PDQvVhDfcCKdTRbF3vmQsJV
1MqrFq+ui6In1Bw4iPI/ikOq1n83kRx6a/HP9ZuilL+TAvVCAGudbhmFQA39l+3QWXdQ/lmNqDor
q5XRzGmpYlhbuHFhQL4en9APwD6AiAoSZLvOg2euytgCVOLaD5QAQPQ/ilNhVs8/CT2JJR5VCLwz
Sc91mx7pNaUhC9hXVbdCGg9lAJd5djrXR94v9OOX0Y4cfOWPr3rw90jwSzGzXnkJ/hzj56qLwkx7
eLnk/PxkRMOmhIwN7EyW2UR/GCt5nMwN9lMCGF8bnphAG7CF2b2jfsmXU1AnqmBZph2FmE1/w9T8
xLfSrYLVc8WVqPBCsD/W9ayKlrifitNv4NmwpPfk7hmXfE+ZzC2v499AAl54Flm77XyyE6GUh6xV
1t/lG2vDILnB03Uu++3gDF8kBqByJLSo11OKMhArZfyEs1NrQw+NTFiZjaBAm7Nxqli3xgo46Uxm
b1UXmIQF5QaUWfICFZJhtXeJaMkeF1zWO4ipBj4JrhHG0XLsORBTDNZvUb8eNAbAy4jR/ZwCnn/u
QeDZn4ft3oqfrK9GrU1S2eaLeFcUwr2ET/EWPMsnc0bvWlj2lNUsSjtOOH1aHxw/wix+YwP/kVt4
D5EKAOGmRm182wd01LxBqojCJgJ6p1U5wnrHEZ9RDvQs7l3VoJs1g6pb1StAZpJaQAwIa8f5l3jr
06J2gc+/w3nczF2wG6MKmDkfFItHJFkvE97yZ+93NeOT36YOaFMqg2wR7W8gYimsXZz8OdcEJKk3
Bcezwqkr7Sy4JyHuiBsKkZAF4XK7oDDVVSajhIPF86ws8pQ2yl53XpK61i/uI1XA9GwskEHJ2rIN
ZEI/87vyJF/x2q2z5U+sp2tLHDK9zrOCMBTfjmlhu4KFscjOcu6XI6v0LOCuc54sR52QFSRISQD3
FT7e5VL4M+RFcu87dDfR4gGs+Hl6dKL4zmAZs+jNqIV7A9/XtTocfkc+zNw3/gsbcQy6w4JVgkuk
cVbLuZA1EKhgmlTI0GbJJZvNhyfNUCX8gaKCZCo6RES353AiO5/1QuiZCD4vdsVqZgVsVn21b6Mx
FOJHdjnKeVzLNT78oNuagEvVQJ7DM0nSY97nIJ2UDawz629NFzoIe0rRJYqbzKPQAHglrKfRZIyM
9uM6WFoHQEuAxX2ifOmqMq3vFwP+c8LDLtOdTwckTQ/2IC05LV7WVAZAUHjwscTNxN6aFMeTP8Pb
RsNILdDT4/pC78KfpmoQD8y1+2qq4g37c7qPrpIM1dTVhfGCJQ7CSgzSetg0x+GbwOlVkvstD01B
ILCGRD0qvlF+8mZA8e6Hz3zIZ4EyaT8iArA1UDRBZ0Wo1W7zyHX1QTtvGnZDypcj+vwoVBDLDxMy
Dd6MNdEuk0QLidAkWZY/0WkdV83e2L8HB+Xl8//Drp6u/0HNHrMkValN+znefvIYnkSt8n9h2dHC
DFEKm0pKKUjAYz+nL70EE5TvEVcayJbFpkT6XDjQkvAaFB2K3oqKSne5qD6XR1UnFo9tGLzchMkI
j+vP49YXnovb2UD7rpo1aq/WNS2kgm9+dhqnUicc8hjPZ+IgweSTH1uzrWILkI4biZL9+lbO9Hzj
OsT805ezbQAIvqm9obRlRGBrCFVfTvbmTtLf2nG+i3foz8dlkVtIgXCvjNQ2lcoNgNid6OZPgTXJ
psdV/zzsWT1EOoT88Q5BZbtwkpTsDK6KSMDiZa8RdI7m3foqK4/sj6Q+V7zEh99rDfHoQQX7/kYP
zdzjGjYfrl8DxvgWkByrd2EuLyN0kpwl6OmgekkRgzP4SbISuwgTB7vw15AGWCmSDrh/GKfUCofB
j0O5OeV1L2EsIXh7dw3cudymmbWQU2KM8R2Hdw/Rrqk2cr8nCir1CP+O1WOphAh2H7+SUe3Mbafj
Z1PZojX5dVFkwheJlVA3EHHdUkdkgZj9XvDlSngUACIebwb8IgTeMOYA7N+dUVkq44wO0Ao8rHPf
Pcs4UpKVTRLWqtQHrJM2/4c6chuXwFgUucxvk48+Iu5avUfRf985R2W/+tcbTPv48MuEkH67RESG
6g499fHUPXrQ2mOrSejkEVHV9eXm9cRSjeKI+BlF/6Opc9Jcpngai8w2pMAvli9gwTRX5NKUeI6j
rRzQYk9Wla22DuITtasZoT+4DkvmZAHJjOfTtzB69eLL8QMT8pd4+O/IqqvaLBoojcmuSL2Ra3f0
C9unslHvwGc/in0aO57+BaVAEbOVqRD/u1iqwlZgtw8OFix0R1A/dEMMaXOalD59XcAUZnZqH1/7
yiDARB8dCasizXs2zgJCFhHJ237chGPZQwLterNqJFe+SgtbCGxD52F49DJ6UfDZCxmTQPxmnr5Y
RtaqgUi90Gwakni0oZhvXF6urLo6zc09zVe6OOliKHYYj+RSMHzKJOvmAwYKGvOTEF+DgfQo27cg
Fc6BWp5TpxEEXh39ezqZ/jNv1h+VKDJ291lYE+63I2oHxJaOdxiAjktGo+DGwJb9KURDmUSWFy1p
qF4TURBopOWz0Qz6PSRM+CgpPN7VYMWyZeWjcmXSZtuWIkKZFNbLGEcKjKqE5UvR0Pps6aT5GakQ
5B93JO9AUVTeqJpE2PrC/h8F06wGia1kEr2ZmIlKy5Zcddg7OrndUNjJWpoxvEXwp0lOfAoOwTn5
WRFvBy5QcUyB4Vnfz0Y80NqL9gfc4Ia0nfWTuqtACkVmi1ChDYWorY1sWzSvLyjfQXE+oCsEUErW
KRUPOcldklSjn1cuIRs/qRzy3lJ3moVKuXWiYlHqaohb7GEGSfa9dezY6nLJSY36Btf4Ss1jMEv2
lSZSRO/8MkHhOEiz96+WSNyKiBokRQhTf6HmzGXab+OaUdZvTdq74LaXCcKVOrCL1N5N5BGZgmqW
p6HJyACwIrSw6Re6fb/Fwi4180wTPUKqA0GsqsuIk6gW89O8TtrBQv9DM8uQ/owFDUW19PwS4e0L
RmJ+oQfOzgMJuuJ3vvT/qMjq7mv2SdrFwFOSGInwdDgufQr3fch1/OfuoEWYDWsYNQjXLUyJ6Hq+
94qDJqABb+yUHuZQdx2MDwOYNCXvPKhcPy2wG5ACK4xHlWH7BvJU++mwJqtOIpfxhjC1AAbfkS7h
A7djH6hYxuO+Y+Tqgch4QfOuwGpuPQwJkw0WP2WnyTQcoPIZMEx7VIHELsncWQISMfRkHeWBaTWU
OYXj+sEaf3e7bfApMnzKIo8D44xujXZe/mFk9unwU42hgCfMaDNU2c/5ivRJjOUM8f2sVXdNX9Ed
qIhXXun6VVm+l1tjX8Wbp6yykht0E5pr/SMRePbL+NVaQ6akog649rJo8TJfL4jLjevii4JgcaE+
A2deb7//eHk3gR7a+BE+sJ+ID42VuaFZXbWaetpGD542A4PNWYT/Ab74Jf3AjaVPqx0pK3T2O3KS
6FT7w6paxn2U9W5d39SKlSkJj9YU7ittOV9O8JsVZE6PONk1ofwNPnet/MzzhOMP5Yyf8J7c8reF
O7PGXRwa5cMsW3qOtjOCjpyI4f2kb7MSN1nX5pGAmpFbWYem4MHTGCP2j3llSXkSHCbol/RWfE1D
VKhcEdEEJG1DLoWEteoki6eCx23yevAX/wXRODex5mM/p/IW8JkMgnZtSLWdAd32mitoNIWhjjOS
xcITZ2t/EM2OLgBDFPEZ7J3Gk+zHGFBJsLW16N15BU1UTHpVKGK4ymk++7MjygjCvEjoTGn7dj2d
KN/wgU54RAZB7lJ4y2srUrpDFog0qF36UP7Wa0xWo0mAdY543zZKKlNIfShHLEfA0CAYAdJ/XDNN
KhT9h6ExIHb4VqixhfY4p8UNGFyhOygNSGPjjmc1QonWFIjyjCrNkiOVYs4FL38Pu4TIBcB3GwWT
2i6oaG7MTYwu4Xq0foL/VLYddHcVqazNyYW3D2QIkgackYEB90EUhbbHadmC7DNtsGwxUKITGX6Y
Cf3uruQr+Cr2123AV7b8AtoVJm+nVHCJmXRnU3FrTqnc8zxhliXYuhf5ANdWS7XBe9PQW8iL1ZLp
LMpMhN7q7lYJQg8nhYRmRiAQ11DNPsoC0DJnLdq/kWAPv4kui+/FXczKDiVM5sfbMlwE10dJJZNj
k28mgScM2WMc6ufIMbJuJDmGL9qNRahi5+RIku3pyPaLWoOIML6kK/0/FvH8ltzbVyCIHQEnZnSu
KQavPpiFdICUKXxp/ssv9bTDGNpYQahVqPSS9DN+9CZtUjuat9V3FmaqlBXLoKPnGtrj+AtGQOss
5ezChABZsNxdz50QncVFsjJZCJgUV8cGt+RuYsfNhj8QYtsSLncS39jLlJRsIKM+PLNwBnmrQBjh
2xP4S+dF6H6UrqSADfYz3v+Et+pvM0kqVrr5C4lf1IGAwMUA6QWzISKYL8z8g8jUBG3znW5gS/CN
iu/GXxrjDYO6DA4cOpJconP5bEnJivDyUmmDq2vILNKhaHnMSwGsYL5GjTBShZj61nLGl66/UsVt
+5ZF4VbNU9DQSusGJeEdm7l30WF6tycPBdSPZ7ik/Vcz/IfZKseKESQzVYlJj+72Z350oZcsCkad
7v6ChAGGD8isxLfbzI9lvNvb+lNiW/vM8W2S19BTaGSAYBshuc4LXuVMdembT3H6+tnYYD+rkxCS
M5/jZZ8CVv/J5xO/OjJBLmQmZpfmm/DI3dQSBy2VhEAODJgJsbhuUd0qC03LxV3AS1lSnOQ5sGF9
AE5jzMxD+gKkB+9VImHM1zUOT8sKEWQwoG84x0QG6VW7LToLWUjL+argThBdxtjCvJWB23Ccf9aL
fhYmgx47bGhTcI/JQkzda+V9B3IBQDXGU+tBKicIUMArFwEwib8gogtQqdroU1yZHyTr8h8kRnF3
u1a719kGxrUqXF4+4sV5ajx4obAehz0EnPqQWyUk7geXo/lWqhMsmSp+l7uVtYV4JH+uGm/FaPNB
9oAaep9VkcQ66E2elaxF29rTpn9EZM0laiZU0JGERAw3W0HjxtpXXnfhldK4RM59zHKBQrV3ZgPY
WJLM+Ag/WCi5pw1s0daNS5p2WYFSMmFGjxECtTkxC0gvRXyMRJ7bdIeXDAn//0MzXeRdBA6CwMXY
sexEQ5KOEUNlHm/ReJANw8gxT5ovCLNxnYTBVHBGQprXvvKXvdVbxvv5AqK8WAkgAwsnX7cDB++C
RjmXGa18n43CR7Dd6lBrzpDP0UWoiTwmB/rJMtAeyIdsGESc/8Y4asHdm6sBCoZwrOV5MWxQRBSF
u7QHLJoo35jdfFovl3UysKop8RGzqPfiafBUqXu+80k47pzl3fUftY8O6ccMe8gWNY0g1sBbA1t1
e6Db51wAkJLomezSU0gbMTcfJIg02/Ers0gQDx+GP3gAHvPwSjNUNZWf9dlbWahkQ5dnB/dWB7jq
njTNCi8OML8K2yqlJy6CbQsK/CI2ZYIDc2pP9y3RTylf75tzpEkbphMkS2wjbAuXcXwODW4SFpgD
YAkkOcZ6y9AsXs6lg3BM0SoM2lM+ANIviY2TqiT9KIhsxM1Sab3/BvjbrLkb9mpNvqsVTBMfRfZb
sVwH11mw9ItOBVSpO5Bn94du1CHtD2WLfh5uPnBlr7g47xh4dfJcXetqDMY7k3DcZbc9kXCvtTx7
VGGMJiqCTU5u+Q/SonoradDqWBXJcOBGZfNn3hom65DYwhiMGa1w2vAOcYaBP92KWYakbAK64uFu
C4/mGd9ctsZbygYtMBMrdugWt7yMfaI3dGK/nCl9SRjbd8GV3ElK1bBywPqxk7lEufu8zKlAylgk
lvgoG2wSc2ChacE9TtMmTRG5yku5jOu6VqXZMVBqk2Z4fEbw+QuvP4dNFqUZvjjS7m8ymeX+XZnM
mrIhP8feINi5jn4Qn6KnJJZrn5c0yN+NtF47L5V6R/NLoRsTK3FQ+WNy4eqdtNsg4AJc9A444/iC
Nhrj1Yc1eFaC5CBT7sz67/nu7DsTq8NFchsxUniGphNEpreIL/fdwbZ3fwg0TyN6wSMAsdKzn/AA
n7Ti7/PjIgeoePJBU3Xr5OU2mrgir4RG7AKRUg2dYbiorFCZO6Cse9z/8ri8tgVz4vZrPYk8yC06
6VoeWS9fQmHATV7KXULERn2/rLwaFx7oTy6cTIEGBx5lVvwlcP71MZxSjD5WuuhqkAoZZV1y6ZZU
rQxo6E/2FEnGP7kIVsHrvAmncLoWeflTGOfoBRQawxCYNrq/msbkvUpSHFqaKm2gm9R59uH/L1k+
8NG5bHF5eZks2YoPBt84MTzToa1yvp7ip47kvYwjlu5kDUaytGR3Xnz4TmOTCTm47p3kugqAc3NN
HGdp0Xf+W37FcE0zh1SzTiGq0UsS8Ok9jzQ/rMJpMoXNyrYHx0j7HwmMym3u6OmRqA6Y63kQprAt
CvbcHErldmmy/Kj7XcxzPRi1DVuADAYv4v2DUBCN21DWjKq8YUilPvgN4ACm7Zh9V8uU1WFyPH5h
7BXqq5zjxziraz6vLu2FGFjIYziXXSynEOAyZOXdltdq46ovRlO4HaRYALJxtAuO2soL6NdVbybV
IGALrND/aiRM1Wudu2ziaxyx/5VQ/LDlsLAW8FQ0kOKkrsEem9+T6StRDnXbuukWKlruhxfIP2+4
kLN/MQg7gTXujSkU2FY8RlkOzTD5zDjIu6SbouMlqKbeZkEwFTqeWmRcmkcJNdgb6BOOwpxIgCDP
iH0SILO6uiq4FCLk9T8z1GTtIaDsK4eO0Ff5U6Neasc/f9LJhwL+syK3zcz3AseO6xjC/kTjahfV
miN1fRA3MIXwIDH/qcQ3NHxaLtPF31U0efIox3qRyPgHbTN5ubQbvnXKERjW2evtt6puW/TthB4n
sMfQaA8g3ixG+GbXlVMlu+JzAXnV7vpuSalsRz1P3E0+KEIXaHKg1wljHUts3HcZZrivwDyCunp7
dem8rMwbcd2RCi3PxDm1wFVVUyUHYtZbe/lQlb93M7Fdr7Mm9djPOEqZGgO48nBFEBOcfUS0gKIh
e9FTfUDWGvznriScRrVSLfqozcesdZ71tm7y2i12Qv6Ee9ocAvKr0Gyo/xbHF58Y65J/GqIV8X3O
DPCTCzSVbWoaC0/MvDrUTQp0tUgigxB4ilcbIoEYKmQyTwYqcb5EK5227GVvQSrGezbojracTjJG
ISRA3/z7e+ojrfxGm2SpyXpFdFRXzdAEhAqbfGv5lY5ckTIbRFcXy4dQj9JOXTOXFxTadgoLREVS
7mnbNtkkabwbB5UiX1z4E71C8ILj+OogL1KFhIuvc9BsEBGVTSdNucMM/VADu+JxJmmve4Lmntf2
xJfaoJoqJ4LnKtNTFqZTpthynev3itWhJW2HBcnELy2TYEhZ4MVcFNAcSKz/LA1T7Se54b4HN0dZ
EBkmqTy9bTQZdN5CY4Gb8zLkFW1ijuHCirdF+TDxwM6f5cQnu8BRwGQjVbbF5UaYInFg8EmZHtBa
E3phm9xjlIKkBxzVMzXr3PFScQ6qXqL8B4A764tawORiyDjT/I5vzsTaUx6By0R94QsFsf1hbLxr
W/Mx5tL58PbhT9Eg2KK02RgQSM9LwbDvx+2jZy1pR52MY2LZV0cbRUZAwzCoQcd39nZ2BbHXH8ib
pgc4NP0L4eOxcWA90rpUU5sBlVhllI+MeQOLq9+MX78xsP6+p1kdnSYlpdCIYpENTU2+zXYlUpca
W1St1VdUMLd6FoDZ5z9I7AYszTdNsI3Y/TsYXDXpXNwdna+mCQ4j4zAWQAbadi0kV+48X1f0NpsG
cjVUkSJmet5QIV+9OgUIzbINtE7K9d4zqpKyY93InaFriybq4Vp5ZeULIHnxf3NT8n5uHoc2Cztc
gaAQDKESU3hlfZSAt+Why+hGSwWBMu17UXd2ewq0XB6zwVErgVtXeqT6J1p8YKOdEWlTIhUKz7qo
2k8le6R1Nqskk+BMNU/he/ZAxO62drlERqghCeHn2qBlJp7a/tVJbSFWDZh5xa9nSejGSU80xH0B
BG5+EMsMyWIa0QFXBcGRMcxn3+Oi3WCLbFZjBF0LIFS41hheAElhSVMMrcMJD7Lyc+azwa9vNjSv
ndjgFYG+lVexhy+wPj4SYGHJpVf7FcPXN0wdpfeUxkGB2aN333NWW6pdSwwnSM8/D3nJUYy84+Y8
c8oJZfBK5/juEcPRqOJI+ThP8GQ2oJ4zu19EqgCr8MJzwHWWWMTH6lsmsf+wb+p+Zia/ue0fmIsq
3vK/7R9T1Ykap+Ib5zqD17OFbWioxb6A4iMRyvbSt+LYNfcKZFtcOFsH0vc4yqI38mnHJ0BzV3H7
qHc/RglYpVabOSDa9qKOHms30S2FIDwMfkQb4EbcqIAjtm3xn66JwGKwSo6iC7J6rvsG6F4NJXKy
A83rJOxddK0yC1cmxnlTsYRC5UJXn9+UH4NFWtE/ntGDnmo/cSQndesdvn4s5RFvG67Eh9M1SqW8
nqu0/BG7wSsWOyvhhSqjUhffNxiDfxmVQPLZlsivmrAxXTnjx8ccbMR0HbyZeBvndKzahYOwjejL
AGDOJC+9r/f+RgSz4JgGrHbpuOIXgAY8hxeuK0su/no12fK2xvRBZHHkfGv+kRB+kTKshqb7qGfy
2PNINJTdQLmmcafx2atGob2zI/0syBRljMJCwKt7rUJ7l8OoYbh1+4Uy/+IhjDlK66neSGYWa0Md
xJkLV9nB8PIj5PaFqwSbk6L6oJU7yMNIHER349l0WFFmhntbQQFm0KJITX4d9i2am6/t0mUp11tb
2558WxB6nz/sBwhTHqqm3f0cZfwmgAMX8hAfSiCkkrv858r8wkf3oYcF8EF4ryO9DDMDZWCEq6ku
9eHjd2loRcHZ/xSOlH+b6YIadYcmTM8pRXM0xwGc1V2eHAM6sVXl9CYSF1Y2c6GsPpgVZw5zyaMi
pQSqq81L3QhZFW4permYOM2HxEebgM3L/KmHsVOEpzUow17MmpkaeqZBUBTUL3202Ayz6DoGROAz
s3y0DQSLRHiuhttedfrNkTgu/35qN5ju0go27oi75S8owonsBPouu9vZPXJoFIm67FoNIXMp4BcH
QtF7FCIGRTHWyqQ90S3nmC4wRouYdYCtmuJivTspk7CFpEM8DsUBYPNPd+JBIlMouPPysHUZi3F6
m8qq0QFWUhCIly1F+p93Vdv6h28owmqEVBkfk/deJTAwcZfjEudBh51G10BBMUmd94z+ZjB+336j
GBwnQX5R7CphaTu8RZttN8C4DiMeUuHYMceFn9Kn6plkc74g7yl8rTgUSz4c4pLa4VsL8pxS+tI/
EX+oPf9qz2H0mN790mAvua6elaUrqdzfBvaPLyb3ANALc8UqEsptuftgK7sTLaVQwkxoH+zesa7M
XviHYiO1mGD4Tl9xBdO+uQE3jTkhv2aOd4HTDwuhnlnTE+Asw9++1BWZyywXuiVjKEj3LfxSVsPA
vY4faxLWCU9ukVSisb7GmTFJ1oJ6rYJTailhYZLF6+4MPYwaKp5wVuLxNoQyxUTArfcrWH2+XStf
F8UHzlbg822ydnZnWGtwN8q7SPZbNOQ6Kxf5tWcgP65Ysfc5+Ws6b4/lldyish9sKwuzvidmtUBo
kq4/TcAblVOOUWvZ2JueW+mdUbQ3fIDw3CjI7x7yLuiZyLeSakD6xKbMiFIqBrogXTomTrcNcf3O
deinRhDmk8lw2f0SdMG75FQtJlU51GjUnTK3wPwmQxMMUKfIP0xVLKUyeH91lAXR9FxNPB+g7A4N
TkCsAnVbM1vZPPEv1ddlwci69/F71N/ErBxHJZ8beSRzCcUxqdciH2pYNOFBeH2ZtDVnfYMPdPki
hGswafyLf42K/4RdH1oQYyABeGnjST0B7BkRlvrQURmaIQR7H6pFjMz9ui8cBevX0p4qyIBOeYtI
Le+zTBhp3AK1cZZLAeYcGOfvcFwj7Ol84XcGQjyYBtnt5Vu57g3dJF3pXTMQBcHxUDDQaY5gg6ui
ZMCXzwyHHPrur5bZdI+luan5zfqiPCAxVl+2AFInKce1sMEZZ7/EF8lwZ7JXgT2FKsrhRHfN/+9z
NeEbnINr5jSmN4SlbAT0sx0IXToRsJ6fhFa+IBI32xlBjN9C5hfiRn50Hp++U/k6hqgexAD16dHk
7MoaSS3pZbRzBMRHECeBF0X4Fgsfnjbks17Gf4KKL23xZYlW/ZVhHt/wZm77XcXfolJXHa6MZQXv
jB94BA6eoDbdYdoov8cV2cx36J8Yn+xEftlHOY36XX50qSEWHP3U3eItCQ/zJ4zPvI4pu18Zr2a3
9Ohw7KVb6J1dAu5od+l74b2PRrnbY5EH5cEjJbBBVhnofxGPQGPoDlwni4jysHMDlAMd6ZS4uAb0
byJlqbeOxQgtwDTut7g7oU0xEZl3fWvO9mG/16audpBg4HYjAbHMBupLJ9JDkyPYpyk7MxNFKysA
0CM+j7ZDi+32966bmtkYfxldgNqmjXmTYj0P29/IUmKTxYPkz3xlrfaU9qz8hscNfgJgM6apeeU9
iJfKQ69wDntOLqw+3aknNoQWPKbjumbGxZR17UyfaUwrWkM2Uky22kaIEy/ms8MOwgOvzPo3GGmZ
JZkYsrzQ9S7Hvbdx+aieKvM7uoxNnTjfdKu4zEf1fIhvYBZOX1NrY2qv0UHQYfeaAGsBieGwR6i8
In+oIdHf+jLC7AixhKjlaC5wxbPtwmIB9m2O1f3VP+vu9051VnVw2wSidtIHB/8wHmCBBayzSLcZ
0UImnBaWdhFLTHvSohScPqJLYIH0pXM4OPmUTGkTgh/jy064bjfs/0Mue/RRXap5phe4Xgizb7rg
eDpjahcEutS8qeSYs0r2uMJNOirhXSHAa0k/0lBhk0QoRPfLi/j0RNrboDrRwBg/O3hRZLIKiykW
4j9imCek5WWpN+3MeawYbpIQK35ZhRIl8ciTtA1hIb6BSrfFPMTZ/9JaGN6j7boaThTPLdHF2wf8
dR2/KDHbYzAeu7SU7KZ1dJhuZnol/4jTfb6bDUjGcEgwBR4B4+3nuUsJkYqD2/JQ6menZIk/s6HE
7N5V9NmSUXTS5kMFZBE/mtwkhS2G3I2Y14OdLHHmeHnGafgxOQUxwzsBe5xVNaer6NxxFozf+Bux
b/MDenFPFhaCTFwUEnqo/W+PkTU4ZlsD1JD8xy6iS9rNO66Ol9wVO8ECSxLI3blWMiw/U/wIaO3U
5CA05q+DeJ996n4IulIa9l7AVjCWEAtIyYzV5qVkz2+UI86tnW1qtjOm7KKWxS13y0tRSBQui7MU
cGlCewk0Vj5gJGwrFiwYaQq/fZM2nABmeKo/PUzH+Qm7Q1H4d3a6pu+Nm9RuzBF9JZtP5X3WwgPA
UFjjSjcrOuqr1b5hdKKikF4KdeSUd5JAKTGQhiRQD+r0QdLQaXf3aBlVckvC1bMDhmI0VH6Fj58M
ddrW9UNqh48YsvGk76W5yLEsfZzDOHUYvH2H+FFYI0CI7uf/ryA43Lnz3zP26fKFZ9VPoVweTZ4M
2OQ4ZxX2WAOY3c0asJSyUJfYZzt5ykywgdeRLzwQF1+gYgd8Huv//Y7KLysjUUnthDBHHS9rvORO
c/rgvxAqf6LT2KrxCK1lX/+6P/ccnK14kKeSxBwI5XExk7saqEbd23uzVMh2kaQXQ/qaGlQz50/B
z0HVTLIIAsT0ps2T1Yno8lSHZxG+HYpezS14kfIsK4g7oIgqgRjI0akIwcONgscXve0QCeYTQxii
vrkPOBZgp88FPyEyK485w7woCCN/Uea8b16y+XPFCTYaUGSbfA58lMYEhHzpKVnRJUBWDsQ/Dgcc
5xU5rNpsWSgSp5AeF0grA/ADHl//LccJ7z1+oT5RH2rSGmGE/KRmkt6IeP8J7H1eCV8CpTM7z23o
hnqrpCfBalr0L8cqBwwh/Uj6C1x33Z/Ucb4ovXWw0b1I1MMGGdKzelGN/saglPdfKs6lXWGAXSEi
Up3s87rVMYWGmldlZ+9ay4o6cPJNbJ34SK8w3940+fB/g/dYCfGilOVOBoT3HBvgRG8e+oCKRGw0
znbBrIKYxvCyU07kmF5fW1UDe59PH/aKFyd0KVZknUQ0bnwTIenMp0T/S43nWXCbbISQuEIKrQ0H
itoyCRsNtMly5q4/e6WyO1ZWh4eFpBU9b/5ep+RTUm62Uw4KlwIywTBenjqhTO9cboMUPdf6uo8n
PoXzgl5/AaaaaimVQCYJ/lDC+Q3hinU7mNzMVs/wwKfXFgkr9Dhup0yHDQXg7Km9rT1n58+edCTi
JS1+jmrs42+yK0RwETq54B+QUVXLHt7opcMJx9p3zzFYFCS2oTj+VLv/wdWswI1k4Ay3NaUKTgJ5
ep2T/OHayyxQ59x24E3HYfmED70ffFtZDsNoDYffj+qBE0INh//SvFDSbsi1IzMLLyFdaRgKlXiV
5GrhX7Sd/P7LHEujwux+8w0Oj6VUuLxkSbeiw5SB/YVj0hwQ0k/zIcbwgKagaCFqAmC9tdaPFFxA
sxyJtp3vYMFhTXbuYqKndMmN3RyXYCe7AUKegKBVM6xX94IIgQ03+GTW+Iteva0BSgW7VpKfEnQX
BiFOk6SGS3twfHJ8tg3JQbK/KBW+tkPcp+GblCxdMMhtd5dLjW7z8VaWZ4htqqL92zOVzEc0V/7f
Jnbh3M2zn1bMOqaEh6s508Tw3K8VmZaAvU9ZCs0dqWCWSKPkZGpPEhEf0sycGj9Gpz8nS8th0tz4
y7OgeVG2KduqBEOwf5f02fIB1IedsTqxPmIblTgIep++aFElNHGtprtgnHudvC2JuIZWMVUXmT0T
e8rGNfyiihl3lUSqAyXKAmNeL4FchN/TnJm/yv4ZBtM2m6wJBbu1WKiHSd5s8FN09QwixJ+hgXaa
JBGGiV58xDYuHGqasx8C9GLnY7TFKZNhue6LtwxYoUVyIFrZEqfUUaBu/mRsWY5Q7khupmfHbns/
w9+srsSs2oHOA6Mo8+9KiyR5WxwZN7BdUbyy+lU3DFNZThTmOOt079/FVqVc3kBop0jcx9a08Sbc
FLWAiz1GDtI6Vw/pH5bw06cTIlBChragIHrE/cEDWzW0HZJ7QleBOz/j0Bx3VFnaQy7vVUVtQ7w7
SKxpRAJmdQIl3mvOxLbIhOa/ob0kAW4u/hTwNTUzQt2bryqbZURUP+oDbbaeO9F5ArzrlWOzfLUF
JFYU8m1s6b+2NvBMLyMZUWql6Eutc5AsUZ/GC80IdXR5sGVGPL2WUzxDAMWrBIWR8CrsKPORaB9a
kmjPdNkWIyyApR5M+nKYqDNKDLSX6mIzGBwHcECwYZy7wTrUwo6VbyeqNKqrE2oGpUdESXHOAR8q
ldAYszWeTs7LPZDq0tT95uBEcpKMYroL8NezqvHyDRnmdkW2GWbRC96Whgd6UeGQjOe1kqblhE4j
zK6mdxc6C4UJ7bTqE8ZYu7s/Lry4RMkcVwSGyL9pXP20z28l6IvOEidCMtLXNKwN4QcUfHSk/Axc
prJVeP54v+uTyZWSerN9X95exLpmNu8BS7mGbrysHPHjHHLITZ2g84Rhs2wbKk/6+1kyrZaht8fs
T8TDjyFjLmLuHSmyr7Kcm0mt1i5fG3VaMuzgEYVDQU6BVA0cPgp3u69SAlBdKn7g7CQ0WuLRlSP7
+IUjtMTanGHSB0gAYvzXHKu/BHhAD5jdZT2mEdsdIG0aqOHoW5Y55D7Scqnh7Cv+1Bn2Mgk0u4l5
1iV9W1cAEw/+tw9E2aib5LzalwQV+VA9YfBXMeCO2x21B9t5tqJw0ZduX602PVUSK254eQURsMd4
z0+AUjMJL+XJMD/1lWjuQjdVh7hp0oiRM+5oCJE5UbA7QGSXUcxYiPbEB8pH4w68XEvLq6OYI56q
n1093Ndz6AnW5KjQOZqlUKYuQ9+1fhFcBauxhBoqjThIs2M3N2QXM1iU4S4VXJKCVotRivjHuegA
59QVT/6Eutrig+FaZ/1OOZarJuKcWp6xCPW43h+hlRcAQGWU70MyZMLVPe1zmptMSyEO4/onJ9WG
nKgdpvLs91FNf9o3I2IG5X3NdtCTbTmrR8yfHmRUI1PvfK2BtFnTNWj/2TxcTa2lCC2O3ewGmRPl
bt2Hd+JCIFYg3f4SJ9kJWi7XwzzRZvrtTIk8vlVryU+bgXDfOPiuzjVsTKpYuPUuW8dtS9irpSYk
0cT4hw05/AJEW1mQUQPOs3+dYq9QNO+TU5gGNKihC0ZEa5BWxecRF5CwmDc9XA2F7ntXNbB8f5o2
kePEjF+H4Ds+J0k0rORxRrh+vqGi2SxuSwK/mSvTOz4RJXYiskhEfqk3K6S8WKLU+P9MXkMztN4X
qBNVE454tcLgusVKwj5saSNO+z7ATlYPxOSjz6SYY1tfUc8QxTrAqtw9MRc5MeEmBIS4qkGa4dUm
XO8EHY3RD8q7sb/9L8V8Bh6bb9OYMhdQU6NKXY9NvpJy+bEwypVLGK6jfBGP0JQUkVFtqg+qJ7P3
LLbBIPufrpY5mlRd8cA7fyB3dbAj2O9LwmKo7w4Ww1rxCxR5RovMMrh5c8HdlZv6OjtyKLQF4JUN
WIlwRL6jvJZjCHJBZ4kkVOt0+/uvy+bGA38bO1N7xuW76cO04n4erF7d158lqwIA7wn6onLkEYsk
UbDynXtGWtzJE0vtrc+wrw3zWMdEJ6VJ9x3Z1Pw0pgUmUGk+eVRq57Caln3yxvMnI3jtKIw40rzX
3s3VF6rn7LY08VuGaYCp0aRkjzeK1JAWYw58DHCelYesnswFdDXJtGhw4su7++VoFJHjhdhTT4ft
Tf1NviAevTT0LDcPrZhl2SxVxVeLn0Gqx5YBKc/8hJlLQNQR3LDfcpbFl0/rBrW79WwT8YB2P3Fe
4jtbfRkPK3BMQOCQIWHyHWwEdPXhlp4n7JH+f7l+2Y5oVa4f1fazU5/DLOwvPjCpE5htsr8JRirL
SZVTpqPg47OBgrNm5Yh/sjpy3V/E6B0ohA2V+SZk4bf+Jjf6/MnmTNwHBTN23mJbXleahp2ayOxd
NULukyv2wu/JodJ3IB+IADkLGUuh2179EOmY/cq5Ka+L3pLvg3q42SVewhZfTek7T4yDyFujlMID
CLYc0zakc+NHD4L4ZRJaeRd/511DWRVtsyEeRBYMjjFZgLBpSPul1C0K6ck0qFSNYuWO36rjyIpd
yWQ1xdjSBYg0KIX0uFUkZzN0j3CWxkCVCSyqZmhRFB0V2FBxTYgYKJ1I+sgMjYiCROM8qNcWPZwa
/KBKgh9uGlIbkgUPulhiRtQkYmQjxPL0KhvAj3e5EuOH7jvbHpkIniXJIbQKT9OhY1bbz18VWgQZ
Qp+tx01JdqUqvZyDY5SUR07FnKRgyTUYJmDqmEvXglNtH2lzSp8kRkM6yCKVQmIUN+0z+1ed2aDe
ygdXjQnpdG4DgkXViMTVwl20rNm6VFOlQ7yRo/8++IMKlrUKJoHUhlSEfVWlV/vuZQxht4UFPFZ2
lXrsX5jBudth1CvhnVfs6ygFcS95F5yPDqz+hQ5h17eHhoBG4pCbF7vWnG23N9tuCX6jAkTyh+m+
LaUn551cAtb9C8xNnfoYGcpRNu63rKj7+SXdeml3Pg8uuuTZ+3QsO9EMxUJZes8LTnSOfQ5etyds
f8if/lr5iObFN1rW0MgNhINa31GgKrj8cd7kcki3D1vpfFeLmiCpSZUbn20kkDf6GK/DOREjzV7F
BahSRtLCweaahLtRSOnvhrqXPh7+DsYKlvowSi8qae10bc0j/pDmBvcKThcbp5xW0XQQMq/BbCAs
DOVCzadw7YOPYoZPwlTtWXuY+GC1D+5Cnau+1CFrpTIqvw0WjSbD6Hcydf8lPGy6oevhRrgPMosK
lzn20zQgx5BelcTw+1hTUUUFThAEXKhPpDZMYOit6VFWBu8zOdJWlMUonyANd9iTTl9j4to4WJru
zqhZvyhm0MD+hRic/uCFI54PZ2CoJqsNco47pv4RGtIv0E3DSugFrR5fSPvzaRg7qihpXMR/oKMT
bBsvLjzWiWjdkVC4WFYb4GL07WQHuN0kSsfVL4NrmzF1uqIAgBDcFuqOOH6cAV3Fw1Y2VTmgMnfe
tJSVlVnod4cFnRODjAVCYJSHZH4EsFq4Vcm2G5L0H8LJtsYwGFFniS/Sd7rym/3Gbqojxf3dSKNa
WkkB8IQ/zSj8wDYeI8Veu1pBx19Nm7DTYsyjOjTgrFEfhrW/gyK+P6eNoc9cpkxix9gkmbLZHZ5D
NYsj/LyRKAyAzi6BDA1K8Hk1ylTNPjMlE1wiILBxlSqckC/dcw4mDszeBgizKjxWrPPegIW66KLQ
b/CDTO8/vOPDTzyfH9JFwA6tp646NaqCWRmtC73LACFUTQPQrmJHRAlRYnfI19fbPHDCJ4MGfuNJ
NBlzdTTLRu6JueXGEW60BtZUnMG+3ZSya0SjXWjV90NBaJ6Wi76NFBYlOOGEEw3Q5TJO1iaCGJT4
acwdIcVOb7eKBqRNe+lT+ENbHCJ/kXb9xcMe6uXyqtXigM5zXWU2ikR8Ht8crqg3VTpaf6lw4qSP
0a6220InDQTCGc8CcO8NQZzl08yPCp+SKKAsSLecNyV6tGaiRhaZtPOEDigSRuTX+EJ+ekOkIZYT
jVKCajwWisZW4hQbgMxV6LOm4n7RxZoL6ZtjkzErV1X1UaHcAxLiT3XWOXDF6V+7U+5TmhArj4v7
oh+YJFF6NG0RyDQaUqTMPTdO5iDmpjkcIkvY/3JeeHKzkVFc2p3QJZNj0bT94kOMw2ky2Yp7eo1W
CtpP6xpniJRELKv2u+hJRPwT2tyQVMQlPxdJG1q8q+ePBnn4+AvnwlIh6wcOG404vAkpJhpRGlpR
FJWAEPrESH7OPuAQhcwnPKfU+9yfbpguJVEwouHLzEuSxAu/Dw0iGrTlDDe9SPScUaSLeS2Lx1KS
BU7k3OBosxg7I6X7Q7AZWV1U7ou52s4UHiAgEopcSe0qYgFSd0qxdQen8IejlAyG4qYU/HhZZ67N
XHGF/9JapBzGQILxUr+lNDI5S7VV9yBLz19BRN0kuW9YKWHk+wjSBKpAs/mrgKZt6JJYi4C5eLp2
G+iEjYUPN5duPEjL1cl8NsfY4F/M9wlPEP5vpsiVyxW7CgYUvo3/3O/cjN7QGe6Mz4fx8yo49vTH
PbzPgpzhMQfNq/IGpbDXmgHzU2HIMJL+jae/T8ZrFGDZuxPyh7kC+HEExyQWNbNUmoFCDv4yg7sl
ebAqZSXG8exgO0eF3t79r9NORDpB2ezVoh/dYJ9GaucHoZqYchcnR1ewM9KX8mpuOtaYumQ3NQAz
hGhOZwdoK6M7cpky1sDUrtx8FH/8PqlXGpGHiWRSjcZOQuwvY6laUv4NZhn2TW49mqOU7ddtBh6R
LcWtosQLPk89nu+rHpE1VZEENQPwtMcml04O/nCZnBssDgwua8eqBZAquL5ywHdx9uXMXNDd4Rm1
bwn3SpoT0pc48UJn/Jz2zC/xaMSEPKHTJ2PITtU+eB5pO/uvz3YfbcXn9ROdOYQS2eN3IuMj2nti
+T4D7l1a8PC0hLtgjHiJENRGV/9C/ga3WFfd0mlinQdTBoZ3kogWQiglBvOIczBDrEfOEVoY23u8
k+CQS/YeQmhmw+5j41p4b08KaaphKlVVkYc6s+WFJBMr3vYgwsIuGVjvfeqtu63LQSA5bVS8ZYbg
i2ZtM5b4mnPcHUkOCMSXGYo/oaGUMV7WYAH8/amGq6rJ3Rz+WSBntLO+B22vZg4zmGt8S1ZdbZH9
MJwKkScF7DxRq2xLjcpA4xZ2bCDklsomFfYzq57dG60lyPZ1NvcawdmpEGYnvkpdMzRwfyTs0l/v
u2LgWQxvcMzqobauetByNBK5SAIWZWQzZ0Wyw6TqXaxJTQVNxzdCBjC9mxlUAUAz9tSxZJpw/s4t
axDOw80nEZAtGxk6osfwIsh3WwTe0irYu4sJ9OlXfT6DyGu4rf0E1ySm3Tf2+kWGpm4dlI3iDwHB
2TGFJLf/Wnlbd0sKkCfJuclgNm5kVySv23LyBa6MD/RJKey1S2Wh2lq6XL7t+umvdlD/t/XedhDu
MN0sjDriPZwF90Re3HMkasHD4H/10NZEOu8XQUstAqVAh0ryebkP4Csndn+ehwzB2yowGJsiBIPY
swSSL2oMuy8RkAX5UssUMvSW9ksHgtpEmHH94naLkFTSZ1zvkHS7jwwxsYhZUTBEsimStcD7R24i
fyxSXoXj6kv6EZ4OU+xEmRJodB7qqVZTSGjO+cI9Vss4Be0E+XU2m70KONqHY1G6nlldvEbsQNh5
k7mWGuRJWBh1HbsLViIHC11q3M53PHb7/zocHDpmox4Xihmn3L3sIpjufjAvMOBU3kwSTaObFg5v
IhcZHVqF6fdXnFFA5P+vfobjIeHQoHJ4Kx3gEj0Wrp1BscdH4R3UR1XdFTfCof85Wk6xxKjkVxy1
LfbuXHPJ9dvlp1l7zMTj5EZJAfe7tLCYij3JBd9TCZPMLUzW9GPO2MUgksyy3YaM8Baws9YVgHBm
DqP2tJ/kpv3E8Fg7768YB9us9MC9MS9IHKWIPG+udjaifBGsFicl3DDLy3cTjCzWSm4qqUiQFc1i
zubyC817zxBbT+3x1wihmcR1gAVZpn/0zFSLTrCAFywFpPbL8+2NDRRa5eHTk0w5kwzAe4WAQ19M
06873KhBZVn4U0Qp19o2UGaL5CdGAwGgF3GPIoKQEm74kQOvdndD+YO4p4LfUJzjyu5liJZEKsLC
hla1jzi9Eg7k5QnajAmHvFp2ufTW2vnDicyMnaipUIIRgGj5M76qFA27kXYZf1OdXHUm75kpjsJ7
HQ2TprSaGZrqCvMb+kXfGfbMUw6/opsgaCjxFBF4L5opDOt0iJqyxtL0CKv2IsZbyOBwSgmSYjy3
oT9rtMA8/6yHIKXFf2LEHzrwcT7/wOJyht80OAH6hE0FMZbuVSZMlXHbYRwwFGGJH38B4SVByALJ
eQ7kQhi+be0aIUy3CVrN0rRDGDyaNMdPt9SMsNezMC8+duCGla1WIUBZ1ROP2vTwkNSZ5NftFP+s
8m+3BU7mVIoESr763i1RwrYsoNeR+rEJR1s2cNNmRmTck8WOfFitjQPAQlqyeD70LJbwr1sL4cED
MiD0+4yFLsj0Xq78p9DEBSxaq7q9HVsYeAE3xAv7Dt2FRDRLa0OdcmCrtQQtf+K6i3723R55Vfds
NmIw2wQ8jnR7uebUhz5rH29uMXEXT0xVtfsys0jqYbSWAKHapFxEwmvcRytnFdJ5f8LtfQcVOvB+
URPpxTakWLRIwkeW3AL49Bbc4EA6JmhXLILs25Ny2ktuPoUkwppN9Von13sPtIFb6a9BZH8jZZVR
90rxRjzdIiVQHC/qAjTwkdUt6BLFmTK5z76+2HYyDBsLaJBpiVpq24V9d9MNofhSxFv9pQGVUZie
W7ijIhzjj4JSyYBImQiHoSSdji9m0FMIX7hzz87vb2zBfBN2q3gDy9XtD4hDS37HSZ4BKyPPHil7
BQI09rVULFf0KlxwZPASU/stUSlTaIOJzB/cQMUBcYJrfFI28R4Y7P8WSxjFtcqGWGfTdAxjofSu
reJU64WZVf/lwsH334hHQpuR70VW/i/2wCmQLx/HUT3zbuJ+BmHAjGqUGZmyWXu7MckdNVi/vr1R
n8U2H0GRDIiNkS5s3igiLHCuUSHiNK2riLuJpx7Q7jLZegY14WV64/yoHIR0koDzH0qtmovGQ9Gk
YMkU+oRL1el2piehXxqJNXCxST4qMJUP9VPm8onU0ljW4YpW7GrxKDCpeurCdapUTUhmZORND11z
aZe/dc33LsNcVPIJ4ingUIWYk9eaqmYhr/cT3TfBW5sYPNT0jF9QHHk80lqklYgxGX2Vdf8L1rHF
RULvNyQ5rrASG/RZ1SN9z8N2LLx/y1uSHttvClsf5xqXj+4sVwTSkmRu1/dWW5xOF4f5nl2/LmLA
iYHj2cssaLOwBDE1PVUazmjUHp6b5qYOReYIiLqikRMH9msNJezqvbaiiGP9K1TwxHi72zKbMXeb
mdSCKxTwQZk/ccy+EmLetWzG8wqI3hX6nuYGtEylVh+QEeHdDA+lyxdFf3kGCLLig8xvWG4dVruT
gxey7RM6PY9sTePc8pLkqvnTPbxMn66lcPo7m9bhmJ1lUd2XLgABNaaZlJ+fXGD68PlC5oo2Nw4P
k2h0MIK33huSFnE9pTB6CJr22LVqZDntMb9FYmzmb991gKfZBtcDy4r9nY7rEL/neIZFkiyqeU0+
cxx5+05j8dmnEdu2uPWakBj63SomWgRJ1BO9tXMjmRZZXjTHUo/bIjLhCXoH13YKZjDM3EwjrJSL
1okdFbpbsfd4i23hlegVnVsYUkelA9J9gt8n8WvTRKtD1ldh1mawu0Zk0n4U/osW3NgyTdEL4DTT
9GjxxUTtNJipXtPZKq8KAVv5eDM2+fg1Ga50tddad/UTZVBN8AdVEdD7t6crbRJcfFMaXsIoBvfW
yp0J1d5aTO43Stna4+VJgdyQe9DBCa/XUnpLQAlp/tQoqXsJIPr4FpZylUYDydhoTWp/DmZ3DKM2
YF8d5C5HjyePUPr9h8aC4hJkCd3xaF7Ccued4LWfxgQi83ZQqUdXsg064SfBr5AzgPxwqgY39M6P
WKzw/PzDj3P5UoXDLImCRkcYp0varQmSNVCa2nHv/W9KcudYQCTRrvduNYKjw0mgeF7+SrwfXFlH
rGsCgYuTItWcqW4lxMWSqnlnsCgOq9WiKjAhM01GClSgOO5krHNklCpkDsgWTIp4nSUi6cwa4OZD
XXdEXFHtkUR+8g0yZqNDtYfLS2UG3DpKyYdUR8dmDFxdxbi0qF5AzwxXTh5HVy7dgx84/QhFYXnn
viSyYceH6kvuZWVFamkqMMN0jap3j+SVnbNLxvDt4xQCtykuU5lIp9FUVZsYRFc0yMBhKqgbJo/2
pKNKJt7salEbKniNxEXxJCkdtYjzcQIaRZX0Km/JkH0O5Uwv038NAbd4ekN+SSjQMi95dd0WTZds
/x+x0MHjKqq0YLqwhbsP4xVIC5qPccivFR2FHrAtfCzHR206nxoftN09pxZUiSjF/1UqmuMXtlDD
MDUeMkJb0Y3EAIeSEWkwn5+w6d0y1JgrTXQPloSZARoP0+Hmk07Ox10PcbuKdsl5rCG/yIAaejji
+FllLFkC/JdBNFxoEz/Pw97g3GFCuRuzcqVnsFwvctLfczlNHpyoT5XcytrZbDXlp5FSs8VWYtzS
f3QHxg0F7b62mSg7Lnhe2JJkr9QuoUj9GZ+QD+hY+ut7mPSxR2yw+CwPVLe9XhgrbKh8q+pEYubj
y6OkTQ9fqtho9A9ECeBmg3RS4Jz9hl724k2Sa7DNO9Im9gzKkY3DuxFh8U1nsrjvMS6GPhK/zXws
GIheotEql6raTlb1J0fEXBT9XQmhbGWmAFSsxcJ8TKqymwNWKiDOSVBOw/44w+C6UoDJYzDlcV7e
YovWYmHz2f2NnDrAoRnEXEqnD2hEp1dgMJke8tpG9XBDeqorAgqzbIgTLLjX2vohmVUbPveyye+n
a5WCKFCQO3gvR8JEoBAPH2aNs6bxwyft56OQeFiFytCfB4ixVAAssqja9DJejqkLq1twOOVtmhU2
VlPaCIu3jDmOIZQb7Zlca7kvsqlQKVdgeLQ/JeW0MMJc0E6mcUEJ40PqUibiZU8+/L7vY0jv1tz+
vGrgjzMS+m+IbbLXpSuC/Pyuyoo65YTs3kfn8eXofTnpLsAS2m61SbKNRX6w0ENHV8cj1ysy3cZa
JmZ+ut0Avi9WU6E5YwR08tyhwnepNg3u+wrHXawpeOp6kwCdEH0+qEEvG6bEt/t/Wfu6lE1T8Lz3
WkHSMxGa/bdeIDBBAwhN1PE8CYHVBm71qxOD16CBhZ3k9HjUf2VS+WlcE55vFjU61ze1TlIucqdE
2qBGFATamwPdtPTIXEOD7WmDPxjoI4g/z+BM0ph9e2qUIpn0TJGQ5k32XbIGBM4grQ18n6OXx5Qa
zavkQtjgkEg+v0qmOQtZeYe1rE06HOEulQe/0X98XE8/lqfqozrOgWuPuVrGz0j6ebJmAEvOb1M3
gvRydX9T+p+joJTB/S9tqJ9m3kR+TS0dRQbhhoZ6QWTMd446Sqtc/imMRUL06URWqXVss3myphqw
3yPqRAUIm2qjEA5u228uIEW9nTk6HmABCma4+w2Qu2XaDw9OKPACXac9io4TbmvuJQLnfxWG95ow
dThWnElKK94j8mlh1ZilecoszoVxFDaz5BtnXTUFBixSV/zkzzbzvyFsiPGpnzSRuriCouaq6vRf
3/mc7dIJEc8AeJuvqWdYtdfrFmRrkHW+8tkH04jtze+UNDUqlSmlm1G5sqmR5P5KcWQRqpBa3Otl
7HM+CJ/9jzcetsCSOffDOzZMn5y/pfDiU6jNSc34NMSokim/Vp6/CaSi6fvCIKAsPY/1wda0hXCP
Gg8mS1a6A2OTFXSgrIPGU2KgeP4LULziPH1EPlsTy2wSVCclqYEaa5EPKb9TTWIQxrP9VIxW8WIX
O1qkZOqFF78IqX8gFZHHQmb0wgFBQmOwgm6ZSmSJ7Ykwqtaeyjf9E3cBW36hNXVaewJasOo40pch
GPc5j4PvQRJQDkQzYYSXhV4JO4ZhGeif/ybz1Aga2lUdFzmo5Qgz2c97hpK1K+xvJrO+edJwnjW7
dF5VWrvijM1qS+ywkNOSEZjEQGTqr7LKHK76XG2fzavz6SgdL1KixpnYChp+AAp2Oxj8GI03V9Ll
Pnr7INR25DjDmq9i7mChtM04NJeFyr3LDYirwsmlQs3BO4vmrwKpgBRFMshO+mRK1/YVp5KqvWIn
NShIwrJU4k4HO3GWsB4DTrHorwxUopzRiSxIgzc/6l1QFmfUScC7YoIpRgvYxm1Ohc/HsZmtUO7O
ggMLdSmY+raChKS8SiIxKVVOMWEUSDE1rtzUEeevmTqysDssetpjTcr6dsoTsHWpkcikfHNt58L4
qgw+hBT3h2klThcEBbd3Bo10VkPvyv2h9P3yoTqpuhYaOKrxgY2d3JDNeqElM6Zarmh5xBPlX847
UEheL5N10XagnIDsBq69vYN26Xz1d2j4rPaBDpQOqedmVU2uUOIwMQXg6LiJFwshITyhnfGCLYPQ
BzWryH2aDwDeGkIM4586CFCWJf+KhHTI+e5VnmZkoAcfdBLHu1+ClLt/UpXOPVRQEANVf4QfK4uG
awpbH+7kb1wuKB2c6qy4q9WtP6YrwgOlfI1uVwwQPKdWu8FOMddHVgBENH3hKoOuZQb3BQm/S2Yg
hIabi3zJ83OD3uEMaH+3yxxb8jyWIII/kHrPUUk4/lUZxjEzdwsId3ZiGFq6nx4IQESuPh+SoZtG
3TEQcQc/M1lWQM4mKfkbbxlEeCxPsyjnNEPlM6KBSXj3dtDGGZae3FJNh8+3nnGdLLYWkB0ptqDb
9k7C812Bxw80y3Ex0XKRYtVQ2y+/AYkNt52ZrTUihXWPa8x63MfethqB6VS/eTqS+maCbrFkk8Ps
a2rEb1iJk7i3crJTIaUdSJoo4i7n2Cgc2v4H9YiSC9Dc9Lr5M5XUM6tPbSfJGnSoWuxKAi/3lcPb
qv9a7qHFyVrg3XEGzz+zgdBExIcmTVzPEd1BYXpZDDe2jfV0Gs7YAcElbOPGzxT6UTzJ0sgBumjw
YtnU4Uebi6F4eLiW2mieRzdHqej4yNdhj2srYYblZ0tmNqIHASxznJVphQ8sjglF5Tvf89UWd6Ii
SCAywSF9Eq1CqKXlA1oCKrts6sSbsakQ2WXkVSK8OoY8/uunZRpiv4Yscv/CqPvaW5HhXx14MlSx
ye/uX6x02N8bk8dK23kdniAXyQe6aMQSSQWID1BLF1yi64+xKVgl4kaUVuJTFZlA4CX53oI8tVVc
wVxLrr0oladv694iYpoCl7hugz4ghX43zN3WPjSfXEpcAkCXOD5kg8O/TKhSMcye08L1axB9BMNU
lifAUTp0Fc13Mpj9Nimq31SejkhWK4IzBMa0Uco62R4BwIg1mHXtTeJZXowpt7MLAYVz6cWPKUl3
IvUbiH2PIbrnFgX9WkB6FzsLtCg07J83eyJgY7UHVoKKPsvH5h4SrksZYtymlvWoQ9/d35vtEqJ8
wL9CRBNaPsGe7NTk6ZLbWFwGe9B2qH5Ac9QrDZpFyU3WkAcMPhpTXenlTrVdieDaBsRn9TByUb1d
2+zqh1OLKt51J8gZp4NPIMTRw1QgSBp6m6mmBObISWCuT/KP91Z8WMtl4btIFYaH49u0jXNEpnO+
qBYb6NnGVa6ZglZVFYD+vXnbYmYtbRWa+P9pFVmD7ORQHzknNVtLoCZ5pHhHdRyLrMg0UfMp8Ye8
wDL2QKds9DcJT/aMbSwikrf1F+PAqO+GAar0X8oJDTJOx43SrBKeYC8bntDZuK6YOmcb8WuBbKK4
1LHGLG/OkDi5MRIP8EMG2qboveUg4xHB/fXIH9DdYmTYK2JHjo/hCtrsLOz0iAqz/884UyTQF66c
S5RYNxlTKkWgeXCDK2jAVmnwXmAgVtIj97dxN8RX91i+/gM1rw0iAo3D3xGEI1ysAByFH6BLBpnR
2RKzgeCWrmYfxFAFXWjBKQKPV+ASPQFg5qp63JH3yJWaOFK7cooqOYKB9X2HBoF3ZTqtFh8CgaHs
a1oYwmw0+l1hpiba6xzzUSs98nXWLY71gJQSlM6OqGXIiu1rLAcd0UN1TodACG19i0sPEXcPa/Dj
rjxMbL6aP65Hk6jHZ/SHwxmS4zm64u/6JtSge9XRKcX12owArMomw3+jH8ORVWdBjo15HqkiohXU
t8S3US/ykfpM/koUGFaZtHsRZ/VE8HCj6tvtUM5wla4/dit/t3QEWxxICXK8kA9HBmSpSBs/ardQ
H3iTM7lnbQyl+RDb9n8Uvp4FV6nknpJL10QcT5Z2rSRBoZXjYPxwa/QmSzjRYmMoqIE1aITaA0i2
pDMVqyCPbJRivBQivik8v+r36Nqfh9CsBXiZ1awcarhkYVzR18sf5cRkV0SBmUuDYDHpW5hYVbAy
2Tdj9jbJSQ/QMzqlTZfV20fof6kgbYi8EAqkOJJfZyrOjeK8qh8ojm71ZVLcEScJNrRe0NpOls7q
+1Y5reVJ+N4lpeirZug/5iTN9AUkty/bdl4Xa1tJdsTR5VWNLB3LsarLptR0+Fl9D0X4QZhBi2cd
xWLPktS9DLT5RlDHXy3Vk+gJkzqNnusNIdjmr38os2hKZS30SoVeymxPzkkzgut9MtlDFKFzrzpY
8r5DRWxcK37pmWVwInyuUfUhgIiYXEsrocH0QszWpPzHWYyo1aTMXbcpJGwuISww8RcK27fRkszC
oxdt/tGZTPKZy/3Fv6CHcH16ymfC1e+H83NQvexF2RLJH5/REox2wAdeDX8M1x151nZ6Uhk1/UQL
nVld6qSIEh+LDTyxFZf3GTvrSPwzY79p7dqMm01xhKOszAHL65kVcyzpUVGr1N5lWRxX4R12j/Nb
DInWtLiBvHAb0mdjD0uMXnxNiQSUYnHcylkuhvyLGlRP09BQCvzcPvFMQlV64EEcME5dkNL+7XXK
UhEcVSGVZsHmCy+coXIPi9bBtXhg5XfG/lEFMDFI9IuUBocJcUjLUjzZwggJkJh3miePFb0a+hxx
+qonr6/YjKMUKvJRsZvRdShXujEx5PNzxkAibF8HBNK/+w1ZShz/6V+/aFpXuJ1YFVo9wBtGp2s1
D/GiHe/J+F4vOW6WTp5h/KrX0sAsyO80lj2KitGqjdcPQ+dv6r0hEOJ3X3TZ+Hb7mmoTGUIjlXiH
9uqpnid2AriHg6//so1KaYfhCtpABnegGWSTi16H87aeN8rcw4h2qmei//07iy8dA51/RZUFuyBF
qdQlwWgOz6jN9LqEhagrlw/3kcVgXrA+Tp9+m4TetyY2IYGml9x/gKziWVnCZTs0OVzmFH7EqMVi
6AoKIOH4F/jr75vxuqpm9qlP0150J27gbzPG0419Fd6deoyqSzjeqWWupmo3vQtU3ZllMNM8eY98
pXNC1G6kFat0XOKzxqM4zyni5DFC+FyeSVXPsZ/UbSdJrXW3xxHRrJZN5DO5LzGMj6xzfvbikdjm
pOi4J7Q9iZL5FRZwjKZT/3VCqlbO4zeFnHuC9bzK2uS7FxU3Z54T56G8LSiT2kj+lLxG3bjen2kL
uoYOdolbj5rkF4t9RJQjWByXaU9nJN3G9nS7hHdFTAOdM/vg/sOuXl+oila4u6mvRt8xII+Ru0jP
qhz5XCV/NUGqhSQ4pNNKvijzXgP+34EcDlHwymQK66+NRlQ0k8OL8aE9yuzamt0W1KT60FVNv4Ga
ardU/2/b4qEojLC68lvmwD7BoHBOXsU7chYkLxMy9eC0RnqY9yJi8Iltb5NMdVVhGJe7raLXqIN5
0e/2AHeDB3I6YkkB4e8IVyPE9awwAwQKJQUG5PnoR1W02N5hGP5QuKfBD/LhbNmLgQvxjnNTCTMN
XjTwPtAGbAtHgBF+Hx7JWY/wZ/wDn9y1W6BAo8909E7zoDA1ZmPYYlkZcCf0dYBfyb/4YxVMCIEI
NnhyoUQ+O6kvXNrPlR32D5JHyflNvnD0AxGueWwGs9HBcHQ85hzDTzjeK/fyvbgzYKekUPv37ISN
qMpUqtoeUXp2rEgBu4rYNqbWxB5gTJ2If//JLXnA2qGeNmU5mjpZe5cKn5L5A45j6YsbSWnz8ABm
2tqP/r8WDdJtBAoh+Ub1mwMA/1fRHbwvTS5/HtmxIoenaxBd1Arr1AYvcfFF7EjxAG3gtS4UiuMv
xyXMg6CuLO1WbB0hwbXNX2SnOJyXRlmXwDsbdVTN+JbE9oQGNeHo33OL1mFbypP6dvl+EZLA5YyR
xvlKiGKmE6PWOaEJCzbWruQ0E5OKE1CA5CCWwX9lffBzRm3yNKKDGEAsl5Gq8lbtzqTeq0tJsxZE
stAccYBAiSoqP3g4Dm3nVAw3ctWZBMoHO2dQkQHmbBB0GWn2jg+g8wE4YdNtRjblRKirhpdRpX8h
3vD/Fwn8lGzck8MsmUsk6J+UnMvQy2lXB5eLL0Mu5o6zK1hYg9bERF3LZaN9TNI6SNA6A6OMHcYq
zDSXsoC1H5PElye4/e3R3TKDIOsXaa2kkw+dAXXwJ2rUUQg/aZbBn0IlMNy5jh0Zbe5KpzbFwT4X
Gviraw33k3vAdBh1FfRLU3LqQwm5T0Q2V20R+kqVm+c7JPLIVxQ+mXssEPZ6JTkd+8uufOrsszat
0ZqALvhPK48gUUpQLp3BHWQ6+mp/LDSez8xp65ZIkm9ewOOBWPrYDsIYS0ma1a4EuAZlTJ9DTeB4
8BkFb5qQI8Y+9WF7MIeuOzC+mUSfzOdCbW6l3VIrDjZPLpMsgqLfjwkg6U4s3fd5VAeS26ylYIjs
SgVdAYCgweExy8IWKqKhv58GpE0n5d4HWgemEkW4WbOTLPs7F2mphuFM37vRJqQBY+yqrr8O6ypk
K7rhHuODViJm4pQhsacwlyXd3E82ZXraaDHj6wxijheDmRWvq75FpAUDfNtt53Q/YNfObrj70B1L
MU5NK8S7fBzxbASzb3Q3te/k0QkTBSoIrvTqBhmpsPjdf5LjYzMQ4xgxEGOIWVlwVxvk+VqjQwiT
YkHOldHdeoiqxTZAPKcxIdcR8zYZlwy3yDWKWDJKPolzLDS/MEnvxlmK3t86iegugITJPZfN7mT9
s8kX/beUIuYwd8wl4+6BAeTtihshEr8y6JVLNRVVxIc2UKq23NjNKH7cJz6PvKDNkIIcbGKqONl0
mkIzvETpQKSE4+gqb0j3IplC9knCSfo4ILh93tba4S91QdxGYcLeeZrgPy0/hmeEEKYG3n69AOKA
iZ9vUv8y3CtsrP6bhe4cimp94cROmfrACg1ZhEhhZuuCkF2+UIu8x+2dh9l4A3qp43dNtieisdhD
wS+fY26p1UOCI0rHivNY7qWCmnErKSSFxUa+8yRdpeIEnymaOjDzgnr7QLFVWH60lbl6E2xE16Wb
vZiOwf2iXZ4jVg9GiPon16Q9CEoTKqiHX/Mxt/3SZHPnyt21mEAlcE8MlsGvmFKOy0QAnhSHIPfz
W1Ms4/il87sK9sKDE3Z/8HTS6JKzIqzMrqqP9cpbLYVn/DDWP5WdR5cCpuiOU85qJ/SMKkZ/WgY3
gvTi8th8BSB7Qbxr40F1Zc4q3qIplIwO/G2jNcHygrzNYsKYgVf9YPQzODtAeWad40dSzeNUIaeb
MXDyO3A4DP1CpTY7b9gOcnWD4IyIqyk16FhZbYXlqMtGbs7yXKQ5tAN7WS+VAdypQm1Pq/bZBlvK
eN645PdXpoIUGryM70bhPBTywvZVfMx+kitWxFDolstM6OeUWX6woWD6ID21jEwn40BSGNLOoGNn
BOQbGFKhfrCtkSxmW7ouJYnsqcKxeRJIvlbfWauYjC0/baioU9aIPQRz+tf7Td1Zk74yHJhApR6J
YoDcEzBS3orrpS89bQ5wJiFa8UyWz2nFB2j4pOaUDRf4H7OxKWc0slL2HLIwL413zryth3KCKsJq
FbE09HNA4ETibxwZHnzORnGE8fMeDCZcfQCvbcwwEGV4HrUV/sUWaXGCuaLCYqQ87/F7E3xE/a3h
AzwlOlop86gApDH3JVYr0t52kvlqFyQG6EsCtSHbWXV8PvTje1Fm5QTHdhliHxdHqVYJNZkEJGKF
2l64E1KVNmOO3aK/1yMfNVosHUYnpmyzUfB/bzkitoaExGC60F4ORODSt34zjlj3pdAsDFIAx0PQ
CTvjMllzZLA7DewOc+QLqRK6mIMH4McCkzcGiy6OJAShPKD3yk6rNJ2sRxtdPWrhBgAlgeV/feEY
QXEFwZ+tpUrVhVSOmNgCapIPz0T2abt33Smmp0Rqd/WX213BvVPip2q/Y86LNnfo7z4PhU5jqd+8
z4J0nZqmbaFMkPepeYo+9DgkS0fDyMXKmmbr5apmzsggxt0rdC3WHrK+wj4pVdrmyzoFHvpX1KG8
IXYQ+V1Qc915/HiMqoZlxaqx/565UShs+yZ7Ie3ImVReQam0myBm0dkR5QUgHMRxFL5HUKiEGKEn
skAgKRkhhA8xIEKN9b2gjyYDDPRRugj5duh8YzD5g6MZHUThEWGE1OrlK0QHhVZD3tgAsJyP6sTS
G7qid8s9mHJsQ7hiRY7Wz9bw7KiU87NJVk98KVe93/9h+uRIPQ7gEbvcLb0Y5vCQM2TDZbRb90aR
XO2YVBWE9GTYn4A9E8urXBY6tWC+4OfD0feVf6JXIYmkuP34Id9gAcP4trclyBG1o1V8cjw6Fmf4
Ps0PZYNQJbdyqznRca0DOklR0HXZTlBP2KuJVOk15apg2GtgugFTI0yC+78tY9jpH8bv705nTGpE
ctRPkCP9TtTd+E5pqvw2ZsgpaJAITTBBog8dM86imLmlvZQeihnPkr3TnT3KMxfe5CcoImbHWINr
4B3pCLFGes/TOP9yIwrBoYpjR/WvrVg53fdEY7fgOg4uDYQ65Hgj3IPWpeNYncM02gWD6BUhg1NP
/QAne6qsn4aWfCRwCkV/WqYSU7pXwrYAAfSLjd4jqQSwnwuHvDw+OhGcaMFp1IwGyG0SVn01t27Z
GiwhWQqp1qBM0gYu9tT8U6IviDyCQ9Q/Eik8e0Cwiw8oarKUNQvoL3H077AfDn0er+LV5HdVcr+L
0X+2kmKz33DRkQvJwJZ3CxcTG3/ZGJeNHRkVKo3n4hC5/synfx4nhevPNUdkoPriokDgt7d3YVSe
PQay2NLVlFLqt/DTX0CPkuIBe1Ps/ZHf4A/wrFLVSdidmdcwkJiny9+Lvtuq3JNYnXUwQak6+OG9
KEuL1q8kmWVwHwSuiX8t5lFTGy3mKZ80VG09VIuV0DxJfAP7Fn8Pu8HWi3t1UGWZI2K2SpaR/IGk
LvprncEcaEK9HDkINxAKHairkh6BZsllBDoY3aAAS79ImjNPe+fIJtUPJDYSPIWKEvm4kmG8sj2h
PM/XS6QaHXudeZ05pjce6OAunTPomaLFOAPGhSh/iWpk21KcAaaM1N0TlGouq5F+S1lV6oIzqOaW
Quq8c6JQ7EMRzzJyK8iQogewzuvkGyWisXM/zMHrOIdfvEH/Mkbbv3WDN/zpfw0nXAggDoG12Itl
WpVIEzG/3IvfO1WoErZrC6qgHeF9NbgwJxr5G3HamwiK813sRv39uHvIQ2DXt/v0Wn2SII+Sqmdn
/EZhBtXn+Dpu4iI4wdoOhy4T5thERSbPH3aZZXfwT2YUNIM3X/fM8yoaapbySWnJmqTZEuaE0ud/
ma7ZGXI3OKf+vJ+gbpwZideKXSoA4Z69yLvTggd6eOTvEOC4yQjSpLS23BmBy3GmCDiQFfWPdgV6
PHBQ54ksoxkp6DZdxI+hLkqHiy8PaWeblMtH6IdK8hg04TAWDUYtex+xFMKKCOfnuukjKdNAmyl9
kombL+yk4nNUNLRUU4PKJ87/IATzIoK+9DqfLJFztJ85faDiWQgA8MoHi+EIeUGnuZv29g+8ExMi
/MXX7UxhAWb5P95+yxtXE2zDFggXYAONP5OJfu13AWSMulNuB1bEqQGBpCCmdiCNxqG6ikP0qKFt
DG2ra1pQm6LpiNfDBHIrkPbflHxHHmYeINp5zjayE9qHybHKo5HBlS3b9GduVWuMfX6M1slV2Aai
ArdltNuFqpkn8QSvkSyhz7m3onczI7IIUL4ZKu7ZFYX9lR59SKpxaBOet0v+Rij0nynCkkTAlvR6
uBZB3Dr1pjE7T38fyWkOosQmMl4VKncNCguL1w64BAC+2QaINqI5ohSvovrxT2mzMKkgan0GASqU
tmfSa/vX+K55yPba4krDfQsF4eUa5n4TLz6LzC6xoDb0hYo7f9jGj7r84yvJDhX7h/0u4fXxjijQ
T29cqgP8EEdcitkRs/rVrkHHtwll8d0ytCkLANvB4gRROQvcONc0LLp+oR2UdIK9GxSa1juNEsnw
RVyf+u9HFAwcAhgg9c/cXqESC5WWSp1dtMIKbcEQpCyRgRRiNEZwn0mNueYosOM3jd03pS1yfSAA
Ap7S2ZOZYPdJ4uvcUTUOD4W9Xr6Zq0E6L3JhKLtOApdfm6HV2sIqZwbPOSHfqlu11dqgEc2fiY7y
I25ZR1bvcCOCe7upr5C6E5z1ceX7B1yNG7ax53DW0skFuyoqSUADS0l/6q/Z/gH9P/1Xn8Swr8/c
nDqQ89alJ8HqrrxrBUSdvcjiaI3N41Jo59jyQVQUzjMGc81YfNGyR8aj3SaKtBfVyyK9pJ3hokQ1
u7R+eiefJ+WNOkktd/dre+W3N372/qdzvLvRGyG/nZCuCgXeQ+75+RS149Mtga7AHDeZDNfVx0Gm
3wqrUDxPWHW4aYgAVKtqT5P/+yooOodOJovUvcwdT/Ft5ISy00+XhY8hG08vN15iFsopoXVF6kVX
mZW7Viv4/31Zt3S14yeqn6gybKbkM2RCJmg5hq7odcKMKyt93BjGOf64vMzsr/cnTQjsm2UHvtR4
mJWuCMtq2HjMNkTNoGpqBJhllc8yTmA1mDopG6MRIGl2YzB7jZAEyGGXhBpPML4ffOZtYwWDaWwX
PUto6dwh7ApWJTB+PfXaIWREPPJV/QW+Saxln8NEy0KAd26l6gORZ3XSV/MY3ePwKHacyAUYUFVT
WVotNCVJwtT33MmFJ7Pc1xXD+eG8mrIYL2zNOtrm6m6CAQsvSGaWPA0TVEygeckcxi3sz3PMkYDA
cLN4TrPeb0If83j7g2NC523gyBUqShU2CNkhUPhzw5jPgy7M/RqhU1HndCRe6vIPm8H71hzAgbUf
w8kIAfcY6dN3CaPBbUV2gpIV8I9t/dax/5ntMRYMSvDmQsACISWuRGlgmvj/AJ7jdzRjUezW5YXs
5KrjCNP1ezkcLcBYwRRyIB+9PAW75iOdKiq5CdDQiFtMSLhLXJag1CL2h9667tbWmQURk7occXod
/H6W2OgINUeE4SjAPKyYn9bAJmYzLOofsQk3xoCI5pVp6Sjq+Xk8iogBfundXQG+Fe6Z9gOA3ZNX
UIUMQXSaqur3hkp/wquYqtHCpibc7oZ+oFyZKX4ZXNmbvbFLHeamneus4dZYc4oVI08pgo7J1eTG
kBeR8x8ruA4RLgnRCLsBGSkUpEnjbi2L1/d7A5ryB5cZuOCrSR/gPcAeipSoXbwvENc8JU3x/yix
i6cgc+9VzvZLv6b/IK4KksSCveaiJikuSbkmCkSU+/u1DGv9jlrGOXkg0vDT/PVLv+hN+htzzQGY
PtW2tasWt1PnJBPzcYO19IG6mTZAnBBHMbHryGa3/HXJByS7w11CslUhruaoGg2MsCvYSiRR5kaX
cdShut1ddP+UHrYVY6/uc0KkpcVfYOKaskIt6abcfA8NIx18OlZbfE3V8VFP/P87Pt99/DTCZm9t
HVgp4rF2jRZR6yFDUbTdgpXM/VchOFafpIA9aGgcrrqqPVXn7rAGlcBX4ROSvNyEQRv9gNY5lRX5
d/xQc88fPrfDhleBYgPINT+iY1p38P+G94NQn7J8Ghxdw8GT6nWiPnHrtToy+wmpel/ZFn4VTHbZ
R/1XnUw7bdqwLzpgni9dNGkI/BwitT1DQuU0xpgEtGJjU7yQ6R2cqN7NRg9KP8gTFeE9pjsaH7s0
jqA61WAJc426bCAvOnjcHo00X+dA1G9v//Rdf7D/fpeevZUhR9vv7tqEWPdFGnBwQZ6bsAUv+QN6
i7cn4t3xWMJjtPE2ri3OPjPV/VguG+iBGWOriKrcwTLwuqSIIQ6RNIPaZsdkPhSIO9yF16Tka3eJ
PFcFMfjfXgYr37WmmY67HF+I9lKBs1lu2SjI0MZHn1dMKrenZz/oWH40g386oSPd4dtabb53KJT/
PIICpatZiJaYZ939/CS0DNAveGe5MiROqhOf1jl/yj2+3vFOSuiclsrWw85G3ZcCzJlSEwL+X2BX
kLZUy73P+8I4jpUENtkEtlLfyCFBTEThjMQwfdo25IsBlgCvrYKMZ+dTEpekvC39TsJbDWwHqTp6
biBxn9JBIIZktm3Gk3WCbE3gaoIzoELVEuJO6Ddl7oOQMbTXdYybUrAeoWoqv3sRIkEfptSlBivN
biZnaMvALQFwbG/+JF8ewGhrcjkCxcloXqJwvb6FwkSYYWLvbi7ZyvFVSpYtAmyrjO7vYQHjARHv
rkB6dCPY6yFRsLnhkx5VENDT1iYJNzgtA1tdKkK82LJRLlVmaLxBnfCEn2oe++UTGFjzBoqLXotj
LZDINiz5NYnTWNr2557PTpzwkRwX3+R6I9DpDzotN7H10FalEQ8JKrnV8gpz6XNip2NBrDiE862Y
86jZYLbEokBrQXhPz9xkKmTLzn2AWUaVNR38fI6/3XajO0eaw3aPkX8GA9gD9ZKDhxCDVzSnxJWD
DHrk8cZXca4EEqH6Hpc744u8fyu6k3Ybl4tA3c9vgSwEpn0dUyvb4BJegJ57mj+6vqHyNUOXnQDS
02NEfnG+Bo0GqtyC+BbaPj1x5ElkYLvGDNxE6OI5KbYD0fuOyL/OceFRq1u1J8iXMLUh8XX8FJpn
MnJX5HwenDCJ56zGIQuohoWVir60hjq+2NpqJ9LeR1P44257DgSmia4oEzBKcXkcsCXUmJEQ9TYa
ac8mLcKLmI2sIxU3a602pwKurC0r/xDYQN5zOpABxr0lbim/gXzvMTt5BCbSKFhVq4354m5vpaqr
qufmMvXhI1JKTi1ExOSl5h1uuyRtH43dpVeYSYfeuXIIEJooY4B3XtIzdNvmxwrNTC9txFaQuV6s
R+lbapWO/S8L9Jp5sgXVQlgYw95Ji8A/G5o7GzSJgdO3cHPUvPs/CYbykuVORdSCDLVZP+CTWXxZ
q7Ag7K1Mlf+GLMDkzKMaVN0TJQDpjx68NfxYeYlkWs+j5/1XezMhIGB+czXj6hx12CplMatedagg
OFL7PUe1SAKn4aVc7gmfb5EQVmqoNGU73I2sSc7Qv939c1HwRnpS1bRZsirc/MrvjPdSn9gaPvID
dmqyZ/xHEdQKZD1qHMQuBxPXOKigZHnXgZiE+O4ksbdoLMEZu9Wv1sDIKLHvDCCLiLoegmDGpRam
dJLM4b5HAtGCpA/zFHi2P1zZlFGM3L8i2qJcU8BgX5HdBNb93kAJuq4HKOZRrN9Po/Z5hpokaTzz
+HgZUEQjnJYmzSoI2apTlTY76esmDSO+7ZCopVrnC7Q1DlJWh0+LN/1El8TvhPpEU7Gorq3zqmLf
KM0eFNqcfCyWu6edZi3fSztL6G5LBWVENL71mRZ4RcsCN9pe5MmnV1+eT4jKO4ak2jMtVh0ofadd
VdCAkoa+9ZzprU7Sz4qO4UTu3MZtofyDQNRsnrjcxfgsRsvMzC+mQbxqo9apTbYEzUm9BqBepNoR
8xAAYlRi8DSeSGeAV4bjXO2XO9Bzi5lzDRQFw6HKLzHwbpXTAZiSpoobNnR5NQwCBMLlrcWdidw3
inyqRpSscjbeDsL2zvENlSvfnsq9FVY9LKrTfh4z+52NA1vwa3ZiQCOl4qmMjzrgY/AGulA3/9gR
CNijOycuLlnTd0wCaby831FWFoTEeaOulNzHBd3EzM6hGssmOWdlKRxRlEZZzS5KybDjIRn/GTVt
XL40tZaQT1UfIkiRyxIskfoQD9CLUKD7rTmy4aXroYocZtL+QA8+zzI8IsQFnKtzFXD0J3omIwfQ
6M/DGcIZdJd8PyuIiDmcCnVWMrNxnLOrZaZEVdHBCoqCENX4du5pC8KsVdU0onjkKd5lukOuh45C
AlEwNUV4AHDb5X67xg7ff+QvfPwRkuiK0XdEciosd7+BuEDaVliBbf7aUc1j/NyOdxhbFZgMYQ7T
X8KV84lKaWkPjB8AEDFyssfYDJyfX0q2rjQKEiOQU2QYWas7MJXrATAx2Ar068WvmHz+id5bffTZ
lcPyFuq1D18/HixkBmXlhoAWX/J2vbyaNLDfitcehiTx2RYhhsIScS3t3JvBHoiRucyshZgb0qaV
pokm82yUDgCi3r3d0xpTFpMO6T3I+ojv93LI5nnWUD7BYWaU6Y+uIsuL68fg1cgQQTu1SgPKHFW7
mNnf+kbP3gO64ofzXgN3OTzNP8EXsUgYw7mrjKOeHzfKLWBwGnzEii1LNF7t9rnjNsKOYns8Vc9/
hqSiLUsz5OIJE53ioc7BQfWtV17dTbJgC6UkXi/ng3hVZS6W/GHde0qbXF0kxK2I0or74bHehUd3
TkfG6fWsSJrB8pu7cfA3ldp+qqOFC0OdcyUQXIQKxRMTywtZjjH4V8/pLr6ZDXFsewnCHPjVqzi8
ZoTZjaCaW3xNh28x8ZsVQdiLuKs4EedA1XovAg7OGNKnxUOKtRbJ1b7LnaOz8/LEFd9eJx6BcYEN
+SNwGOKqcbrirIOeQYwzNg7eWud0wgMkZoINkts2qpIIX13EgVcb6BapnrStuhaVnV+oVC8OEP/7
nx1tTrO0S1cp8HLoRJzzhRxN/FOgSUH25I0x+2MwdAMd/fBAJbAm3DILLkZdDwslmY0Chqc5Nv5j
PoLAAePCbTNpLuyjakGBcDBtymD+nR6cfFISVm78Y97hDBzgJhakA01pTjjh8SEhiB0GmncezPeq
KpN+CakSYW73TD7LtG+NQ0guP6n2ggRX1RJGZlORjzuO/vX/3G30QmbcEhVeKyf5OZE0J5c6Kr71
BFsG6rhL/ZY9RjV2GvISoR/q69LgFOSYxR5FLueBmBpmnaxMdaQf7MqtBkHbAHNW8XWxx4L1Oiu7
43JpB6nmYqE01YMUIaSwG3x5Vp27eKDVlFEL4Jz9bqmMwycdJ/dZ8VztTuknteLxAepUnbzWoEpP
Ym1MoKAqOWrxle1UeM7KjRDpld9Cao5ArUHTidYROrSMX6FxQl5V9bx04q5u9RYzm+ZdJQIK1rwO
7aIL8RjUBCeil/SYU0WPPTKOe8FZacTnezPHh7vuj9HnY7ozUPMfFnGpH3HGzyOxrQ9p1WRvNTqR
lzzRVAUkWb733CaHXtfvB8zsACypW6msrELYfW4mOuuhH+xsAdl6wNZf4TaUBHrpQUWbekctUS8H
0RXNty1nl4ILf+eDSqRVIXP4KyLftjjVyJXzr+ONgZ9vvzPaSm3haHY5UDhaaOP2urdKOUZ4rNnb
aLG6BGaagjWolofZk7p2iTj+KunBSE98fKvfFP7RQXKDh69x1KOyYXmQIo/2hH7aAg6HN21z6Iua
AsoJ/QkV5NNdDGIyZrDiS4hdJH58j6N6Yhz4AVCH4lQr36lY0xiduKuSxNODxq4+CbyVvq54ZhFR
+qbls7EOT01u0gxo7LqHaaeq5IuG4E9pPbp1mRhhsiMSNoB+2xo+nlJ2jkmD0WJ7iu6ZazS+8g3Q
V1PTqKr995zsFiWNYYnbQJWDg2LsFnLS804AFXGWYFd9XVPLF1jurI6o1OBTgzplnHldONE1uBjc
s0kGBjI4qoyc21NJ+5TjJfQGn4mQwvUx6tfOb0GZok0ITAKj5jK3hPpYCUbnUqCkmZ1MxNIf9TrE
3uTt20CBrzkcehShX/IIfyThzPLWYmkwjeiIUmmcxvZOMWxtthinR3s/ZDotWJUwnp62O55BsoNc
a/EcKYKRS+JerquYyS0I8rqGxyBecusS6dVo3gy8S6cJM5g7SkcOCMdc3JCHw4dSezeg9SYODibY
HBFYMTI2dulefLJakYALWtrEOlO35/lV7XBfifov9RcDQUQP0vgBWTy4cODpKmUpv6V+cuoBjyVs
hmjodZyWqo7xxvIuSCUkyuOBWmiF+tDSu29/VONZESGTLuX8HGsDhN4iH9FvZ9i72hOLyfM0X9mp
skvmikRmqWKqrVgHxtw58xBp+OcEbcVN0MGaekIC9wrbrEpV4x/jKrNizQxucCEKtpxOlglf/lfi
da+BRfvrSeaovA8rg8io0Qa7oN0vsGnc2a7Uj8x3TC5cFeg1b+WXgDdJ0DfwME+dXvBo5aWCj2GS
f+Uk659NHUoKBrp2LeJQC3iiXqCEEwuEbxgafIObMVHNA26VHDuFfmJN1R6z3MzR0i/1rMP/BKg4
ImCl97mbuGsl4rbyO864k2J1h/8AKcyIpGz5W6laJXONnmCLcWD4YG9I5wE/6+i9hjRMav3pgsH4
5GGIYO0AiuFR4P/A0W8qmb/1Gx2+6/EXG+BrZHJQXZGxxSaIjZo4wNv1CVoj/4irCWXTpHqRslKK
5Eymxb/8Cg/FJAC2B4k8X780sPs5Dp8/T017lEEZDHLvQlAGZBHuUsbl9G7RdHZOp93fopDrNbxX
Tz+/6w+1wIQ345/2BnL85FSJTm9vy6Eo3V85sDozz3vLqc570p6bCZrBuuctBl08t9boiGiOawZB
O5mo+ATL3OCLxAhc/R9NiWLt5Glde0eQPdkZsj91E1rtNUvB9WkNTjxdh3aK62AIX2STWSL5rcFy
gXoVvpFg+4cCegv5Ka/70CZ3nuESjDlMYKtqEUnhCDLM/aAx7FJDzj64z6EH5k7GO5R6xqwVVKhU
r7d75pcQLgk94JglPIYwOIxg6mp3gSZFN1vwa3BBrP3iR8TCtMFrZEI6y7UPMlyZnWGtjNlE977M
vVJQP5fIoNyFwv30g5bGrgwL2/dv9DNnCzUWwZpuTw7GCf7ZyozWYfquwRgMLPYjsBttBmajPnLC
k5ORxwM1pQRcaVPpFn4/kMhCHB/urDLnUHpZaFWTATjWC3CDz6EPkoYhVtwcwhZKDiFzeALZVMkE
nLNkRHNpqijGk9QqT0fgv85+4bLiyccSx55A5oCWdaQs49crsbmJ7H6WTbP7WYPvl3TnMPuYr+v3
+dkAVJRIT9C3iERi0sTpmq4LHDBpwrEsKncAOUhueLskq4b9XP7bNlxl7lK/VCa/s7x2xLxSM+I6
yufUzwohYW8s519kbTsWzWY+KxNDlWIbR4kni8Y/DWkKIV7VWBWihAJrdQSGhwWZhsPgiad3+AeP
t6eWbYmPcnlfVEBHYCvSH38jqB3GD8I7VanG9Mnde+uU9FCKN7n1A4TWvf2U9xXKQBRvjVupBb3Y
4bKGy0liLkgMTrwUz2uwO1bcFVZYo1DSEv9wOQaCNoZuV05SSm+zmYxAk5FPzRB4zsAdYyXssdBM
UqgAlBy1Tyhrob8VVJwW3kMGFonPRx8zKieaBi3tptn6CovBtoNl6l+FN7AbSlXxgiDTFa7sQ3MS
O5hDkWuiZ6UdWMZD6zblHX2YeKabv7Ifid/Rl0jy5uLT468uThZ4VZnietv+1MsQIjSkRTFdfo+Z
1W+DD6KNT64Rj7C51/khcYpRDRj0Jla0cT+CfAc0bQSFllT20yTQ4tobacMEC6dv8IF3SVs1IXr7
J8DFNguwpkQS2x9T3UR6o1+ArSmCUYLVyulbYb3Qh2ak/aMya/umNQgkut0I2WKaIpbtHSlByolJ
8qzDzLMwLGetwVxJ0mCIL25HXvDjIckGM46AztKYhIfJrAeHmPTyydAP3arxH6pyN/sv0HlwS/98
SMkyVgxkeKvB6nHdIX89tAvUFRkBHzS4F5W9kiX89HnfN+Wy+bW9BaZv5s/K8SpeRlkoX0CEmJp+
TrDi6LzXgFTvsLiRXB77dFknpwWdiVng+yCmYJWLi6usBU2DCeDXvoewruFF41uDqQonQ9TQI59X
XurrfOWZvKkMXTzTuLnBkpcp4PIs3hvmogrdEFrkIyGiB/mVwGkiuqvuSBM6B6/nVvrUPDHvMvjA
XRwmOEkKHb4UXP/GiETwbJt6sFFaQnz6zyv3x+1SjAS7wEh/3fqJkJXorlSVnJSvfuVzl+2oj/w1
chwDDhm/vNMH1BrBHgGAVL2niWK4LF1YKxk57PhTixE1hmmfhgbsrxEAv4/4SjEtwe0tD4rOCLiN
osa71ietYvvdKL9vfDTyTXTtTLfPPmi9w2bumEUtDQz+9f2NLtoYd+PaoHn7ilqSRKKBrfrj1zMx
QJZa7l3WbSZns37T25K1MfEIAuVlDX/4lE2zRYOVGR7uABmjGNKoIARMXEcSQShzcYO91cgFqrYv
ya3QCxxFD/oaPsloQ2A9RTgSPyuwyim7d/InMnB7uDJjU6kdGErviGXyZcdrWih6C10bF66YtWKd
V1IssaDXr2dfUUTHatNa+sGnXJ/nuZVHJkxz/BlZ3+WR2F+/0pSAUIlmEmmtx6+Kz3E7glRFyhIv
PNXndc44bwSELGJqRrIl1tZSeU6Kekfz5JOVbiPB0Iz98yZoENV4ajFCqGffPGSucnhvMdVnBbNz
gn5Resj0irco185ISldnDHmLRiMOf0oMjeQSAMTFjlw7NSFZIcyqSKLfETiQPxzuRH2Ul36895VL
bqQ8DuLOSErEEH9nBmQYOyPvQpKct31xIFdrP+pqSJwaQGc0VTn04qkUkdHOlpma/lMxE3ewQOGJ
eTJLMBd4unOD/l++scLpiIzHhhVLAntWxsilKnm3p3D+dqeD/gWorXkFdcBI2UeQqv77iWZEVife
9zU+e/T2cF6Rrv1vIk+/kn9fA8XlIC8Da6G3/FMMcyAW5R2+B925i8lt0/EAfpvKmbdX1nW5oALy
mfcMU6YSxmHYP9gIwjUvhNPMDKj77rumL0DdhnmmKccBNAzH7Fxum76sWdWtKmiSMEKjD4YpbBz0
YmFDfo37FpM4qL6sDQ5PsfmvUx9Se7b9v6Q4XccvKtgCzQwq6AedKZ38JjPRm+Q1aZPcO+WaN142
1vluMnSkOmUvYKP2SU15BJNaQTsa307F6IARkLgtnkNTiEXplZ1OMQ5uXrNxZZm0dqOsJX94XVrL
zZSfoeteZd9cNfvmJmeKEZkOi1FehRspblibmWGkhZm3sil3pmIddKbCmjzWK2DXKyqNkq86iXTu
/4p98xGYe8Zw0Tb57PqrHX+Np0gzqjARtRfkyzQP2XZQsmttaWAD3D6suJU+fdRqQqDbBy8gLv3N
BJnVoJgURKzwiKeqxD8m9VlA03NUgJQkIFJVXAW8TKx/2tU6ajX/ABbbhIKGmxrtao/4zDB0bPhv
8AaleAk1xFPGH9u4ul8zZqOiKnWOS179O7lTs6CMlAwjKIjmf2GHXGYW0iGcV5p+/59LIULPl83Z
/HdLd8Wh+nlV3yUcBFMFibLwSMVKJUm1QesKDnTZB0YPLsD8CFSX60df4xpPoYxSi22c+66sc5Zi
RYSq8T3PbGeHC8MClejl2j9d4NmetVPc8yrYkaiF7KCokgMkDXAge8+aZJ9rO4pFj7A4ABAaqfKs
leqrwzFmrWnvqKJKrr6iCWZL3Eurrds3Jx3ZxfZGsKqWkhItTmdUrdheOgM9aGsSyF3/nA5prNMG
lKKMGCn1/qPWKYR9tk12YXt93xZC99+xPd3LmFTdnuvMPBCKgOt3P3l98tcb66nHfj7g6ciXmG2c
ffRjzdWCfUTR1kEyQHzqz+RmDAwbFhmIK/ebI/ALSDP9GnE4T5HthT65Xi2cdUMPkwUcmDIy+wzJ
Qr2gCV2x5MRCge5LE+3LZRvWQjBcWhsXjg4OgNlQS4f/CTI7A4xgY9czpnp1F1E/bxeCjvn6PTqy
JxcUBDYh/c9e7LEwEM4gclm2s3WLp4qmvueaUMJ99Sl2WQ4CRfH/9nsRWjF4JUe+cXkIGV2Xjgoy
Qw3R5rjYlkFmty64xwXk5Z31Aj4wTVZfSZpbklVcrvabHIBaD+ZiapnXIG3YQAJ6jDaVR5NfcLc+
kL3c7olnQSo+JkQZ1hIXdXvd/aPs1CCjICT8ny9kRuLRr/AyLhDpaD4AlhoIO++T6yAuF082j7iK
7Pjj5j9GiXQkM5OOMYZIUZH9yboF8iUbUyPtHTfwM7qM1tLW+81JLU0mamfWwLh4s/S+mHsnb0vI
dptkQnLlpHR9CLhR8uXN/IihFNTyNJidDLs/DnopgzVTbkOvLr6bvyk8zM7hWYrgIgb7kwcvqAdB
b/WoYeK51ft5sCBECaRHQhubifosItCMcavgrPU3iVP7yNENQaJDlUUWV1Lc3+a6ZMYoyUK+9B41
IB4LMQgLn4l4dlAHrQVxu6fvrf6CRv+ml2c6OKuuLxGG0k9YEQzkOtU1SmRWG7/x+f4jQ+hjU6W+
efJIKqqzPxACeFgOqxuWJA3VA3mmTJIALH0WokjTB/BEpOR9qu9NXCPsP5Rw8JCbmoSDe2LBH7b6
PVYlVsZXVdgpglRudmUXSqCEZt1UGYmmlhuF64qFbJgyD7fk4fijxWwPIvY9ETJfcsFi9p1gXBn0
cUTCy8TcMmexXeCAqpGCVobjdHH/lNDMCOp8KsUdoQQ4obCuHCcaIejWzSv4115f8Dqi5At/NDtc
RN0zL+4R+vQ4/Y18m8hpWxVWsCQeCCF8XovGHupoICGf9+9Ac8eQ0SxfQ/pcgOOEzjd17iYU8ydf
VFTMzPCBRqcIJJ9r+HOSadocVktnTqrw2bqs1OM8VI7/dtGtcr9gy0yGVKbWKlRdaNCTa62nPhef
N9+kb4diYicBNkhLdX82OP2YkRCRRY/TNHlKJENQENCcImcoV9gdPqlUtAINKkcoubYzx1fGApZL
pEdVVFj1+9NcqLJ/DAPzp6pM72O9xcDaGAjGPvEPlOGz8/dCiDhvb1KdpBcfGPEKemNqLpMVxHBN
+itB2FC/X4kuLiYJhmMGDkKelJOKcN9E05BK86gDOXyezGdtd5loK3jDYEk2b7uAsvyA3u1LVJ2j
QM0M7dMvOwpmySlGGM+vrd42AVZUuMdXTSv0xil7fc8GUN6tU2+bKOe8jJxxvd0BwzYWU+TbiCzU
3NSsQFSgPMIjlmEPWbmK596xP3Ifv7lpVZpWT+aeaPmjsUAddcsDHemqO1vpzDrnDWp9KUefGslV
vkFdEQwn1F0OQ1VELyTIJJ4kJKkk8ST83KT/kXDi4kb0DdnVKCjOhKxQaKfYBewcNdoX1miOZFM+
FC2bD1D4uHiq9LacM0QpFrjhRg25UjPA4U5pXhI8HSqmIZUpXUVjWndnjtoFekq3anjeG8rXnptr
K7512eiB7AJDkrTNavktUF2XFS4CbhoIBXpeBJQFQiXFnRIVXpPz2FJxMMAAN0r6j4yevi7cIbSU
voXMsYKH+6DRddY7DQn1ALMwOFTlbjrWl/UKjt/S+ccDWw4/e8Kx+ZGPizJJ4Gy53cVgsQ3Pryry
HGy+/4c/FwD01u+B96nSlf2kgUbWg5JrFA5wbyCI+cvRH3onasT3YV5MTG7VsO4T0ohX+gkpShQi
yyf3n1FHBJMrPNgJOr5s1DRD3fwW9uDJrdVtiZuuRYrxmTVfwBB7oLHlK1A5hapdUErrsH72osUu
WG3VJp1fiZX5ujKczTt1U+vHdk4LdxY8yfxDHwjuuzFvlyUgAs2deynJDHoHoCIwzWUNGMCMrzf6
ENREUEHKpF9QEFdOrHxwSQSuj2C88NtVm67/fi2oXsAIuQU43aEwOsYEj4uF9YFk1ZPoiYkvzCnx
upFrolZwzAGMd5mYboQ1kvxjyftFTK/5stnawAFomAPrd5R85yJokHv3GWiQK6kNDSIhtjX63mEx
BaXSKDHQ0IyJbk6ChxA4GKyVNU9ltuGhf6Geruo/iuGzMnnlEqi+K61w6vtQOMc0qPSPXkf65D1P
HlCEeYEkVUKHYuEK1J0MUp7AmvAiM2KbIBCAox0FaUMwQG+3xlbPeRnn7Zqg3ECiRPgD5gyXPwQz
QF7LklXok5Uz/6g1+D3FkJfkOEqdymGDd/xELIvdaMb3KuH/Cy2v6jy94BIZVk0SXubkyhQ4COwp
b83hg53GEkE3vVo5yNWh4JxuK9ZRCXu99O9IPyEpGv4LwAImjM+OGBi/Lf3w+u1mPn59G7IXWR/E
5mM6l1cYqKO6MHl8JBZwkrW31dfwqI4GLCjQNPYqeF4lvwCwQOB2iLHag+bkEhCKZFbZCh5q2req
lXuAcTDeSVyl0vp6UppZ2hqzAP5exfC/KfJnLkpWZ0DEYxTUkGVJRTb7AwPmdJdNGJ452jrFKfrK
+Hgzxsh8kkVEKMkNphMoViNuy9mlY8Ccbs1uS5YeFsnBNd+1JdBczzGz19cY8KDYU+Lb0ta6QFF/
UQpKKEBj4dCzMzHddTqTWHMQrdrD++dK0jpQqvl8sqiE46ZsaoCzI4ZUcBrkJnZEDLU6KRZ7i+VM
Xgs7fm23tWZlTZKWsnSzWJyPvQasqVg2YB6exo6YeXyIP1l5PisVvrCaM0nHg81/j8O9GstU0QEE
E6FVDXL6XWIKJu8CTjuyVsBwt/X9K+9guReWgH/JXg0lAxjKoisXKlUMb+Wa4UzggMqWdDliqItW
Xwk/19zw6VUTPDIHUKF8EdpUiXJuz/gX8XLSJYKIbqgqtN84LE7YTLAg+6/orLtIEhL6IYRchq4S
cNPOYdJ0CYJJjtt5y1dtyzQ4Hha5kPnHYDE4UnHqyTdcwmy+UknWHLgK+cIi2i1YmA/r3DMAaNFi
XKa5MATKN1E1nMgfF9lFMMdxe4x1VdXZePPHSgegZ4OhEGqbCTooRQUqr+tkXe9v8NqTdaHbZKr7
1i87yVKIJuns7TQ/jyUqyZAmKzDZXfKVstmTDd7l3qmLvkU1hYuxTzIWCp4LvaCwvFBVIKDXEqQ0
emVwumnNBIBSFlptLU1FlTCJjXGDXbrhfegMt0l8KkLR/EqQscSeh5Rmjyp7+ArD+Q9XoJjAr46B
qPzcO3ymvMwVUs4JnM/JMNBKzojHT2aevQSfGOPhdnV+vqAr+Fg45ttnGK85Vx4gybeGApgvcs3d
vDlqj+T74nWiUfjhXdbnbom+c4PWOqTwIcW2VzCu0gkB4ToWo0xNbWzod9PGfXyM7Wzd9K4X2hzK
9J2BAJ9qchpFBL4pvy/jvyOg9bw3oOFVrMGWoECfvOMch6Xcqo4SMohFReF/DlIHApZB1/qPj8BG
j6Xh4U2+6n69vHlJ6njFDGf9BiaKJtge1mES4eCXFivv26pE+XDVuPK4AVJt3d8UlOD2yBch9HnZ
7uZxhbUd5cWrBuP/tggNU99gPzX9YOCOEdeiGSdMtb5+D4FAYLvc4asd+GRw+70kvm4TyBkMedxB
/9sd1Ym12jgJdY7CBfCkqgunR9jp/gAsWGlsUWBErs70Mm1a317H5Xu7K99fs52AjAQRwgMT0t8w
/tqUwUdMYyeno+8rxtJBIhj4QXfmgDx3lKBzip/wU5UcEUcPynu5+Txy1D/f9LDF++m8YYTvWTrn
2V07GfSTpBLw9NHiWmEoMQoqUdiRf7VNrq1eTDqX1eYllTTxGYSxTQUnANYz7GAO9wOD2SC84Isy
y5NHNxnBqxPiy6CGGoZyS7WgttjY/iRJTvqflOZxgPaRj+CYG73Ztjr9i4kav/Uept5z7jJ0UKbd
oNpvGeZ569HOE3FimdAvgT88EoYvcddqXtYP45hWM/PAlhG+VNsDTzr0Rj36MpJ0CF61mpejWUJL
S6DGWGp0+Bpvg23BLqvYGod5wI+QlNfyU7c3aZ+UKZKIKDrknrZvelfO5zW4NEeom4sbow2Y25vN
faO7+W0pzdZraBSTZd+cb0H3gIGavaAtPB+OLhk1m37At/sTwQ9IzY/GFpEdQROv+mNhs3/Q4kK8
fyqT/fUh/ryeWi8EjTGLULjPe9iQZ1l2Kno7xA7z5V0W0+MbeNI+Ez4hNiTe+GO/KroPknMg4cEN
+bnqHZRhLFy9n6smvMsF9QEjpqBNixYjt3NyjuU1W/ROZ2muSlzWf3jEhaxzuCSdKhWs/w7R7txR
wqm7lCiGzxa1eLeo8i08CokpqpY5dQSPOgSSCYkD0V4MC25ml45i6D7q9YRRXAtcRPOnmv0oFGMa
IapM2ogR3UzWLerjrDZKwEYgWHLquE/2gw3kvYJxvG3y1JAAbOMwA4SEZ81nY2xuKSSOfFk5HkYx
KGF7CToYqxvWb1SezQkUpv/w1xdM8zcyXDFsibCXSzzEBGUl/4CAK0uPvbDxO033Y3DH1maELqZ2
Vt3izNbXivHoQXF77l13/X8eh5/RoZxjn8amB/Q3pFoqlXb9RJr/f4z9hxdX63ywEGeW+Ao0jSQ8
/HPWRTWAM3kLwerCJoLR2vp9vipIgQPhxMiuTqP2jYkqX0hgyCa7TRa7hfUZnboTKhtpgm81CJaB
DNhRqHG8P4Wf+1WOOZT/xxFNLzdCFx2+NW9EzH2MAV+97PlHDc9PxbiJnW2ZL1WWGX3YAktVKAFx
zJ7fHtVgjoxUSOICZJKjPI7p88XeWBtG6qkcLm1fPpVg2yVPCFYTa2MlGk/htUTwI0wuExwuWnv+
jULU6+DvIOaiSt13PSyL+hbgqaZnjhSquyWQr5AVvHzuTUCsgvx3hMMDKuahqYKrqsIvwPzeD6V8
wluhRawYB9W34CMfOB458uXR8H/++tlAWewsWFoY0qNgkh6cIHu76+di35QTTqSTA8gu9wplduQy
+3+a8mUNnVUMcvLUSa0aHVcQyhZ3N9z3I5iYqFft6MOxa1TtaGJKcPZQbne74sxUBxO2FhGUIEa4
Hnvb6BXzFRk9bEj8jucy62wzkbWajjEyHVPN9NvqZozjgKc8Ot+nPwATDklevJc/XxYK/ms4ZTMo
4jJ2zSo9vPEv3qFOyAAF9NgSyNmNs2ZY/kwjHv6zYRHldtm6ErNNd2t+sfkquU4iZYFBP4nHwbM6
Mu+pJTWyln9HN8aaBW93UY0AEBMuItmSfCqaUrmxkjnhK2X1JTWWrHeRaN4lyj/UB8rf/LSASYDq
iLrV4i+3DOAxAbOS0LjeLmXE2XWKGx5aYm6vsGFfeuHGt9f60bx3IVZ8+XB6u4dH9OFNqW9s5Eby
t0A9msWyA/jagMO2K4guLRuDUP9T4VcUWRKtumVyPCsS96QrcU23J/s8mefshh/DKJqX0MgckqO5
gg2rpA68ETuhvFhuVvq3RdMeFpIYh4q2/aD0B/jZfdcG5bI6cPikA7uoe9BR13GoAjRZoyrR3B4v
oS8fO/dh/gEd/oaVIySs75CJSyU9YgJGQM1TjL6xy94DwYp4uy7tXAM0kijdnhPDz+/7pT7IEcKK
l63U9yCSRaSbt5qisIn8cvgSXUjFL/eM0BUJigUtTNv1n5uWCs/fCT+smTN9WhPj+ioG54dpH5uS
3LoctIohkUPBmkyJNkg+NKibNGMm13hCCe3S/bSoZF875zXFV/rQT7y0j2ZXiyR1JYs2GbieIjKX
iB7mGWq2lIhgvD6/9NT4td9jfkwT+oJY1X0nCK7y7+d94dxBK1ngBDkPe54y/9KfP/lFNWe52IVA
2pfH8PYYRWHcCqFK6Uy1xVRhwyeyR3qcsYsNJYnokINjK0BsvdJjLdu0fX8xMbDtmYqKlxr+hyI4
RU18DLIqBbvPFjMx481XpouUrMH7HOYHUXOXPm7zCyewklQopYvIzdV/5qhT+JNfqxFCIX5mX7C+
Uoyxt6EHW9KrAB22n5gpOAPE4RK6C5zczyu9nZMRC5S9eGWr4znvAxtCe817Mm3wX68d7E8yHn5t
qR8KuwPOR2TAuDot+c5td5w2rloILxmeTYN9ckMQEF1/VrsxrFSs2uuAz4Mqp12CkeRqBYmQ78hu
2zoDyXrzWPKAQ8va3/DdWc41BCnchbbLMu7PpJb9rejIU3ZKw6L9yIOPJ/gFvg5uBlNfKtgeisPE
dNczNbSK7VbsMErfreh7udxHZqGU2FQdWZc3fhScE8dEpcJ6dSjF3Fe+tw8gVFgnNws62nOnvjas
J3BTNSHAXx4ko1ZMD4t5IS3Ry8y2g7TURjFyZkTUTSOPSwVP5Do1iImUglEy2+cOuwnSrfJVp3lv
sA1ex+gro46WcApYGSmAvt8qhyX2ZqIiHurbNtrYlBgqbUJ0AXzlwexg1wVkLn5AXJciyUTOdyEn
XgiKU9sRDe1aoJiMRaApO5E6tuGVWubR9AUhgU9bdZpfgx43TmHVD1pSPS8E6NUz5FtYz8d3S2Lu
vpzjM+SKrB/hfS766GWkS9YVyjU8pSa9wr4OZcLl923oyJnFQcHxAqWTgJSlcxxresYLVMMooSbr
e9zaBfOxgpWnht2Ch8OpoIEAqeVIQnI3F1M331bOVrqPNc96dhk+LRJkq6yBiJQzpNKt4C7hybgM
TaljFtyMJ8ThUW8CXw6b/Wg1vHpdgQvNrwJeCNCLa1HJhkWi5im9UPzUjKH9F8qLpFRw4Mt9psR5
pXYZR7DvMnwlKmKk7stGIagkmVZOhUumULQ22VtfwFcB1lwCIdxq0LTiOBLLdRWQZetb9x7Z3+S4
2jqp3KUesgdt8g97Rcxw07s7GCqkL00vmKZKwt2Px+bXKuxB0hPuBdLU5DFpL0KT52sD7l2Ygkzg
sSi21pWbTcWyb1I8sQJV2Fj/XEXl4YgUr4GRpLvXrxri3jJthF4rIc28Onba5pSVTlQTfFrq2mcv
xBSfHKzX98Ea2bHDITcubGVcrrbHPzy7y6qro+QVUeuft5cxLXrwYnWGk5vF+u0Por/jn9eZslAV
tkR1VcjsJvqF80bAKkxGHsNzlDNpssW1Gisd+X86A6rLQ24YnhER4AVSUwSCy5aCB8aAd7CTK0CW
dX+vnmidyIGyFsxc7J/wA2sdHLx5GH0HB03uSYaV0BdYq+Ggwopumqbq1UKEilMWpac6F1Lv1rdz
DgCO/oDrJhu4GLi+pbmYQAg9zvVsK3mx7+UtTdFn5SAYf+5IpNAnAuRCfTjPpznCHdZmeoS2W3Bs
+D7W6AO/rA/F7fgjQxWF2xzM7u/cvdCo/I71G/t5ZENScnOm9RQz8r36bixKfA6jxrZN9kemv47u
s4vZIcb9X1t5tH/WS443nYzkAwohb1UAcjcixGlnY+sRkki7GpL6DlP7p9onX3YElSiJzmc0PdNf
JRife3t3J9kQKiRvdM+CCKfqSJZNFaTMNn9Jcf/wj8WytQdF8FTio/UqNEr/1UA/KZO4U7D07M05
+juN0ZGB8C7ngVPLMqn8LgHEmYyZ2QKppXxA/8ZwVtNXj1q6tMhhCO9Y6bXpcncOXv5xJZsOsL2V
Aiqwo+DXCVdRTtId9jIeMambqVkjIKQbEToW2eMuFmg9+7O+iERSLG+Bz35CrYuoc4BccaUIYBgk
wHZL9TeqHkD49NNzyhENVC6muFx8r+1qIuXykDaEcd6OqO/58JbNXniYm3WhSpOUCWBsWprptpkt
evpArYz99L0Pt/WjSk1mtQnbUF43l4d9tJwSK5MI+F+JjqD8nOjsmQtWBxALleL6hDmAGnUaOSVg
8CC8k85w5jjy36mlWXWa/LbzKbEo+j62yRR//qmNqwrVZg1oyXkE6pCQJ2IZF14WSljQlkg8Mr3J
olcU5poPczZpyBxyoQpSv8mJi4UQcO/9B+MlJnxfwloPulCWsCGJ8K1X0E/PU0X1F4tAwEYRe1j7
rWJav7GGeUT5fq1eyYK90U/DnjA7H3AoVY62Z6ihUicnYg/n9IJc3FIPT6VpzZtt/VUrHiXoaEY6
zBgMHx3gv1a5+gP5mNvZXg93vPxOVz4/Q3v3lqhOD5zygL+ZJtUIuWqw4iMm8dWkRYo07ws9N+tv
Qlw+5+rHFNOAvHc4pypKEg8cdeRZ92UyUEWCD0rXS4uMZ6GK3FmiK2tUUp/mleZH6qiGGmIpDVZQ
hovkOPBBYpvO6dVevkyxuI5Gzx1BSiQnbsbGiTIcCmb6pwoNwusJ3Sn4DpZ1SNK4Gyyts9s54Kk5
gsqsVk6CNYjE0OXgWo0XkLGa+V2G3giu/IYvv7h7D7+MnOOXEl58w0fSbt/4Hqvrbv/KwTJ7Ijpr
UWcO4YmrGv0BExMvUh3jn66oK1QSzmBUbxnSn7Oke8PxdFw7xEZs2sjng3JsB7tN4BkPH5ivUIz9
m6riloxEcX4YtuHTubH8MqzpUJtRk6gOS0kprFbXK4xR0qAx+sto6w81UVyLPrE/D7r1SL3+XiPf
g7awcMWG/43y6Oq3L878b8Ly9SkbTSgN4dAWT7ESzZlK1ePrtVS3JtCLvG61WyyW31XUYE9Waynr
ngSMj08w/SsLM4LN3tMRNvzvgalM/3M6PIOKR35Zn0nRcLNhzOE/iql8pI24vBzT6TpxBPv6TaeC
66FTdIrF/IHgAWnXPhMNT/WP2QzEtFlhs2vv9BB4fMN/JrgEk5DqC3jE2/P3IzvGCF5bUeYV3J6Y
sDsRVCCPrHIGoF1rk50S+CflV9dv4onA2ab0n5i6ufS/IdGaeBSJLvNxEVJj0etGGO65irvkrBmu
PW0vULzcPJ09b7nqRjaNqL8f4RK6QIsjrB1EkbXNSLoMXIvV0d8ViHDa2uKvIPtZL22J40N6BD+s
RohU2lo1wcFbnj5niwZZF8+KrLIutA20hmdrwnPzeqirCQQkbMsBLJnjH2nNp8oFJkCdN1jXCgWG
oh+IYbhhRaMPAIaKbSTMAfFmJDiKcEKg41Hv4nAqX2r659eACib03TVhCPL1dSmKPpc+HLGx21GN
tKoNe+fry32q4tQEUQm9MpjEDluthlgplje9uiwQrqeNTJotg6x98eeA+SQ63oQUTProANr7sbx2
0TMDq2AIGabGIi0TsYwl4GLkbvnSfpy/s82ptHGxFFgrdcCvarNeUSNJ6otN+7UfiR4HQatIfyZI
yVTh0TLv3NorCdd+sOouuxMkWntMPJUQE/8y1r5Yu3I01qBsX5/ifKGM2GNAwbLPUKwOjRidd+hT
tKq8Sc/q8jPhsXzburYJBoLRpXDV0JZEovoF2dTncfRmdAx+FmS1gWC/op1+/JhiPThoWBx602GI
8t852cHdxIkP7mIYQ34RtmMC8IHw2NW38pMVQtutw0+8K3KabNnbxxGqJFqLrCWjMQ9OxJLiCU39
0NEEiY8Jm5UBlEtpGxh+2dvnZXxQRyD3IwmtQoPsOc925sXbnfl/AdEpbHNP5XQnXCv507XnN72y
1kAfXD3HhI+iUQRKdnmcVBYCK8GL5S+iysADWDk3VpQ3D/Q/H9bY3vXwTt83Lw/t5qTKhKrqNL2w
/lFW7Qgi5MIRuNeNOntdA1D80q1L0GdDiG5yHoZ2aUonjdaA/Jj0c0s3HdIcT2YcwgqUAlBAcm1L
xMXP95/Tf4OT5wMsJ9rxTDgwFzfMpjJzRXBzb8dQGygnHhV9Zjwz7KTtFLx+j1F03BZDHU7Wja4M
mNkOtynCf3p7owlbBZjQfmUCp/SAdEAU46hC8lvFklB/bqTcCE0TR1vVGtLGIuG4bRTOjexCdcom
59Wh9saek+wNprps81gLK7L5l+jTpaPWTPSgzM4Y5MWZ9HNc1IGvY5qPY3hGeZyHohtFqRAsDCl9
Znf3CqCvwK/GzgaDbvw+CIDztE55l0QLbXYdrnaNFIjVab/jsFPwMTqlBRvnGeBmZ6aSIYIemoQ4
ltvOcD1tMc+GUTz+0pHhsxSBmqYw/K0zkKkzpEy2iTSTOq5udzYNu/dZAgiMiFPmDVwdfklfYDzW
DNzYlLM+k4kRIM2C+3wbce7UA1D5GTwD/t5yx7yvcyWNdfe3AEFMbUd6hcElhJOctN+lKYLZcKen
j2PIhLVzdIz345FES4IFo9NW9UL8DOGocJDBRPMwgI3shiMAXFukjDjIESCHJtE565A+tNP2NFHJ
IGvs/4FwLJ+/PM1RkvOT/VypKZ7CkoebGkc3k5a/Q7Ld5sPMN2ZpJZQNo5YvmprxmU9RaDaxSpRE
UHbdlwo2AVHA1J1Fb2elZjHcScdw0DTz5t1bgrqNOGHYiESXkSjHFKkHeQDvlJQ9AUtIVSqg2hMq
aJ/Dpa4+s+kb1JrO+qbrmSugtLMFTvADFAjNl4miJS4wVdf3vY6C3PBZGFABx8/Aj8G80TgDA/C+
PBmhlwrMICSJXgVX48okWpamioqlqOcrc+PgWkxedw6wm4Cy7/7639R9X2+4s+hvXq8pt7CKL62e
un3CXcLsybgBlEqJsMtd3SRVM2ejENGjRYMT35Q4XfX0MavT4y3N4yiIelau9VT5UOK6LwCUtiXs
hsbw7Bs/PkBSf9rah3UrLMCRt7pWF3Fuva8uyzJ36yoovYvA/C25P+20YjMbQ8YfGaLH9Jct5ERx
9uqzDKXrBH4ya1NXaMn8NF38ZwOKkHBlbMasa/2hBPRwjYnrxHpHuigYvPD5ZreIq26Y+uB/3s1o
jXXOouivfY2si43T1m1umMT0hmSUfKWJE86MrKOaCYn2+F6sTadoH4niWqczex6fUSKxhoGRxOpQ
7VDZNhbBqkZcEokSxvGhBBbKWPM7cC6xcFL/BXOJfTnuSQccWoW62ygMnziSi8QpgB0wUWJGC4ih
gHJhLxE2eLKAQjiSXu339D9fy2ZcODishvICgMNR7wSAJPHNsMoI2nab9lHjthH0o3BYyylbi3Uj
wzkSDTFT9cmoC7s2SIgZ4nd8/FkIOI9xt67wwWzvIRQ0x5PY9m4y47U/QNamIANPvv4TLv+mhbRO
KCE0klFWr9a+3iIG0e0cmloc+Sv2t2ZOhQzGTIqqQBK6GN9RdFvFuHc7OjadepjIgDwPTJK9HhNB
7oV91gbI67tY4fRgiZfrlFLMTtNxa7eRLq2oB8w7DoblZg0NFj9bFVqQscHd2hgQmNhUkmuj0H32
dYq5gwCzBJHPaLfIObiMvPwr/Yp9fW96zlwtdSnsEAtilkNNbtAK5+6UJC6oGmm/xSX9t8zXotbf
zbqTAmkw4TiCTQRW1K/wIjv0aTp2ken9B8O62rwupli+1JKlv45OQMdkEY9qUDgI+zzUHDKT0gk8
j2SLJCmM/aHamPI+EapD0EP7NWI+1jbX/IvBi+M8QwNJc6kInMVgcEJVd8X65IqhWNWnoHf7WheP
pZeDBSOvyH3qg8cwkkZymo9JcerA59PQl/RzenC53x+pehF3JHnxAffdkVlKk75U+hijH4JdpfM8
e0nJCaQPw0u8td8yjHsMLPKY9vELUF1uSi0ude6GuUW9o+k4xGSFhtWUTH4CNeLgKhVor4B9OSYF
zMxDU6cACw+iysfaV9HmbfhwDAgE1DXgXNhBaQQwxZKIFC4djHM19lLq87jzg7cFHtRNJMtEOrB2
Rg5MkA1X7Fv1xAV+mWsnnVUJgV0MxjWfN77OOYSD1/Jr+4PnpEKWx3XdJk3A8Ra+Ro03uLYGSsw3
WZw4pTmsIpHF6k4wc18U5sMvMZWeW3dhUMymz4j56Ht/pQSLQFunkYoD4Q1WjsEvJEml/sk2XKdc
MXB/FMPLsqg4TN1zwZllznAeTBOlbNIo5Ba+/+3pKRc2iQzPyzu6gJRiXrTTCy/wm9uoCWvQU5L5
guie+6v+zvvoMypMYLEdPqAZAbuN3usAzyTPucpxWS+SOvTq4/uSXuWi3xeZGJpKNZXycKhmfb+I
rcTMMUZk6OvPkJ7m6F4/9cxPjhjMJLnnXjNbpFnKk3WetzTN2GHdlcyjKfwchpxVmzlqu9ZMffgN
TAHANaACgHpjYnC9pKdsZ/KKW0Huu4ISPmiTEQKbpXOi9ynP1cbdbPkff6WHlDgsv89oQE+RXXLP
N1daKcjIse/N4MHw6GbYgC4AiJm0jwX3+Scq9VIOC+5FZk1js6AfiMdg7dhOkEE9YEm3FS5qJmdB
G6E00gjak/yCxm0QfpOlH8GFZAyHPkrm12W9Ps35Enov358NEV7a/VYUhJj51bAHGqbAyoIdeSSB
6l3RQZvRR/WvP7RKwd99idSeCUdI1fCvaHZOcebbtPmuXEU9jbezNuAS69saKA4A49Zfl9h429SE
wK5oZ+WPm2+W/9oryRFpZGsb0jcc5kwcsqw8N64ObfLFT0DjNWgJnI8uuTVzChtBXMy10hPVZakZ
Rkb8URjcHAHHZF4023vd0Rtka2SAY3HS8TR+WafSdKck6tb6brAdd+BN3BW38KvYK2MIYP+SUqux
AhxpW3ToodlilF/IvML2RDHJcPgqYiDUf6ElMHchTaIRdqgOY18bhz2Jz5B/Ev49VP1cWZHZ85QV
n8wuYgTBM7xNtrJoCqVwk3tnHMHSWCDfqFE+PHu9R7blc5Qolr0Tvw+0+3P95px7TA9Ghxfs2X8x
DNNoc5DCoeSrMym65+4pzISLWvvzmgCgBoK+OKW5obZFn/pZdSel7QO+ksV89j51N2FLE9osgZKa
+gqWQahyGE9O8LuPKWkVJ2nHqRDb0YdfL+aR8pprjBt72n2Q53cZuLcZ7ZbgvQeQ1SpJ96aWw3wt
nTryNqclPyypeXEBmi/nbUwOMB1nWuODoaiqzHqmvzQ86gEyBVr3D7iclQ6ttg5eRMeNS/rcZMFk
UDPc0Iql9vaPfgYkDlNpuGRuobhzx/PVlvqKtiXthQe6z92NssPr918Vg0Qa8lh6S1emvEIOGGAU
MoOAl7rmiAfXhFvBtUZkMWspaOp8iFghJ26y5tVHC96TPS9SKXTyUk1NV+xbdQulS6o556Sh7STv
Jg2a35No4npXJPRDyn4ZQfmIcQ8/iMdmPTDLXEOi6SHvdGRvvwqKoOuJvxev7cDw9pUj1NwE68uw
UfEXaAEKBSNwiVbHiYnvT/tLZzB5en+/ntvFCJO2Z1XqRXB00xwL3h7ASb2yoWzcwmUEyn9h+DCG
HyytzTKrzOd1H/3S0gh4fnWWUmrerALxjCxzAnvF0v8wdvJf9dcYWXd0MNEUUxYSBv8IHu3HwCNg
Gzhqis9mFJcvot3XPosoucsaArVLOy0A4inuKqY1zyzi8y9gIjT5ijCjii4E3MG+z48e7mjxzYHC
LPwJqY2Vx8VPncRdm2PmbK5D3/vgPpuTWuiaEuZaqWtnKgDzFX/t1PgfTK4lKw0tIN18zBEbU56s
nk7hRjC7u1R/wsDFtfJaueUT5OjJ0SkU4LPmvEi+TM+5YvC3tbjSTMHzoMHiaIbt4trGilyBW26a
SoLIjVTC6NAZnnp4RTblHaSCdy/muIgyjYpcOcOAK9GqqyZiTYbWMQo51EVRNbgDcupNP5nO3KEY
Y7sXfqREPfS2mu0pDvtM1PlLI8Jc3gY7+8CaguA+L8xle3yQ6CV6/mh2UTWdH9IwedXM0jYlcTtj
johEBuipSRAkUq78YJxRQpYjL5S3JjJ40JlpPcbOFfeHlG3aq2XtB3BIojD9W2SpZd6NiTmhst1R
mtJpX/O3DoKIT25wuj2kpIOJmfDXBSTP0qFZSda/qyiMsWLyZcp6n+eNFUDjBuD9cYPj/snO7ysb
gRUFvEHtDHf8veySJuuA3aaECBIjxqc+zuNMSCnzsxz4PF21iewlvPDJh8hxirXgvXCtdb+TLDn6
xjpSaqnPHvcerU5EKH7BakwLN4pBQ4NvS1XiUyo2DeqD7epWeFNhkixyuPWiRjLl4zFlbL07y5cL
lbSK40GAz8osF6YYD+wTLWbwkCqylaNVjsw3p05KmykCK15BzRAFIbsT9SnPmtG3tfC45NLjhvBB
yB9W67Ei4Blx73tUr6l0fbDgAITnHvA6Sxu3qJR/QHyD5SixIZCYmPnzOcu9fEQ8SclvifRK4/UF
9njtflwV8w0o8RJWwB7tAQ055uAjmrNsbGPi4++mp5/SJPF+gWLkg5Qq8yxLTHSZGLQdwLMESDGG
6CeIzArJkM7oY44u4yJtG04Ubu0+DO3zrM6/8aJFGSr5uyGB8CGyyioMPBwVJcACwN+E/LWvIurC
UTqoprIJ/zjWMNeQsf6K87lVcZaibSiU4qyiwG03rHOrtr0s7tgG40woRCpOsrhzQ8uLE7jJ6be9
cb2ADOLYhULNxyyealTptFi8WtN4oJiiCSMIQYdnzXC9NNrCDuEY/jBqx95Cg9pOvaKaVgKD6vyQ
6LcK+5i6JR0udd733H4SoV6Bckj7CjvhSf+4mAWsgGm0uMpZweAVwD36UJupS4caWSUmEm8zr4W7
wn9cA+1LKMrLTT4IijwtC16BxbNCJb4l0akaZrou7hbqLJ+E+4xbMN3epXoFdvF84TrduniIvgUw
/NM9sQ7bfJIEmAdERYqQvGMgY/FK+Bgc+wIYJepUozgXbIKSaqc0+tkCs0lbk8IO+bfKSMpLhlOI
vFm4gsoQhavmsAeKUC7izYJ8fefoJy3zq2IfhDUAFrH7QbY+ui6wcRoLdpyUgFPublBUGiQCLLfc
ectG09wceJ3hrlBAvz6V8XzX2wvYxgXo9mcCUQLDguoQjG83AfoeLmtJ1RD0jeXm2JRLG4v0LnrF
sEFBXMrAjSL0SSMBZRrRzvQaSsvpgLbam/XNV+11izwogxK40J7C6p07yx+S5GQ7pSf0PRVluOlZ
Ss2rV0O9vaMWTxv1GoiOL0KazSp3BV9s2yimBJh1+7hze2C638FtV+o43m1GPL1r1UvyljtRyhp+
NyH+exXYqzi0VH1LsTWbENzRJY9h9HSFopDw48MX3WzeLlcJjYa8vwTQBLShepnI4w4KtScOrTYO
S+dboHnaYO+gS9YwSrXLHu65fM/ZTfynUG0vE3JWvQuDg8zSkBWi8Y6OfTKANkPPXRDE1kJzKHTi
xjr/VlPYiTzDOsYVpLEONoQogby5FiR8xTe3q3V1LW7l1uGkMbWdTnaH3TUzZtea5EhSJQQBFKm7
4iusG2QRxedthS3nnRAHa2qZ3FApwftAqB1M9/5EmED7vrR7dv4ZHzD5FdelwtJ68+DCLnI1rUN9
Li1px1bVDIYssyTO7NLwa9ZGhBOyZTZO6xndC1XlBN0Bc7jF/bFCIox89JU/gSp6P/oxtZ89i56w
lDF5Bs39MkeJLwzMhbfLAGaj9ko7gY5ggjYRMh1APM9AhP0zVq3d2/ALFLUL4t/TK+qg3DHL5qDM
t08suo/5QUIx0eSKxWHL6PO6rIkYGX0fN0eY9asAALSFzCv7LQmDrBVisSsTL6nMKLYhf4Mdoz5y
UPq1xLpoO2WXZTZJijinSt9yoejRmK6JIz/ki6Z/H+XVofz5+AVCMMWHz517w+UlAdHQrA50gYbm
4JVvjbPYSzL8GnFCFnhxgrWb+mLGZv8qOaRW/lOJvpaJi4T2ECTyE/f8i8QrddBK1nr77gi0yb7Z
NBo8+VcS8xjkQEyYs9tYwM9KxOSZkg9TVCyrtBsx6wHmxyMf7m44R5K2cJmCIZ18vN1rL+ucQJUP
DMQWnuZRCEA2ChsBCp6oz1iENJlM+3hFnJPwMbHRfnTA3FC0LHJWuCgtxHuQzLQOdH8sGrtd11y8
iDEJ1/DVh72dz7CODZMgJRRyiWys/Fl8TQYe5Ws21riFnQb050EUvJn5sS9xc/clwX84JGLDdf9n
70n+7LytZq1czcOVmUdY9iFJkGbJvx7BoibJx1q1Byb+whKXTvIfkK1L/Rc68D9GRX+CQHUSYJnf
IVnPy2kJN/x2V6mCDzSxKgTRhvuTx6TbzU4v6DvDn2mVtoZbmR5NUnEugSFo9tXKMVAVGPmSnWtP
sKK6xCulmZELrD+xeVJHbTm2fdsnRNd54psmzvEZbZ0bzeDrmYj7LprhtLEK04RYfrS11IoW2Dk5
awktpYoHMh9KUSsVxaazXjaOCDcGkKpVuUbzXwKkFR8UOgxWT7pkaP4bg0VN7j9nzXLmQo96deNU
u3iXI3W5q3+5o06VxgH453dZ6XtNi5lxJZL7W+I0QDhkqHEuUz7+3NtJIQrhGLZAB3ARQ7foGuMp
HYuzfpbZm6cNuXOEbmJZtGKbNzllr+CWR+Lwat+h4zdRF9VwkvahlOZCSIbH3X7o/pBpq5t0Bvgf
a1bjAsTQWmRBInthtkg0WbGWUsj6dNPL1GKABFjVnJhvrulgGzR+GqJN9cf8F2/sml+wd6jT4+3W
PbJZ/DSh2rOyvviA8Iwtg6Ti8vI8q7pHwJiZFOdTuZ7crJzldZyeZ+sPBTFxhbF3F8bFCkemYi4n
dbucIoBWSdYsyQ2iJMx16/fJ8X5eWaOTQNhjBoNMvB19Zxk8pphCuIcf9gvncGtIV/zvZOzdCdZ2
w43o+v4HMqZU7UH6Q+PfksffhIw+yPw2MitlzB3QhO2FLPKF15Eh3EmrlwZMqpV2bi21N+fpwxHH
SCQrMm7Bd5WP556pL9u/iVa0de+RI4E6bziuTMdQ1C/WpFub7QlLAGJ3eH71lIl1O1/QqjlwnnE/
KX/GpeQb6YCm48EATAPajBUGlx264YOvWTvqWGNdaBSOXYWM2GndrdYnZ4pfzToVXt3m2XuQuf62
GkJQ+D1CVr1Bx3OKDd1/zxQhAd0KLvDb7kdovlpPsUpf1FGdQG8ML5eTc7/VmbNdh80KQHA7yUOU
iAS8xj8LxHDk1YUT0J7zu6S6YSj29yCWK4mNCxm37mp7f+z808AlBeIioqis3p1kOz2SIqA5LFlb
S2cDmOyGkdwxgXAYbwZGbSDuGBLSbLLxtllubyTyOwvOzc9IDX/v/Mrg3IbxBDvnqF2PqDbmFWIj
EZ7KEp6Qj7yKOLLkWPfw1hCBUuzwOzalvymy2FUPqp8nwxcYfiEIhaSnbtD7jDUGH2bqthB4MGnz
xj3o1MUJnxmNa72ktXoo2c7SpHJKxo+SID4OFVl4D2FIIUb/yOES+9AwFQSc0SDdUva/hhNH1z3m
5Fx6Y8HKLEecoMv1P1uZ/S3gCwp/YcU7GOD30qbp4l+COaRs1M6DlVHKNHKPL6Rc9KEHT/FfZKsC
McQRD69IVf4BszEjz3PqhmyrzN/lLq4ROUg5rKslgXrifiJliMXvYxOKf/OxsDulVWchXt5vieUg
Gw5cZdf74WuCsh8AJOFXvVMPVAZApN844CML05HWy+fpYUtiQzxDYR0sLbWuhFuJOg6R8TTLAnpB
1c6VSjUQv5CuYrvkxF55P/LK0VTlI1u+bxV+i/r61MH9Iv2bcklG+lf4ycnelCOCpSouTdHKsXbL
s7UX4PD1I+5pD2kgsEmZTd7E0Zsup6I61AOe3YIFqUvjXShzS+pEuNke0chTTZuJAqWA+J9o7o6+
apqj9fmIBtjRfkNeWuuTFawHEqiQZndpx5FIrIPXnruxqSNghp8qtm8FzvJOB4Uz8F3TDIsdaii+
NR2Fq2xDXYzXlt66OSY1VJb+5p6sAISnswsDvRKJtv3Sx1PFyUhrj9K2JCaC1CszD0vloINGj+55
HlGqab6+OtjvdnUVLZhFt4xDDC0oyGEYSdF86LiljeNxspRv3/8nBHJooU1MODIBVXAnqzhalWH/
oDKtMRntF/yv+MuwMhk5aHYkg5ML1nnkPLN+0VbZgNpqjs9XPFjbEIbBl+oreDVnh1n5PV2w4TKa
7DFxyZjR3+o8jRxnIgju/YLpJ+Q1vw8w9EHAtjPoFcvATWh1pqiAwxY+uiEm0Q9dkxqTWL/xOHMB
AltzyLLMPtGEp/dFlrz8eSqxHWxls2KekIURcxpT96aekSN2y28jB1hFmB+wIyd2SWifmJbDICRL
R6oGyvnr5v7hCwovrEYJD51swRajLOI59jHJSIGuFqEIA39Ow4uCQr+NsEs/TdllPn/imZRqCnfL
4awRajLWkPK/NT8A8lmkF7n3m8c+2Rv6Hgqc2rmEBVdEDDDUNv/vkqZFqVb1WSCmOaN/semCwawu
qzVaLXJe+PDLlbzRej77i5IjwS4q8rnfZu916eAt4VoNuMd3uUniOxGM+itfXdw1tt7Nkm2kBYrW
k0pFRIrWOy2xXpoJOmK9/uAQ/yYS6ZZPIAykov/YE+vt43ckDwLg5LQNXG9oC/pjh7ZR4SnzV3VH
kKzo2LidkUSTSIPCGPA1KRAB1GPEzs4jI9PWCbfucF1lkZi7JAGwEVDmPtWJLuHTKIWMFcvakj+K
elQndzo8lt6y3Eo02sMU5U6V6QxRVyUTuUwjW2wfxKPebL87cyKsNi+CBOKYrQqNe0qCNflfV9Ff
31UUwXlIBepOUO6+dpx7hCbd/RmSHm5Lbr1z8Z3bAylkAeEEmwrAQIbZ11zdIYTz6JydSu0PIvs+
nfc8Grb61dGqFt2FVbNv63vl0tUI9psoTr39LmFqzXBSvkXUrT1OM47QUQKr4yDmGqYV+XYRvigE
ioZ00YTIZpnhAQC6PvYeXvELv2eOP89CSgJEpK0wuc8unBKAvw6nidHfzPY8fRe6/zzntbYb3eTq
37BO5VmtXpPrHU6HiX7u4YA3tQ+FSeaRI7wDJJnnf9dQzRB1smqLKx16Ynr1o2V8hOKwbEB2HeMA
z13FSmSOAyxuwpPX8R40EvAVsTreHMThqeRBKMKg+3NrsijphAXUrg0uNWlCD/EoaGVCl8uXssb3
rPXuOYJVGzgOvZuO9tqZYecFN/PplbqnB6sM8CY9l0b0STXvsNjJW3vjlZ6y0P0U11F8jPERkNpX
wO5eLEiPVdhJYzwxd0DCabbv1R3dDOWN6Jp+nXhaAJapO2IssPUZx0okr4kSwnBE/eeZ6CkFJE+N
vfdrGq1yXTOfQU1xE4It1kR2cA45wnOWRUubVN6Ic2X/J83Eq5XJ6D8NUI6zAlT7t+lo1D6ocW9k
ZwHz3mzn4d2bPSGUCYRtSpTT6pg+N8qzRkQkeoLBj/+Ys1SZKAfA+kxTdUIChT+C+ayhRJ/B41dw
FEBWU5AudfrpSQJwNaYekDNvKx/bNUA5RubaEyyO12ARyiDPTO81xDUegShzwj88Eeay9a2fXM/R
7oCKIIct37GTdaoaRJH9hyDjTivKzIWIUQbcOZNiULP7iiI0eYT+m208YRqpeZLGIHKkXGblpBpD
Cee4BVfjMdGNiAtT2U46W6okxsHJK8owLdMQuw0WJttJQZ8KmhX01Ql6HZJETMUW0qSjGRe0xySm
y2xDdiU1i7AIwQXslFQb9GfBIE70zo6TUFgb5n5oN5Vh1BxofmOlexIVJvWSI5xclY8v7eAwVsIy
kKLTiCg6hh0CN0lLSvNj7YypAeQhXuWPh4TVob7/co8sDH7B8A7OUT3f8N/3bqAObBZF5LoTr9JV
hVm5GV+qHE/EkNrF3plRWiFEQfNxssOq6Cm4Qrief4jbdjxrK654/1wmt9CkDQA3LsSR8i6RkooQ
f8ITIYciZj683XZ/C6nn4YjYmYtI3QaTTkZeoGgTy4DXLLzZ8LEYtGHU3ghIhx/Toc9be2fmYxdY
NUy8+n9pk7xK3gUYRkC2KS6j6KPgf+J44ZkhLCgNseJBFcrk9nFd1bSwXbKIqxS8/xQqLS1fGZ1q
FslDgflDyJJA4lr1vqxFBsNskuH1wfHx5J10AHDt6dyEg2GdEmLexTq+OcOYpV6B8VE8MpdPRafz
GNMy8R2R4lkCWkf1Kgt+ylgDYNx1BO73uhux3iu0+jfLhQ+T0rkiydwrfx9EvEdxJn6dfz9YWcsM
OIqE6mSJjBo3duy/jjtUkT866jNgDcAZhUtyzMDNz/nJNHKXxeLZKBmVPbO7XwXzZgI4MP8c4Hfr
QLzn3rhinu3tp0NoKkGfTzIp20Gipw4zcZ6jW/DEe9bhBVvZSUm9NI5V9rjy0NFCgEjs8RcqbWuS
9oXqLstMY+4z8FKfPoG/jTaB8nAHLbMcUdxZvzYkoMbEVarQmXk5K9+U8SrzjBehi+bqcz34e+Cp
Xnqag7SLc0pYFJ9Md/yJdXE9uL6nAYAGapQ2grUuASfG6JCOgs6MdApcAnLOxa4CENa8pOn/TL/v
oS2Wu37pQ1lmpqgs2EHwNtt2r8qLbYnZ6sy3XkS5iMPX3oosOkRBRdlTpf8mUCC7NQIR3GAMmU3O
TfNb2qYjNXiIFQUBAXIcpTz/GyhT11nWu6c+b0E/cksuUQuMQKE8cax758wKY9BBIY8YFNYLUSts
tiMlXFAla0lLm3mxdXpdTFl8bnXxdntS8CJvtriYdDRtwmWhL+AhzrcN5lOt0LbUD+O1POYOTmxC
C7txNqJbm5zYIiwbm2s8X+PwZL2bVPJhZgoQvcb8BzPUG8PzF1/qw0QuN57zwokw0Zj4rHHad8RJ
8QCtHmdqljbfwQ+HMdV9eKtejmi+bce2uVMpNXpiYeu9BMxAAT4R9DaobEsv05rrPLGeAnwXvGGu
k2mCgMekL/vxiKYYiPHVHgWG2LP8PU0sSLK34LXdmj6OrU7c5ypR0cFgQxcq3shNOYQ3G4TYH2oh
ud23gZzbOORH2dKDXDhwhXLKv5tvlHAUa6wKI0SytdeflsM+X61stUB4VNSCPvj7So3l7kTilYlm
WtpVuJT088cIP6Yv64PGYnpu5I/KF8kRQcIEu9CSogcNczWVvZpw1cVHgsWEgspHQside73b+GmT
8/KSHZPxb2nJVcN4Ka3e2oK++Tv506OgD1GatOXTBNrfW6znuAZPH8nqxwoFwsLtGvQ3H93Bx+S5
LfgsP4IwoWUQ+NFaCvnsbgihKj4NUXBfSYGu25xksytHEid7bZ7BflxX70aZAkYOG3UC1rdpg/GP
QIuYTQeAPa53ANHvg4SKvaxiEzQgehocNu2PveCXJpbCPUlLQwmgCztczjSwzrpCaRyeBrao/FyE
eJ6PTZ4CljQXa8EBUqKZ9UcjFVvJrmFe5cBhe6dHXU2TIHC6TJu/jGizQta217IdUAfFmLB4FFSq
Kd/axs9A1CibuIjOUq3xZLjeKdy3p8qfxAOIowXeB6ZRBgWZpqEU3QCWxEMcrLXzTD8eNcosu03l
azILa0vHI7KZ7UheGRIiOwxk6ZBScOWoX0BRO24KaZ3GANp5ArQL7bea9zZGQbmBF4MHE8gGu+iF
I/EYH0pSSzu1O/xsWGub5HSp7nO5Y0WQo1P0AfXWyRZg114ezZT6oflEGwLF1EEVYxzQ2x5EheTR
XT2J6l+VGkNcV6APHlMqPF1p2/8f504nli7RoXJDj+LRK5N7e8Duvr1ssxJ30Z0g3/Vjwwd0Jst2
Ah0UityUeQscOcjW6tM36cumKUGV9sdKCo/C+hlFhPq//7niCcQL+y7A8+QRbBxmrBNgc6vWGnV5
J6JO9zSAHfYF7rTT+tSxdqNMHhMzVRKbe+QAJs27mXl0fPvkNSvHXN7d3h9HEVPWEN8vCJ5lVxpA
lMj97QrCeY5u2vRN1ssEoH2umqkc+Zri3hR49rwt+2KEh+xlbfX71E/N5k7sq5Xuc0kpSZ7+1SNN
wgvNNT/U2nu6ESXIhLG1Rfy/bZkGQPHH4E2/4WYo2L4sJ4gTSAlOClIMwRYwUDo90o5NxalDFdbS
JBK7pvUFd8yC33HA2Rem0wHNtKzNsjmwuyHA3UW+Ng3gGlJMeCL1W/TC7LU1wVIJfoG+eLrlKZ7x
o7frcOr9MmTNnTlMu3HVF2fSWtqhLYsq3NlNNA743NUYONllK+3BwHzl4dJMuP5iaGN66n4YhWzB
CRorRcAS870ZhtSSLTtWej5kaVbm0WWZ7z4pte9i+urQgpOSjkjmexbGO+PZu8hH9Mfdaw4PIGp/
CRie8rCF1O/dV+UsLZ0+cMjadNt9cC+7NV6KAeKclAoDr7iDGbeLkB0My2lIfEZaH6VYrP26fw8L
ns8wq98AYy2QNze8pX7wK3hB6NkJV7Jp38TJ6wzn1W/gKazXmihzX1rwb8KUs3/UgOteJY+Bn24p
9ZN/IGSETFKMuu86cdBi62VVEkWIYLcfkD6/32n9Gzcuu0Es66zo3BtKlI8EsmeMh/1cKbIMQLdx
Dm1tYpQQcGhb++HIuLBnTYvkKr/lLAUz3RXF8gC1bN9gRlJJ7/pygIWxff31d9dhP72CZS5lVbRH
4kaOGEEoz5ihYsNpCJgGc1m+ZWJMKvPmOgrdyTW64CsxbiGmX1qTu32AIpmr60WartBFX0PuUVnD
apLPRL8X9cWo1hNEtzzTOps/0OTHno3nlBRmGFS7zTrn14lsJekhyUm6TIZF4ZR5iXbUk94r7xYl
uVLrZWFTj4hF/KwNQqaxqTMd+thOaF638z+miq4HUvY9DxThgCuXQ/lTbgWWkEuiH7bkzbcSFqgl
xHUoPLyIrFRw8ADZEBp3fVDD8aouxfdBjm0eGhq2J5dc70ij+5Spc6zXgDweXEh0LiGtGb5ZL0bM
u258Z8RqkSiJy2OQeTUkm6ZfXmzyvc16RMW3Tw6dno2qN/lt1b18eeWQXLMu0ZjUvsUChFK4x4pz
8gftigbMk1Q2oUI4bSb5QqD3HK0Wd/gT7KnCEYBnz2ZGSEsAKnVRyf1Ie96+4EIlzlhffWAGjt/k
h7QvjndG3GePfO97ffkkjgDo5TKkzoV/bHDluGK+H2piJoNurZkitEeTVl48CtBWpo5nYZoeZp30
u/fFXvHgjUpkgmfQfMpcb6jVavY+Xn+5hWR8MW+spykD963T2wHQikW3tykUgixZpcWRMmmjDQWJ
epOoWIVLBZASbHJs/XSTOBGCJ6JQWAK/q8gn7HXkmvNywwgA0Mw52MYES2sn4E8gECWF/zYV22nx
qln0RCKhiniChG829HHbt0+xbVpnA14ehu667b1dNeJEtdQfE6feEzt7aRKY0wCGPIJ1ZyFTWmzM
hRbR9M3k0fq54WJx0sXhNqgm7Be77eVcZpvi7LCLw5QKBlnUR5jP/huKzTgZNLxjdHyzQn2P9ORK
6U4i2qvUYPrVmybPcZaQ534yARGhTX7Mn1R8BF8tBChqJzKQKitD18brvzWoCIspU/evFDdAOaHp
oZmRqvf/XLr+YFedLUDsfwAwiXymTQfUAJGfnG6ZPlnJuORvGfHxU2qeikJmr0boDJV4n0EXVJlf
QWOKgUvZiTRzq4dOrp9KpuTbZIugAQ0F2t+v0rMizX1piuFw/4f7rZEtQqx2LFy0CbTUOtrAR9yL
apsTzAuqwGoevUajycun1Mm8EOH8Q6S2lsSf8Lt7h04CQa2rs0//3Fp1vKkt0YMePVxeNDFOI9Uo
XKODcmkqzNsvYU21VgACb4W8MTQTZW23bFbMMhMSuWe8eYz1er682R1/pwXyvcigSIpSfmHdK+lN
AwxYHYkrg5oFhmovJlXmKnZVM7BLerXqzwBJmVNVGmSGF8/J15CUFIHfd8B/tf3AAa7DMf0RazxW
/7KQ8g5fkcfEVgdnS+KF/y0MyeCAWypuvmT7zWScdDxAuee5ch0Fbs73SzUC+tKH9kSjAhFBkifY
FNpITb5nH5q9m5kTwka5q4GAg7+K2TbKGNnPaJ9Tb1465ZR4VW8VAL8ca847lUfDPIAtzKZcPCyF
CcfkWgzq86Yy7WjQKBRbuCBeb/JYCQX+ao9XWo89DLU3FSu4/wh7Xcx8n/86Ju4o+HDbdw2lAvFf
D/gP0WeM7V5ppuWKZwv7Zben9qCKEyP/w/i4vbd+vYEkHNZwa3l53/7+om24YzmtJei11JiyXPf6
neTPlgEO34Oeft1rQBDHtU4ofhQ/MGIhVtjp7vsNgFCF0FL3gnqmfzrkeky96QYQfPi3b1/Nel+3
y7EZluIpqNqOdY/IZxWlBV+zF6aamxJ5e5AHC6H7OtEUQw3dPf3M2aZ5DNHMl9u8NkKu7X/aF7nd
AyGPzBA7qKL85D3XYwVKjXrY373NIJ2h811GzhwkaXz9KfQOMd0/SPQmXDn2ujXM8qi971hcKcXa
xR7ytgT+WPsIbX6uWK4T982GqQ4oMd6YjmsHIYQvKwhlm6O+MKdc/QMC1x10LaGacg0h7LJgYBnn
OC/y/aBDvvuVCfJc4cF9Y4DfcNYpKVwVhgD2t7ogqL2ez6cvysVywrZrCpEhE5ZkGJzrrLLZpl+O
VJ14+c1Zo/Y4yWAnWDbb7vA/Ogxlcm1HKCW7hjTWHwQsBVdA/8NQOH5PO2xo2myzzPzDw0Kna6hH
Ui16eCCX4mz7w59jHUmAlrcJo7Y8gXs6hThGuAX8hkGw2gBcT6QTIv4aTNPzKoeax/Vc5QD5sOFz
LAUGBqD7CewaZZpokPzMuBzXoifOCMG7VXQJ9hn1EUdhK469hgcrL5ebm9wDH530W38LVBHGu2ON
ptlEP9fQoiumDnEgggviWV1jcyiKKFpDPao4M5a5Izf6ykg1rN3haRpI0qkhGv+/SjqvPxAAb/7k
OyVeIw4gByZTIDmROwfoaJp5LAzwTlaJBgKRfplc6OGa2EvSSeaD4ZK3V+VdKFCTCvfSW4AdYl+m
PbGI3SzyAnm3/bMtexxSPQG7KM7FHnzndl62D0Dr+3HeWbpXZabXURORB0fn7QbYrbokjzltooyx
yuIoH8cAd9LNB84Q8TvgjyDWUGOTgz1GIlDwIMIiELmkqI6UKdoMBQ2kDRG0KmhAuO8LVwVWOT1d
d/vYHmvEREJphRQ1VMGe27rhG2kw83oof7GQB9Lb+NvZ9rS+6na9ZE/1mWFpFFZ2wPOETsGTy4V9
wz8qdulzozOF/J+pAS94F9aQrBs3y9Bs7LX07uo9wHOW+Jtlo0OmW5WJfn76j3HDYYV2fMTaLMC1
bczQRbyY5OGB5TkSlPpiTyIHhJihn1SgTVnRVBYB8pMkzNFq24xiVOupNkxxrip82/H6tVaE+FiP
zooOb8V/TKdva/aAXHzpc9pD/aoG7BFMVsw0M3Xyk0/mEEJWQbCPoqgZGxGa5XY8+BYNtc8bFIXt
06WTfQlD57sRSg+nfKw+jxI1jpbA0K1D34KzUJ7v856AmSymnIKsB6WOmitEAXYdw+rAtj184Tpw
H+UauSitSjV88eErcTK/Y7glvllgzIisYeA0QqJeGZmsBHCo3CE7bFJ18OHqZaGgWKleR0dz5sF2
gQJnHQN7Xy9GoB0IHyPJ4vVZhsF20TOluLICeJ3bv1ra/onJThkQuDkRQi2fgwXtbPJIMkYCg73y
KYSPQZLRtShT/GCxjWxtiumG1rym9SqslSAsyFiSv0Si91F+GWDXs5jtZ80K1pBaQtVtux5h2G8g
EmnAVmqcMyvmvKgoxGZwIzCX6aounnDwiNNN4B+bVGvHqSF3IhssMPfgms/z747GgvYkeo5gn42L
jOHeWBzX5lMKp3rNrFKXG3ZgVZXjiokmlkYjP8UMSUNtKVU1Lhz1VuRLZ0+zACz1n2EdgJWXQXoZ
JNsONP+ASqGPyJWpUsSE8N42Nozf2cn7yHpDOo8d7Xchh1ebZdu43bmtavgVT3lfPYvTjhOYR7vu
Jka5P5HI19boTvGDQNuM3iJmcK1OClG4Z33/+V2wZT0lC+pRdWqoZz/IQ+LxlNyRqxamg6nRzsyy
5A4pyEty90A/5aobkrBAe+0w/nxpg1VWDjBtwml76NrqVYhxY+BLqBcqWi+yCeSDEmUxkn89xEuu
YulCIWSRtR8VWfdJsWFPG+gq4g3GQ1eyxFwVGioOIVt++HvF+VTJk25fr7ZBJLAqnFl7XyT5q8/9
1dBKaqhdbY7+q0FUcrxYpqqqu/zzWq/CLcmLgWCEIyWNgEsAJkBxVzL884qQ2WHMaktVKbTPxjRR
aRWfyVJE7VjsQN6W+qHoLwKBvY/XktYZLPMDQ54YkB+hvQEsNwIilzX6g8j9PYO6p3Co8usWMP3U
Z62hQIcBYPYMkMN/nmiARBdVia2niQZBqmZw0RZarek5UNxDm0UHAx7Q6hNRfIoYjlOorFE6rW0p
Q2dGGO9OfunmBeio8zTgKVKIijobDqRQ88pvZgMHI3oMingjwVZhWnO/vQHuuNXlt3INz+yzt5me
CGY5Q5l3S6egSmz64zvehxdt6Q+PNQgzyoitlEIleM5tfvZ5W1ign1IuQgc73o2X1K9TQprMJ3ju
MS6U/oAWm3GT9Pfgh3Thlh4Mm3LHjEsgdbn+UbSSRUgT5qt0d4Zej1TaUf5VKepSLmspa6SEGVwi
omoKOEofDmAaKREJwn4U2/ObG93Mq6/ZvPE24d3EpOQZK/LLsvinrb8VqruQL/wHCdse8Me4aFz1
xUcUZZPgnVMZtRqkzgWs+omAmG6QJGYhFu+wAgLcHIm2WjS+BHx76FD7PFuRwFAr9BjBRNLrvGpV
ah07r8LnNhck894ff424gCT+3PpHOb2bwQwOMJHY7ApUqZXyYMv+dXTn0hq5A62h+gPH5vTfooeo
9EzNf+lbTks1W5WXV9ffBFNykJE1twzBAQaIs4MwngJzp/t/GdAxDKs1+tLa9WaH/toMq1YdqsxB
tHCnGpJoXD1YDPaXFESKAnIMpawA78+KDJcKUUFEc1+N3haqhu3VvWxThtP24bRDXD1vPfoPavsY
kYQHHXY8NFu8oQL+vcy6e8CGHrnZkdPuEP+dOdGwKpoNKFhJ6PQq0hSzhYnEa7jQfrpyYXnrDYQ+
hAzeVSgqjlAmOECiY8oFXdE0gGN62wP1/DK+8GBlBWSfwQGXV5Ta0NNtjfmaL2XC40sKx5BB4c1U
6mvCxo8ZhGbbEUcfT+Q8dU7uQktn/A7RRG08RjcFyOHVcdNtzxO1Y6vIWcLZUDkd192qE76fMcYP
Mg9SpDcLVMbJS4S3iMXhZ8UsP4FR18h1e0RPp8B2DayojZhHUHekz/Z4YsyMdRSHfqXAFXcLKxu+
6srYajP6wxfN76e7SL0bNngWJlHjZGjrtgBTJy23VcgvBwpHJV0DRht6kKOobnUegp/1ksf915vC
GXAbGVfG8SSrWCKYYVKeSpAoidPJ0n2za5OvQ7qYwVClHNEl4U2k8NupKbboxan/o91aJ+FGsWbr
YNkOBYe66m0D99QaeAJzxL7zy2hXBejESxyXCVy5CpmYoBmCvkrC56j+rZwkjQyNLnqKqMkyw0IL
J2zQKlKAS4WgUHtRx0Kkd+F/JQIQW5UTlmx0N+klCGB3GwLYeXaDzotFFepHf0c/HVh/0ypPqj3Q
mevDO7wiGVCws4B9h9QBZihUn+jmRu0p8dN+nBCMSa+UytkNBZ1WI/mFq6H6Du1O8LmuiaUUjbf+
PEAodGHiYP5PvJtA/JNoCIm1UrunRjztwvSM5vDpPSrv3mX/e8QYDMpPGW++eetWosLJam8GqpQ6
65DIwE8R2PbCepUiaKKcli+CKo51JQwa2+3MwA9aH4KTj8UDp13AhBXSpPc8MKNIgLVv5YPmyOvg
iLR7K90Dkk3EQhH4H225rLOoTggpF3WbLrPlOsIjyHn1xvw/E+VepDecXAzOxQtFk33sIYMq94DG
t584xs3X4AOecZNmeYxApn80h9eFqCc0xoQ/ukerkkIIQ1DR4BXmMmmVr6uKEfwlfBVkYfWSq4Sb
SuM7IrdpnFVKGGewRO4PJPViPTsU1hnlqpWubCSFehaemYQ63ByhfDcqWMShBlgOj4rzalAVbikW
cu/kmeydj/8ZpdTfqRcOmR/sX2Z99JjJm/npenXVGTu98W2v6uT/0PihqHTWTgq9YVwHKZs9rmrN
DAs+//Yl070u+XCYPJmkhThJ6IR3r4dJWG38zIGjcSm3a/ybm4Vt3e0dTekDaQJA4b4/3h72bC2b
6yJFVQr3Bmj3FvaZr/FON5IFGjECsEcptXKuPlbXh1aSEcJITQYPBFBaTKIBhY4nrht6WITYsw5U
QBTg/nUxPj0Rrm5Omx0LyEvZqIKEIQxB3NiHiFed9N/UoSEa1EipNVJki7tXknUrK3cUXDqgPG95
qSand/DIAfkQlzValnNT2G+G7jSiKYVbpnsVc+hZzo8yw+tT1aVpbJAq8ejfDpWoF0OpeFvIoY6E
z+0Xkoc64U87Od5jh5k1lAy+63vC14PB7e+q8Z9WfXPXZaPWUJnhDdUXpoYrEWxwwEStXQ6xe+Xk
4WZNBs7jh58y/tlKmA64CbKPiqQBYMrLuPeJqEWcsKrsGepfyD6lywwcceBc+zXfmOyVIw6qoxSC
2WcPlaV6BT8LH95cxUHpfQ9WCp+2E2OPX8/NZ5dOwvu1+Dd92+1GSrQcqXcpncfxncoE3QJRkK7t
8envsC2fpfJtbDVQEU9AMX/BtzxLLuO9kbS960R0YlKd7G48CP/CmxelmmkDqFG89GzJQlmOJz8J
L6z8CDFXbqBblIqLx7M1wRRH9GGUTvWhnj4JLieXMI0Gh9HETuMbIOA/cntOwRPVn1H7Kx5BWdVl
w814csfZJzt1J9ZyL/PRKfON/wDLyIGeuveSYdBB0wSxuUhN69YKT71IN5AEv6aBZtoqh+MV3pxd
l+3D1ReR6T3/bapdPajMfVHr3vPvh3oqef489LGOeElb/K5MwIXAQoNnisLuhLYetnRoS2EsYVEK
nOEyj1ML7/n9c8ZPQLCYXcDutF7mZS0CF+2RFA0KD7Eu8EIXLRc39z2CejLQW3qidzpqsCyWmVri
rY5gADalNdsQ8UZQsnPsCiyQ3rj4fNJAdC44vVhfSmwrKSw3OCLFTduO4oo6lb0HBFuktmcG+7j1
FopFbY32h0Gt0McKy28ysymhTd2I1jb+IDKT1/Gyqww/Idru5yZ2TqXGaayT8RApv/SWpg9UhQ5u
9+nutxH0x28FqUixmH9Ej+nJdxR/ZRbGKe1WqWMu7ld/a9+oeMJdacZk9A8Uv7Hl8kHO4lvhiAle
dWiiHrjcVsux8BklGU038gMi9DkDdxF9OozOztPe+VoLUNluMjOq3VOEvk3YbIOsELrYJ0olAr/W
NOVEhaAm7sD6E96SRGKFJYG+uD8XsDjkX6cUZPqaRVxe0DDAHgTszPFSv07Y0/XN41LE0AIcz6uy
JATjCmIHVKvvmoZzfJqVWCsVoINMvRVP41tFtlWcaBBh48yBIqGfcMHxO6fa09EwqeL9yYq7AsfY
rN23bC3XqtuhKM2PxXvdZqcQ6AmXrDJ3C5swLFppE+JyIx+fbBmagHXr0pw5ai7OMl8ML7ys6chx
OUk36YxFoSf3tYNgN9hFhdfJlxidECmggQPOvuaPJntqBlny5ewJuT7RsLaXiVhv4d2RPapWaCkt
vW4suINFPiWLJD6yi5BWr8thTtcGkJWHCEPGEt30jynl9HK0RIJ9+Baz9g0d78uqKlFJqGTe9oa5
/I1F8Vh//dEJqB0ZszXPMO2jlZTIYFulyNY0/eSHT//UuK9d/oWPHP6u2V65sEi4g/UnpUDWPVxA
bVzgNGYgLB28QW60bfelPGfwcailpcIg7Ag2cV+sHepuVKbzze9kekrwtPSXYZFgHfke3rxhYFT/
etXeTf9WEhxEesfUVI8/6ZWCiLERGk5s7QEsd6coWBZcsVU7zo+GTi6Am6SiuivplTDoFT2WWHxO
kz+l03KsJeDw8LZbwDWymTvjJ7T2xhFyiBa2yKzoeTB3Ce7rRl4RZpZPA6uigXbfSL79ZRhxBrRy
Xuv+izC2Sips3LTJpeSTxIihsNnBtOEJmS8YSBymA8IHRGZIkOrYNIXA8vrK6NrT9MeMjKs4a6ki
Yjwzo8PFNh1coPTBbTiFlYp2Q58Ow6jLFFB/HUiWbY3x0K4kIMoTK0EkaUeGhV3EDlD8PoyvwTPv
WZ54Hn9pZsVochh+TIfvSQx/liTnkIwdTJ6w5y+ldTObTIokrzFmsHoS+rfF8ZhtXgMpIV4WbQoB
kxcvvL8OY8g3AY2c8ZdmQqQnOhzy19kpR2RXgRup891ZcIGZbQn+R/GD+aWcyPevquY0Ng1eIazZ
5cBE5h18e8cjTWiAv8t/ZPCI7iggY49z7fd3orE7T1lYJw4gQsrWX/16wqid1DsA/A3Lg5HsbnBl
WGQjwNsF2TZcod2Cl93aaBhXXNjPUxX3corzsaC0zPe1UZhv26/2+32oUjU+xk7lfoXFSrFwMOik
bufzXe6Gcs5cO4ZBotRTSc+hMQoqY9LgwpQiV3XTveYgAvE5bbiRs6bvwKNurOG3YoAhqNJHTTxc
8R0x3PXL8UdQ8Nll4fspRxULbBVwpc+keCslwkHO1Cgs6JpCok56QDA1M4D/C0v8pN0HQl5NNxfg
5gaXIBkdTmWg0JKtwMk5GQfuLcaivYeUYZimqTC6iZnyuRu/8zz9dX6UduBlNz38PM9m9rVAw5vd
CZ1oRvIOsbEU2G503oWiBUVoP/bwRDDLp2N0sNNrbuoG7RfRk3vxD+ZWbPbC24oDZdl9mMX4YnCm
T23D9EOIHyzLg9q2qu46BeAe10I4nIhMbwwP/vWetwRdA7+CpECr6kld1dLg5yIEGstf0FJQxHf+
tNm21yWujRMkVCx4CmBEe/nP0CYPBK/KU1lPAYPZUI7/w8qC1f0xdm47sJBFj7AQCVo12VkPs1if
p2a8gvJw9b05iWUl4a45XhsqcbOBm/5dSWPA5HHP/poFM3dxiUG+qBVGbrje4lFExhZPIhjXlAuz
C6Ya5Eq2aj8kzL6HNdKDHwd1nKXbLoXfqSn1dGEVo2ana+2gBWbpO24l/66c63WGuJyga/vnqFpE
fmuMi25MesWVIAibM4fuoixVJ+Zk+eAuOJ3TgmOn8I/G6uT4KxeZjbY3xOtRvwMFMant8Ro7f+o8
sGSojyRfH6RO1d/lq/MaGPrAqRsfvIvqYkXhuKAdBiXSSk0FiEuLcLnxsLIWvNuw/VrHtqUFoeWN
2Y0+ICvW2oVPUAvx+5FUE+CpO+vmBOGRDi2f9sE2Ckr6rnlWcNOoOE/5imeysb9QRK+0d+c93n0E
qX2X7x3INQj9HMRHkxsGA5MiNLY8RLkF52CZL+8qULiIg4M4yn+Q67TsAVKYGoclPJr0wMr7Ddp/
vlnw/z1JcSIfJfwEZ2sHFHnSDtl1YzSc1t9b2pMsaGSDVp/hX9Y8kytlECbVZ0Up6obNAZ0YemWL
9UEY0gouTqkToNFuchMeFViCP8oFgsfOz+BCm95wuIrhnEWur0gAtTuRwrLJe0tThKbA2TXgtScG
l8q5PWxXfni9fD9Gq+1I+hqIRKtLyRTcyLOGF4ASiKf0n1Qh222ZThJdmZpTTe0J3F6xCDFpTFlE
ovTLyqvZ+Nr2n7VQ+infMxOkeUjlvQOZ8MVE/LJJDtlW6T+vNm44EKSQ2IY5aCrgh0qL0riOkVhy
AWutKK3um/9s0cfyiC2Fmy4MbY96mN3aH8BYKfaS+r4W+OCZa8uTYYFmtP3frQqTmjePpM0djHg9
Vs70YpVIU2pNq9Ev04V8iPdNbtkSAiCTp4q56g6eqsbUqbQQoW0R1jrlCWzyUlIiRCjzhwQkIgOQ
tzUWsTctQVY9jRVSOS+4bH21bssb74CuCNgTCiOFk7zw6mtz0CG9YUEf4CEr/KR/VFR/MrR8yg4H
zleAGIHXab1Dv9kEBaB+aJBmn4E2cypRlitV6/6DN13qjKjv23xPuTmkiXV2paLlYQqk9zCOqanp
MD0/1iyygPqWDJtJ0GZmVerdX5sqAGRa7FmBbkRoLBQQ2j6arMfUmKnb3q7Bn9yfzZZkwTJTXW3n
+xbzkUmZrHxyga4WgtoToPWklKEUNHzGP/wjGgrRWW+61BVhAOq9ebtqJMCZAOCOhgXLVVzzBksk
z0zh6ScndNZBNFHtjA6PgXfg5EYzqzkxKbH0ciPEjIzbGQ/sWabITdULcaPe2mOdxu83UzsHjEtV
o75hBrtwiHC0ph4f1+MRRgg+jkMvUIvR2t5fk8GoZJVHunGiP9x8gKD7hD2a0dcqaJJdFO8s2nLa
EVDTc59e6M0TmrGQuaV6SApQTxKER6AOZLndfTDjHuebHxYebB6tVCn6vold5mSaS36Wjq5Io8rw
geEtMQ3iRThdketQdgXaCD37hWMXZsa72kG2xws0PpSrqR4z8/GAz/okAJdxZQdOl5DFc7Z3ISrD
FGQt+yBd3egnXwD+wTEZzGuZwga4VKrtSA+ceaWGGfodttht+zRzpVlarHN0Z6Os72Fa7cRwcYem
7iPD1ujCX7vXRbUBsQEFDeYg9tGYlcCVEyWzJi27d3KtgDefj1841MdJmbiwc+UGWfKCES1feyOa
PQxvLQvBFTqDikg2wLxC/GDxGpW43Dapf6rNHzckx7Jysz0aN/BB/6s5649Qr8rwLP4gUGb71e8z
tNn1H9PdTJROO/SRX9VmJzaJWK9unTbVuwR2lFPhXssw+VzyWX4WUxH2uvzGZGuLgRlHF4Q117Ud
QPdZ750wP3ASyxKIe2QSYfBb4EMjJZO1RtkKc7IcDbxUIW9wI4fiEFw27HO1AWl2xkMbkrt5rr5R
IeYOSTKVPQDOM+pn60RxvZ/hExeveEHc+DewIyuG6gTIO3gEZa7d3ub5XcBy2nZi84mB9zuAIf65
43DLGr0tKk+mnFpn9QuEDUIaCvnhaT6RENoGqgoOY/PL4d4dQFRYuOREYqRQkQImNmXk7ZiLayfu
KjOjSHkr7RmKhuyI6CO+P4KuhrSj+MAXgvDwLaTZe2q2mVKwlx4SJQYE9a3+dkgKbr0X3jfX6sVo
aVHR1iX1LQFLHFSXbv2XZgCAR8BvVFeG2C4h4WFPrM3dBhB5sCipk4tdz3GCKLcH+7eHlzOOD6GE
vzH8Ew9BWfm+G00+wsx7MyI/+RoDgG/txMaojuuO/ohdYPAk2KoE3pNZiK1D+05hrCvinU4IRl8W
gCUo442ZciFrfjkNWH5lGywHZ8O6IpcTTigjMfsazhnCrSqQM4yDBS1NC5qqtPcCPPBqMXgxjm6O
yHyJRP3uASrAmPWaFLQHXYm5nj5JXCv4H+nb03PHQ47Mh2PW2UhRhd4j5cPjxWj2Z7ug0s3Nf6q5
MN7Q5xQ9Nh8DLNfOdronkbUvPPmnMb7gZTnZew3KI/hFqgAGrT1Zm9X2HssBiLqtHbOV00xFWuFG
F2+lR7HiTXT1T2C5Jf+LkBWJPDMo/j58iUCCYXNpwKueTBqf1OmkrbKMnQ3SpnfawZK+2SZ8qjU3
XsKlYCWhOxgpNGKUIAcpDjxSLsAqTxG06kbOBvCnvGfOVMxIvy7DOYZxix1qrhERv5eEWCKl+Cog
k2s7Wnydmp81qpBArBCnlIybkxajwFv6RvXdZCmC6hSeyxzOzQctXtTb/QBgTttTF3KKclbgUmf4
kMmAXAkMj+g6gl8fBIz1ghq/uQBmrkoqqusZU2MSqFrLmKDpfbnExDjSO6Ybg4N+Oi6zELCYlhfj
dPW/hvwUJIliXZgsatLGDX/JZlp4x6AQK5wl8Ae3n0pCXCwPv/xh79hEHhHiSGCT+P5b8ImxwRWp
oUTQ7wzeiWuoQaNHzIoNU9oXQ2eTr0nr2IBoGra4+PgLkoARIRzSLZdEuKxtRVAfP02jidbLf7Ks
FzzH7gBm14wiQ1dqqLwi6amvXFBUyDsYMDGWkYuixYCbFTfSefAyIsO9VuBdk55zzmyDsMCOi/fX
bdYtLe0p8tNsgpmtt3vxe9n1pm7+rttrQYjfzl1C1B2F2Ak+gI1nQuFwDG1t/NcrPTg48pMl9/uZ
OPlNfa/fZNWsXH+twSG3R480X0ohXrb6zCr/rkyrNKqQwuhkU0MTc3QGD597m2ujAMSPsQ5V1cwh
g9hcL24trCcPrUpL/bWJe9FWFSv8wRxVVouKAX6dltcWNJOapU3c0O3CbzMHLkfz4dJ0zFpzcugX
LF/wmdn8M3GcQhWB7sLuuSBYx//pTDsdFAsYwLixsikBKe97Y7CPG0AUSbhAt0zYSIi+5prVZIyp
7dPaCYPrd+IiARnw0lu1eqLgH2Ii4RVY1xwPbmEkzGc/thzBSDAXnUubz9xvgXnizy64Oqx7P0ku
JnDzOyUx+8ECP6fcBGspqsWjav8BHbdt23x03No2gZ1/HOMmVD6ly4RsHig37SXn/wetzIdgvK7N
tH46xwsEgjruXCCpy304LSVYExYyMMVOij0hXLbLkB76LXXM2RixJh/x65B+S2irqL3v27ROmaLr
AUOLr4D54o1bsK++bnXdOVQr17sfcufN+yMwe95q3A2b//2HcTva021WMJ15bCSqbzpCw1aRhJtr
+MWEMCWTxVnTvUbf/VU1jGyHC03mIUWSjMey1VJR5hL+iJ8z75Qhgqk9jHqDDE5YCDxZxXJjb14V
lmVj6NnRcL/1DY070PnE9WDipr61YRTh8a/pYuo5DT/t1yfcBTIDZ5yPSJkrdbUyM0MeksMJq5FX
913DeQZpQetyRmppRd2aZD6iA0ZkIk6DfD11Lx+hlW0NDm1udVV7B4LHnf4a7ofi27h3MX+Z7rVO
cLdYp2h5ucm2oK0nYsyRtpv/nSRWv8r77YT+/AZzV9FyLZ3EaXhYFOD+jnjdad2cHuv4zWz2KucH
Q1g5qwsfSQDHmtDj4BjbJ5623ruYw+Hno8CUY8RaoxBfk0XpxTqNTfutat7Z8wXpKe/PVgvf5FOa
guqX5mX/25FAHSniU9vZghv80GAr8YR5e7D/y0gnaVCJAC/DqPZmKSIVjlofSWocDZti9YakLV0b
1bQJ0ohJoIE7jdOl+BcuykQTECEUEoBxKaYDSxBAA6LeJ1vN8ehN6UnzdfFpgVyoMHJIPosVLyPe
nQyxvALj2Gqu2NHE7dx5TINAUZZAyzXTkRKM+jY3P9G+ZMvHafT2UVVElVibNKXIvsX/Vrfk1x7f
7GPuHVzqf3cx03n0PHyfyNjpgWFp+K/YOndoda6gjsVZnSTsqkurwsmVk1MerAqOM9euA18jlIvR
ExH/ihZWB1hJ+BUt0ieMqfJy4Mfsb7VvUmNONbbqaQXhyXtmz3YrEiq346sclx+SPzmytrwaLIcp
WpEHFDXqfGUUz/5G9528bkHoEIC9HI2OxicOJEzoNo7ml5ceuvOKEHQ9HVOwDP7oMOfQhY7GAUCM
XI3sK6jZtNbLAQv4LwjNp4lBKUI2aV2GMQpwY9JmGFlHcyKzmJ1HpzsgCTO8YtLjJFVA5Nuzczfn
MuC2MzXShLqdU10/D78LSCawNpBOw+5Y/FfB0vXcQyAZR6u9/ohSCiH2GRSvsJai/R1YkS62bkXD
9sxozgGISx5uKUAwV7sQYWuoPWy+k1JI5Tx7GlwxCnti1rMPgvF9NKQbAiILQwzjomWzI2HeJqDI
cyHpKSLHEJHvipfRtm0PboYS3v1T4+Y805hOnMwCrrLGGIRAeewhtLHOG0oCo5+FKQOSuLBWkLpB
mqDtPbYrrBkxtvHSWu2Glq5mZWIKwA0KZfwm8NN6nd2vvkPBQouHeFvq7jf2wexuf1b+jZY47N4r
KeXGaI/CnKAqXqAtoVvOUyp512iTfbDpG/w9ct7JlAcl48M6iW/x43a7zNO6sTzO+9A86P1eVmmX
Y2jzbaGAdEIOc033pUxfOm33AHIsB9DvxjVOwx9OD7ORGj0k3EWIIAmwvsgIMZOfTGHdb5SjSo4N
DTtWvRR4nVOt/VchzU6wyHdpi78lBHxhHPsrFLJKsqWSmyi4N8LnO6yittWWLDZPRmWOLOzcgcK1
OBGCMpiJBUZYxEw3hpDNaxXAeJM9eQq/yGcFk03vincg85RZqL4WlV1C6A77E2jf5PIhRXyYMbjh
KrhPdllKSrRVW0V0EZvWhGGoy2mdRDKR0KobcBE8g9WnHPq1hdPM/7T3fz1cTNINPSNtBGAXS46t
9uznPx4ysrPkIuC3uH6nNhJQrqGmusiMoSfuPRaRV+Q46KJxR9gISXYunUARGRnsmRi3sSEFxztD
M+Aom26+yMBv+dskkFb0+E1oxFEhif9oNoipcDgS1mSc44QilWqGlcCzjDNWxM3VqRqINgmtSEFY
IPLGtJtLNAzaZzp/K4TwzqqkWSf01tBkZikmilLJAXncFFjTmvi1NynrODChAvTszIqFR1L6OFge
f7G8QBKz6pVehan5Xy5BrjATBCJw3OZsPsFhfPClwthlAP9ISmThP/G/YuC2yJ7xGPONzS/mmByw
D7K+KZiMSbOyKluWfNhEGd/ZTmbnmmpMbrIhyTvYrbtJLNtrHYPN39re+LH2P8/Nr1KhrpwJqFdE
PiD73bQbXezWE8JU4SJfZtFh6MI+ns6rFfGFKJMH/fkyp8pMWBhFBma9Qu6bRQwDFQK3uW2z3gbz
7zdR91yQHGHvMnDaQj2MPOceZuWneAELrr+hs4esx5KD/sm9kUjWvRSVoUqZqXCF6cjX7wnEpvXK
23OLdsUftWlWZ0nDR1DfUrfDGkaj/56R10peSe2nv6KpePHuDWJGDS4N9DhG5U+PfxMKIbGi22E/
twEUwMaX1Nf2LumXZHu89reu3oKz+Y3Zr7wQYRWm2/KTFgOfYidCFdM/DtMSU4srOwF0ifTms/O9
bHLSHD4s0HD1F7kpZmmgz21XK/dtZD/MdiyFDRolsStWFwywElJiJgD99VWxmIdKa4rK4OIkBwcY
UFE4jN2/60qswrYQG8c7tM/Fzkov5yEcs5PG1hub08a5IUzSms55U6iIQ+VKOKOhhrtDUayCwm2D
WWfoQjn2glTy7fdy0g6+wqWO7Ikq8RxjVAkbRfJY86sccQ3GtcqMak14D0jUk3M3+t19ibiTTStC
nDIqnC7oXP8jvegz3f3p0aZ1RvQH0PP+Z2p9N2bGAxvdO9i6zKIJcICQS5qHXO+xSvzLVF/GSE1R
P9UYJ9YMXWjv9QzTdg94I/HpLV1A9pVyzXCWzNKDmOevn6Mh0Uo9O47Cub7kLb1PkTSq6nUflHuz
XBN2YQp6PpQgOCX8sC4MRAttwJqSHVAjp6auTXk9ld+h5LuVtWYYrtEHl1MTH4FUuOsWZxE9Hn4a
4JNtvQL0lxL1uu3aqncaOFjY4QCXGgovDKFXyyPgOtUJ2mFaYbZoVXl+uYff7UMFd7ebcN7e2fxL
UQ4+lAJgCkOYib3HoFnV9M6kHa3VF38DLw9IvcHODQkAj2X6rd+6kJXAE4uS7pLpYxS2HVEx4Swx
Q0u/kNtpbHEC1+/w4MLagJZeSsgiDKAlphHrDWeSqydWjLQQGmR6rnj3pE+gLjeLsdGpBERX9m4K
sAWpZ4+yZBQNp8lqtEEh5d5in6QQtLYKvpIIg/PwuMUQtu8qDRqGX1wt3k8Y960yIjidPYuUYliE
rb45Hr729xgAMbKc46xDhRSKBcRkVW4bJgbE4j1Gh0sQm7H7ToGTYcox7lC9STk68tNPfh+8wriz
u+4bFRNUR2gxisfUOvFufIQHbaibI4vI9tUC3ci5dhE1hTUqwyR6MO+641uUxcsDvNcvEGGqClgC
NHxZyZEpg/98prRajjIyg0OcsP3qLy4nfd+qFwjfBaSstasAFjKqfzuB0j4F5qeasP0SyfQ6Vqb3
1WiRHYhTR5CwwYZhrpZ0TkijzLCHtpIK/EBEA3gxCEvWCpNZKqB+34j8j927PoeCydWCvNaIFEUe
YsDH01HXR5p+1qb0ZfhEHCnBlLhK/lz29DgADQZ6Mdt4d8fOPlpcDSvW3Ct/B7FLQFnWDoPBkjM8
x1IIAEwgFFojFE4wQTssYY9fKWsGRELOO20SqRKrE05jOeNAXUGtgxbSoFmEt4T9i6aGk3GrEa+7
f7ZKZw7PMWQEn4XP2c5NauwfCXk9QiZB6QH3In/s+f/1hcEOyJd5Vtn89VV6MKVy6GEgtjgLjhOJ
uDEw1XkN5VmDlp5nb5Bp0fAt/5ACEbLPRGfGg+T27T9LGBIWjW6KVNqAoCHOpLycuKoHoNTpPF0+
DxVs0/kHsKIxyl67wWzs5a/ItfA8sVYOXV5Mxvmb+tLvONmxFRhiUN/wLUDW9DeEB2GG3QhMIJil
S3dkQ1Tvh3qRib4fc1gz1sv4USrZPNYxw4p+bwRQXDc6V6zTi1KEDjprgGOPmi5zFnQjzUd9uJS2
pT2gJa99lJNLfceBDBGyPTB/hLEykQAgnnxNhvuXu3FcHvoO44YCgZZLQZN+GNK8vb3I4VQlJESe
QzOlsCVbheEFArcUWJ8vwLbs3RYNooSE81Zb4jmzVFRFg2nbBTF2qXLnQ7OBIDVFw1QWYq3QUwDh
EStmNKd1rMio67FWjk4l7c2izi5F6dH+UNQ7l6wPEno5uA3XqapbyWQnoYJayex47X3PzvLXpqe3
vstoutTP44ld4GutIqATXY3ZYPcPTMEBbm3onI45IIYvKrpblZZcb9ldgFl67eOz0BEUhAR7OZeF
tMLkzPY1LClBrID5Gw1WS+L6fNAcAxHFD0SEGhGdC/FFQ66EJm9+cchCGlVdMOzt3bb2AfnjOXcV
rBIhFm1imMLDGOezz6z6DERQlpHniZuFRwkV4RQmc5sYfCo8zw/tI0ziH8+wC4K9pF5CjdWVjDSY
B+d7ai679FjSD9z6Z/2Aygzre+AOJDT2jAewVOXV+esrTs0Nr3H5BLeRJMGM+HY1OUOVvD2Xb3oh
WtZaPMpddZvbtJZKNRnmUYJSpXw9tQj52ILiYK9Co0FZMgWVofY521mPYdW8vitpSV554wpwyLHT
Jsuei3KB14466gH4ZiUsfkG7aZbcI0ebZ8OYu03YMYJL2WO9YH0LD2/OgNfRPO0Uhyp/4AzgoNAT
R9oN55WWijrBPssHMTspIoUzNE8x8YABeqhWIU2aUfxq4v18XPW/LEYm4B3+MibtFdL1D4Jb33RM
S/mtVobaA3YYSNksUbISvuCUp0fw6G82pQJPRCmmCENpBPJQ8nHHJsFt3tNRC06gyP6eGSjihfSI
T1zsuLnk9G73zL0n0nsMJdPcJsag7jrtLacTLKKRFCCvUXa5gQ0B5w4q+V1mjjZvnm9IbWvLRXO/
2zU0nKiPm3mZWyoUla3wWqMo4l089aSAY2q9fzAW012BPhAMw9C0sGlGYGxjZy7M/xjOpPkKUUNV
sIV6yfh4eTIYNTcYNXOGIJo4o9tE2rOg2kVhjHbWGp9BO8IZWmCJbzLILd/zbIGYHbE9ZjlDxzW9
wIGjEb20duG2yZsP4qMgjxB00jo5JBjbeWaDMHoVC/CWVI1emIXpuNR+4zL1tMqXhKLWHipyZtgz
4qf6N/+7aVWADlSfQyYqSEDt3ZKNSSXs64S/kHGScBV20c3e8+ECkG29x1YQrji+zHa2AMrNZkVB
YTj8ocz5t7nF8K6hlSWxLhJphhEbOgrytkhT956GUkPyQIyumaCoSQWHdAggS/J25IGcdebXmj0a
2THqr5DVTWuxq9OL5bCBSa3PCVAqzhkv+y9EIjNxIGZ+R/ArE4CnaWFiJ3Q4fuEl840Gq7CO0Au0
qW76E18G5fB32aPB2BUrOZX7OJUeEiOY/KrAoR8l8hZ+nNqRFj/bIVSjDg1NCBf6G4707RbJPsPF
DLqmHEYa3WYoXrHR/VzCbiLo534y6xaSHzz3EY45HDnBMjbIZO8GQXCEHHc7e0jb/98RZTGtWKOG
7UQPpzBWPGFUxSfUophG8aZG2QskCp4gT8+5I4t1RekfvfSkQrF53KJRyR0ZLBW4E6XbpJmddvhX
sR5Aw8MX66maRZJoRlRaTb+/7tDcZ7fdM9x9J0WGcjrQyog69GeLIXDurrSzZ1ydmtx7nOQqbhUE
HwNx0W3oX/Imlc0ZSZw0Cr3xFyBGHHOMrcMOkYng+4hKU9PLVTfFXsPo+2qBZaVnIGLzG9FtVKfI
bPEyC8hCPPmzMEHOFTMPpqu77rzzt2bgf6zc+zLU1354nJJigjdAhORDywoWJLezS9Uam45e3b/e
MdXeTzqMAa1eicpHPLByFPUs+QCjMZAlTcVyAFE154njJPlKzrvKCnIIW++IOjjHUknDSkDK9VmM
B2WoFhHeaQhOh3tUxswSaLsdB8WPtoQrvQPLOiWWYgFNb5djW6kzHjZQh1onxjZkE5vPhp+F+RLs
J/H9/zc4J9B0aPC8SKBo4axs4OohUFnVjSUliRqsAHqVesyp452/2/AuF3fpj589WjW67mLbuGFo
T9IIEVP9cqIf5EzYg/8NXb6rGTAnBysBBrMtSXO8DZA4zpvPXq5LZUDWejwZ1/5DY7/FpaSry4ea
qZvxPg2SRUY6YET6tG6D64UFTwvpcsR71kxrl91ekDIl3j6awFuSYqNwz8UOV9oVU4B65BfgRnFy
wESqMyfWHGlCZ4AL6tIBx3wOTt5JtTh+FQf01j5dpjBtS4AKIZc/iqtZ70kW12lPWXS6JvmRZFDe
JiMD7ebchTZkphkhqepB8MjxAr+dSUOjd/FITbd+EMj0IFn4ZbNK75MBHtZCrxL98yAw6abADYV2
Zc/RxE0m3e7i7CVLaol2PSKHlAlKta0pplw6+5i1vxEgYRz3NVufnoOCdz29zDT+i8XHjnPbZ4Nf
srgZcGGdTnp7DS68dhWlNrbUUQ4yoiSwINx9r8LRYsCunylMNJSxKQOzexe/TeNJXGpGaOmtRiqh
gOkkYAxvehz7A2c5IppPBBfBdPfJuJVMOewYE3Cx9+REcpyfA9GH1/p1r7wVT52PG0LCDFlMmumF
iU7ZOKcaNckJSOwTJMJSpYD/xsGPivGHMnZRQ0NLuxZT2ANI04SZL6bZu0K4M1Os51dYoPFnmGBS
uwbd5Ua/Na7oV2k5tyOPIw6p2yeydZHcURIqY4BM3o02JXu7ZUf/K2PpUIzE+m4QcdtZs8onCghR
H2nbEAdMh9Hb4WFHYBPZMjBoT9HdUrivNo1hcuGMWG3Ego091K7Gl+5zqJO3HI9EwFtTrQjw+LXG
ulvUbpPHCMTmq0dCrMNyxXXd25v+saGAGpbFtFoBEZYtaE/DFK0PGxw0yLMVLOQ0r8lId7FdAJ4d
Gnf67T1iL2ddu9OOvlMOUVpXWvQO74LsueYtJ0+AeY7+/xbx6k/nuKakq23wNVK612/Y/h9yYsU6
bWwH8Qa4E5PXnnUDQPLTTi4cMuagDKoUkqhpLEPXA2efnVa5uMt4i2w25Iqk9yp+oGu5eAx5jDLQ
v0S7fViXg21Mzfb3ZZAthQvwgw08sdXxXU8LDbSt/MQb2J24B9PWd8Aymd+jXRKbEZW5JmdEq9sE
sZHyBN1nNwLsr6SfiT7BVV8tDQd+EH/zdVbJi7YpjRCRsbQa+lEnUzcqqujLEJ5Np559xXke83NO
Uy4zidyAObkDZr2BUNqMH1qoHnHv+mhceFcVpjfseRfS/xsHFhaVhURrFoCjLf4MLX2Az8FZo5xk
0VuEvMRuytDAbkIJHA90CbaWWs3k6nkO3z0wHIzcUfkPFBQX4YvzTWcvHpksyWtmiA255xAzsT+H
jCjXejGU6gXBKxq5qEl/fws3RaCwxFz7tNTYTlVRv82C4SLUygada1aScmcqjXVEdjcHBLkwbwIM
3TMwLBqeWYAHPQHy/dwuSAFbLneXAdceDZsInfaiZKKRlWdRmlfyL0GTDJEgvhJn4vR6KFlXPJxz
obt5bZTJPbVKPD2XoeCMeA2Dl/Xw9s7s6F1Wzknp+zVfg5T5sy8TIywA8WB6G9xLBWxR3Y3okIBp
SdeO/TD+sL2zN7r/Nt8Hi1q0t+uETWzJNKKIaA5OEVImOoCg8x7DGlp929Sl0n4mEIddoEEbIU/t
0bAq4CO/K3O0VXklcsxwhzx2hK1kfl5P/CkyRpusLqxX9BXjjQ5GPrB/AShfJMtc7O7cZFQemySG
nbc5p873KUZq8T5cauBGkzQV2XhwaeYxwCjwRWxMjoF3OTRPbJc5HdaCvzybAtkiVcRqQtw+QpOs
IpJb3DSy1+S3tM0ONoK+ghZB45cH0XLS57JRtlaSJSUMg+OKVmDSEQdNw2x+iB61qMoSOylgfwP/
1FyInW7+j9hVE0xom5keSR17C0TFiUl7mi2FvoThuzZUX0gkax1dRj1bGptWXHuQeo4GHzdkmIN+
DGfPDZPFHIQHWVOZPWPAdR7lKP16/AJDkNwNqY6oMJyIM+M4dW3d/rvx+7oODBxbGCrLkbJrw6F2
IEKx028DqFS48T3xyFNKZ2/MkNTdFXz+GXAYlQQlRCi1S1ISz+O/65OCL3x4vbJG3EOLsOL0tPe8
9oWpJJQUOwrxiyAYfG+2MzuoWh42VBqNEFRumMexFp3dIndRCle6b/1enKnaQaCRh6ZHJdlsbqmk
ehaZxN7euuOICv4Siz3GbsCk3giUEsla5tsnTihIszCwmpfKBYMbx0BPyNukzCGdz/597xm7dIka
uXpl3hsNbph10AZHQbariK12hyZkUXZXbCLx4jYUaE7OR/Fo8cN3vQIZsUl20+gpR4/dMu6bgmPK
9LRY626TSnjB0hnPj1Ta7e4RGAEz5vS3JfhOeXGn5qAV86Q6wDys2/06PExdwU941bJegE4ZKajk
c20bR95RMx67NvMKsKvwtczBKAGE4NnbO8fgGJgHS/Rz/xa0Z+nNhQ7k3QJaPptwGsjIeYGwadxK
NrX8Eq9YrNfUk6kC2s325qKBrs3XOcSbHrgPPYxhBcgPOb8QKBmDFhlPjG4wqdjdIlwzNsr9vRkj
mV+CRJ58pRTEeYwheIWlOmy+pmnjhngLgHhiSa56m8br2gGJ45TQPOZ9OZohL8JbGbiXwdCKuhut
NpUkq22Xmy2xmyKxtHOLtWoGzISJv4xwsrRaD4fCjoJL49Qn/PmdfeUoBT3k+1mjc8FTIwO9+Zbs
bwFcvVdokIhNJsGjNjdJ0xMK4PnRe/YZ51wKXt5C11QaWlX8gZq5ba+paBXAeVAYrnytglil4824
nIeXUT2SEjsWtnw3MBaI3ktcMkm3iDt5zCncUypocaWAGBPlcUaQzAf9hX9yO/Qj96cK6JL7ZjDC
DYN+wA9ZcIGzbrK952AwIioGMnW0EgfytNek6dMO7D99RbKX7D0YGXWKIhaeuHIJyrLmgefr2THu
GtD2s152YZ7fnbpOuodBgnHVGO2HTo1E3hj+hF5TxfF2qeCC/3EryPiJR66Q3AJXQ1iF7+HkrGT+
03LtADiyl7FduPnu6hmFyRUea+dL/ZqM6ygoHVCCb6qtflFct8QFDz/tR0vn4ZVOMlXhRGle7WuO
zLHozU4hNq3GOwRfX6BryvNVnl3cAa9iJ1fumlQNxbgoHWSVFMPEE1t2WWC6sz3/GBQ0Ww8byOMz
hyDloYaaWoXfd4k5lTDKypaT3pmWAKuy2s5pclv8SQCJLu7vzPT5/qX/QttZ4rK4Z/4J+vQwL812
P9Ldjsuz/H47OgHVRX5pDGEROQiz2P6T7cM0HMiZ9ud/Q1p2doTTYu4UJNefGP+yFUmIEh1ozrrf
z3wVp5NF+ue6plYZ4VxgQv3XEHoW1mAukwmiDmzZBonT8SHKvhtlRvR6NYLMi62wMLpqP+3K1fw5
9h6ucDJBzCz2/Cvke2CqQGoH2+rliSofsLFiOUXz2n2C+k4ord+hl5YcaszK9VrwjQpRBiNP8INs
0hsbD0iMHH2YkLRyftvrqZxr8AVFe9MAbzziJyFYaa842ukJFXBzXZWdoL+aahJHAmnJmM5Abh+n
5fdT5J1K3XDaW+S+uIrMkM2VC2pTn1niB2wqprVVfGZvRkGJl+FPHcMDLHY+iBupJetEOdIdBIwc
VfDF/TnUHgLuL4EamJ4XrnLTrGID+snv9jgFi/HRdbQbWjiLS3FufL9vH6YzCKwpqlrMpAG+XOLs
ANj4QpyReAmkoZrr0OOfbVDTQvs0H/D0DcK5d7TAaeOUtAwjvd6/fufy7cApxfJys9UmDz9Za0tB
KhD5YgtTCX2G9uJTS3nOhQutEITuZ4DjgGMrIYvy9iuCD+bVh28ZExAyVblfjIL+AjONSsPuE4Ap
AaL47QZG8OapqWbOY6/DpD2OE13yYTX4eLi9qocdxHrEo/2NBc3S7vzQndj1mBac8gJLTVkiffK1
OCSJYqQRO8Kmgt8OhG9oWW2f8xrOyf64jnDYU34OqRx+QMVHSaWoXnxHt+9L/aY9nat93JF1y1ap
Cb/07M76ZVkmGZf62dWAnQl8ntqnBGYzDht5mOtQb6C0SKUPcyr5I6snIRgiEJzja364BaYaFR3v
o5CW/KwaI6dQ/i3hD/IRaul65CykdtanRHMCibeNVybab4WW1T9nT4DUzGlNpXy2w46GZ4oEW/MB
O9kwZmZ6J7eiv49qZy0L++DAdX2qSV9MYF9ty2Bz5Zpfb4VRzcKHYSF3hBpYto6AYu8QW+IBgRI9
5g8t0EfjGSV9Feh4jhmOe600wcIpD7Ik07MpCORlkqHzyvlP8YKINLpMYtgANcsx7vBvGTop2YXd
rEI1hoMEffgS/qHLVG+aExp9vmepGNwzgA8LjC0Xl3LmcfqikplOyvHoFEAeEF0RRbS69lMNMBkJ
8wHBlWHqXGqBGASWN7se7rD5bv14vjZZRcrxaXcJiE9pCnnzZKN6aNjBAMiWqLSY+MFvxjjpFYpY
owROEO4/lILLI+1snZI8E9sI45+mjT2PqHY2T4J/613jEjVJC/hwk+rLF0FAFn7fqfULow5bC8T2
KQvg3oICTTDa/iFOtv02rQfzIggL3hI6U0bURjna2y22P+GCao38Mm3yDXrwX920/g83dm4ZFmm/
aHbRaaKRhaP71MzJ3/C8os/Mint/1BFaWVLiOsYx7ckR3j3WETqyz5/7FtCfNULCheygdUBmvKfv
I0M+r5wvavfApuU4S+Ukeo0u5L02ZGm1itWktT/gOmsJP3m2wTh4U98NgN4QELP7kSFR3UW0OLHr
KlFB8LR+oH4QqHoizKDENQ5t3dOxjrkqxRHwBpomB0Do4L1qI5A07f5z+PnqIH2Q3FAgiIpbEl5o
mJ4pys4hUUpZa41a68/n5QouL85lZZZU4teliHZ2YiDHm1DhtHOtKRxh4yos/BtFaLZWjqdVKDux
gUtfZCkIEOB2VV+DKp9li6VnQNZdJZ5IdnLIBRQ9pnonJ4b+OWsoEojtpEMwvJfGPCGRt9rSrWcg
E9+ENF/kKvH9/hLrMDzj5dtnHzZ1eDfdVnD/7Hg9/r/ZLojnD9oNhkTxwh90+zpkUsODDH9Biz8S
pf36XaDeIIMgwS8mcuk2z6eEcYxzA9JmpGRK3q4fsxsU10OdXHOPmtYOVo98X6M/7m28aD9W+n9P
5PY8jQNfColYfGP1JuEHmZEzKkdID/Xd2E+TVgNIPPnB1MRK6vNhd58ZK+/jX3WTWf3xZG1Nsn1I
H+4Pikm6jwG+HTH/iGsehKpmKHTkXEOsIZsJOE4565Mk1mmv3MDG0aCnXRUX0jNYYo+sbPpqurHS
TLE68JDlD6azoCoeFA67AiigpZ3cu98lRv3jqecBoz8B7IQTfsbgqj8Y2TLDZ0RMWlUeHppf7dSr
EXR1mIXOWhD3S90o2cEVan6Ky3mJTnbztXAUSMkIUpjS1Eu4FZFwIZFTD0zyOK88+Wba6fPAUt8V
dgE40xf9vkHS1ExQTrmeReEcPcl0BXLOOmNjZC7umTwCh+QxZxr3oRp9FSo6ZMIE4uu3lhEQMDzH
yT2fA5JtHFijfyANK+TRmU9iraBE0GWmsg5B2Mylgv/YoGsOtZJU3opNhpuhsUTM0+bLKvFIRC3V
UIMxDLQZ8Ov70+aUsmla0COqp5mKQ89A/y2M2lNMXjEO7RVS0vFE2Emw+gwgYgyW4gRbXDmWT+Ix
oSDvLGuwXBW0d8v0falVLd/qT166GAhmB+xCJv9SQV9fmFwncpcmqOR+Ug3Ygh04iOVLiHx/0LuT
gLO8ndH2Y3F1wsi05WKAcnUk89yRI/4AyBYvfIdTQI1iS/BABAZYiPHVY2OX3c51PiS3q+A2qtJo
EJ6E4z0/cdCjABUsmaEHeQdxr++EH9XDYs06v8z4NdCl9srpslwKm1NhrPf29a2VF0cEnClhArbD
O4C+th+v8w2QkyJbsM/W70d5vsN5xkws5+0fofXaL1bq5JnBJM9Z/RJeJtaWSF6BB8hJxZ0tWMfx
WdLi0Z/1Ze9Nde2wnV6CzBE9jgnCb/Ww13LyVWSYBwnVFrJyKDmyuo6vZec+TtzWBEmws0xhd17P
gr5e0De/652U5Sb3wdsohKRn5wgwE5DGI9Ixt608cykX/YI3sxc/deZYVC0feGbk8iJgn2wEyQwp
Ye6DmGR4ZYhPTBU0UjuLTI6QW42PS0OxZlYW7l/0G5JRI2P0PDkft62fFxAeRyqAuyV9AO3oSpuD
8ynmEl6WChvhVlcrls77GyNq9H8xDcY/XXei5Q6afoAkHg9FRJdfcdxmK6l+iactaQ0NKayFifyV
3Q5WSykR5Wvb0WOQdnBnJQ+uylQglK/iKtrEM25k9CFonJ0PRgsGdQrDxa3A5v03wkALoPQFDIS7
nl4AVNPLjrzBK48DuW+F85iBmauXcIxwUMz8IM5Wgi21/DU92/vPCHC0U9WE/xRWAyH+j3pfoCs9
sH9zOTfuud4fK4qWRg6eUq9LcIA6rLavnaqqWL8aRyvaWsnKAZ0D9LBm9iLpLOnR4rSPL2bwP19U
AaUPMvn2VOHrhoUBLZ27WBxatJx/ns8eh31O4dcuyRpkHTdqxOpPkHFuF/jG+8JmHuL36rsDpabg
Uqlq9lQqqKdmcabrTUv1K1md4FzlzaH9X3Z6/+TWKV/PKqjmODfWNv55aDRbgaSbUg0MDbxFoOiV
INIQRuuUyWZCujB0PtIbR8LlkStIRCi572+phXxOgohYietoGB7jV5EGhl/xWWJ4tlUtAvWIJx78
PFc3NoklsorijFboUwCw67gVlC+uZDy5BPdWJN8zdS2HVswxYFjrdYnbWe7jaJJY8PzmkiI8giyV
hcO4L7Z0/j3FhZk2ILrAWKjXiPIPh9NBB3xdIu7xgTSHQ3rU/FJvEskcMdtwGolaSJzo6yySgz9k
RSExBocc4eJpQ95p7Nxerg22zZl4TwyFNmwcMZb6SIfuv/4RwRlmIVG/FNuNJFMnq4yoV4uN905u
hgAr2VpcN2383TB2bd46pEv+9IUmkNZwywW+/OYZLJF100MqPFWAWlY8SaYMHk8XhLrnnx+nY0JS
sNrhGBGrz+mL/O8Vri/PQlXjMO5CCW1KVUZSHHDwS+dwDImcvSnZ5N5iYgP5CdI9ZUCfobNloxAr
uJBfaK2zkTOxF+HtCksrLE/jyep7cOEx63loRKO2IOmIiIS63YSxepckNk0Sl347hH1EsaLaRkNT
OmjzE3LthcIoWiXa04VY8dfaBKTAwnuZPNOabY79+fJ+Imq0UPrbRlT0LtZTR49+evAcm3LPrNg2
tzrJsPIvimOUBgZMOT6v0c1pI7w2sbuRjtGwXCPY0kk9WSjezo+2C1d3S/TtxVAUgA5k8eV7/qsF
qm7uAdrf3qRBVaYKaF72A79fFGOzEehkooeVESETv4+qHd59yB3K/P0KeVw1fZcTWT3VhsMA1azN
fu/SWkRWyMsKhDaNb5OSExbxW6BpTadVhBOtiSLMabsgfQo1zNdLWNa96QBp/QMWQj7Cog3I7vwh
jGBepP6Xag3yTu303TRc3eetBzhBcvoh+QupnWFeaN5ZBjsjYLjc5zWU5abiltaC8Z39lts7Bz2F
gUpiczGmtDWJe5SX5saKiR7SVBqlbW7IRxN+aFJbQBxXX+WGtW0eYMpkTDvQp8uneTl2kvNT/KD9
6pVhecukkmabpfJM+1tar3445fJf63k9QN6L5VPn1ZfpdExvRObFU1k/vkiCIOcQbyM4dBl8COQe
nHqBUx56UCOi9ZLC6A0KQZD5++Hj7UIR+hPOJkj2uGyiM3QQybK9N9TfFzHP8WZ/dM8cfHucUCVe
6cvtNhmr8KAVuT7ZI9ALpqPSUHZasB+UHSxrDTvvqPlEziBmi5y7ct0PzTFJymALWRygi6Bb1td8
iUfseL3j7R/sqi6jYZkCTspLVLfKPumyoo2UfR7k4gP7/P3k9GMcsn5srAgEAVx8Oh7jtLgkI0SW
hgs00vNgnUr8cLMnG/XvPIXU8my+YVEDCdfe4QwJ1r6HNm0uoha3DXmmLqi3ik9UKcjn+D6T2Bsw
yeBFUE7T47JjxuWd87ZzH6RPkUkdCXT050Y+CKOcftuFENSBLtB6mHrs94PNibILkpBdWdolBh1S
jX1UVEyGu4Zc/uP+VVY7N1XlsLfVq3gwyJGLcblDgelRqQORDf+63EnaJ7dzjPnb65bYjG5fASfD
GZxq80tuT8WKGpzcsqlxcIj/GJNnvK+Bb0+qVxXbzDQbdySyd/V9XmjFeM+YryACcy+zEvAmO+wi
r7ul9Iu0DXcPIFSXnN/5+2DDevHvigLSt1W4nFsKRcWW969RRONUbnY67anSupXIdVlSJDp03+Va
1Cnfem+YI0vid9xbEzxyMx9251ekmxD+i3fsPzUlpdLgYreDMy64TQt8jHn9FAol5ZakmJBI0VIr
PEbbShiVO++bbg7MkZSsIvsKne6Vb34SGRfiUZQMATUtcupx1Zg7S7GU1Mdnft5oUQQ3M5qvehBF
XfQitjOeRzXf8AIho48GDTecVdP/tkxeble+lfd4TxtX/Pgqs1+Xjw9Rza070PqKduNXMU24IU+7
/8jtffLk8s1O/NduAuQEGJ7wzNSANr2tm9eN657404PZHqA9/3NMUMDfEHpjNjGJ8WzkxYo3Cd5s
Ibu0/DW4iU48zjslX6JwPV9q2hZANTaOPR5rica2R7ync7w74BmoQScJS8pZPfcL5pESLICPAnFD
AJL9JdWhj5MhjtkdAixFfuHvCz/qNsDU7C6tANOWfs0MbpBvAaatro9IFHyUvooxs3c9RbG73kz/
B4Ok47yT0vyebf/eRzn+sUyKk7wVBqy0tlQfpyKxaDCe/gjGgrjFylBvg4H6t0nNAeoe8/Xse5MP
pSSNrybB4W4z3OAQuoApZI4esVUb8CGf26TI2qvvcKEgU1Hvm7YUlgZKuPvunYH1dPYid44Kb4uJ
PytJQUWgRhPbKfqcS6rSTswamuDUnEuGPFSzO7wauwkvO25I4RvngqybY6qvtb+8EDke8Bfds3U1
/a+5qoc6+uFva7+mpCCJHsZ+qzkXmINoj4b9PTfbtIZ3hTN4VTGQ8GIrppHv0go76qJrXkG+vvvh
31EqhX9ZzHI2F3eHnYgTc7AnA7KUU9fc4Qui4VSTmdmvfSIolbQaiGw+iIFKQ8U7JL+ZB+v+Sqvx
L7DjsNrpS8ObMyLwKNM2ZQ3YEsCrYfRsccL2x9OEeMYsQlf38W1G0wXYY6OhEgyc1y2WhGVEVokC
HLs4MsfGWnlaRj4Txg99t5UL5qlyLtDbdURW7xgIfrqdFTnCQEbQoASFyt6HuyuVRH04Q+ycz8wF
M7lXB0hwvStT3Kw7FzrJp1fJ8OiAmQY7oQl+bBcfc+l4RXkx6JrL1dI2pY+i5Zkbw6NpCHfgIAcW
30XiMqYampr23Gxc/8NdsNW6KoWX08AWG4xgF+UsoeYqOAI3nF+Z0bIxG/cZNmiVOTKGrU2GfV8m
NVTsnZ/1w5jHNKxvaIYbG/HhA2+8MFqXaa0J3dtibEDPHVpKE0RMxT+6SKhBJ+anexflJuwx9K3i
tfPzfnBBYVp12M/UoZg2/V84qgLqKLiHalbFH9PKT7XlwLNw3ibsjdoeGH/7U3KCqElzl4nh26om
L1tBj9e6Zu8pPlHFnrLezfQpcUpMot6Efu46YC7icOUo6iCiFKpUC6TniC5vYiL4sYJkAMKj6oOK
4RhNyKD16nYxHH2Ujs6LfAhUB9CF96rRuJwExO1UjSQzR8LClDekWZl1PUamq+/ygbh+byenZff5
xstDXwTRNoFV72nds57X9aGHzAXb1PYFv6+ZB3ZQtNnFJT6+3pk6slmj/WFwutoEbEhqGcpkrQHc
aMKsJwywne9NuZmHJ3wcgxWj1dVMFE8pFSgUZg+br1NTEY0Te0Djdt0hob4oCwjW79PIfvAOwqZO
xVnOuB1W7WNCVxzSpDojtn1ftUMtMh0ELldu4k1/nFduCp0eCd3UyL3G8lmaPdnlI6hcLDnDVQaW
ZDP205Dvm9WWRJ8cVczmfZe8h/nQmLPDWBDRz+b+n9R83EaOEE5sQGblWmfh0nvSPHnkjxg7yPpy
eHNv2MZybYEpy8tO26ediLQplaOfjdwV5TPD6N0egc4dWIhlic0uTUvvrLZFtEv/dY2psky3ISBQ
tOhFxmfwf4jpmvGP48v1DWX3WLcPLlsifUK9H3TOXM9SNPWUofTx2rX7pSn3t06hQbTUZQz1OBAz
knQI7kmDb92MMYDzikT/I6NdHrsaRX6EFzYRMOco4/XsDn3A8VopJtjRS2DDtv4rl58hWtcwrpTF
5zf1yts6Gop88o08If4a7aq6/8r3Hjr7bj5M7sxeJknIz1SO1RdyNs2Lc8xnGzJstH8SyN37X0BT
UWcikZJAkn57A2AIcP334Mr2RuTLuwlkYVXa7JCc87eUkh6rm64EOwm6cdVXqvFY41CmeRPj/ZUo
8aOCJZJvHREcA1L5p2zQc4vINmO6sJ3JmuzpT3tr8H1lDF69xokHMr0X9Yp7356XZU9dN1Ji4vKI
FEBlb5+0N15aSMR9uv4VpVV5IRgqbxQxf5bmOa1dDIzb5jS6Io9vgP6fagNYCGKu1+YIyFmwCqgX
wJWIS7aTXtPd5aSpSL24ULZB9LBspAbvA4VqwHRy5KDw7o7BaxXrLeYjDUHPp/M/vaDQpMgwmuQS
VUcHfwbHE6c9lh7F261NmXiD/w/x7ZWGEzt7kLmMPbo/QMl9f19iayVZKbzC9xjgNBmYJLXXScu4
67HCx+ovcrothN9C8G4b+l7w3EoYizW2kUAyEQDqJKuOdMkokB+boOCgU82VlnC6Q+r6AHohVrOH
Mb/ejbpRCbHKcNnCPRaWhtfutEsYT6FwNz9BXq2fXEIoLh7hmtcwEW3AZ3LwM9cCcJfUZDtMlEXx
WAEqgEyg8Uij1GMR80xVhuzMt6fRsVDDmZFZJpcCfSTG2Z6Y4n3sCYPFOb4sDv1qzYiYMi4jomPm
9hWuOn1kNOmqbjv0I+RR8qzX1HXYYxOKb6LUxMgyOSfi816OQrmEec/n8+W2V08JVJtVdvZCLqhk
pL7HpKZs3b9QUkDVXdGqhrZw/0T7pHyL36eILAuRrgxQ4+zdOqd8Es/f5ZNTxQpRGzM2A7yPPfOX
98O1n69acaXQPvaliZPUbLMSh24xUobSzCIbFkQ//GTYQF+ua2/bqCwSGONHPKWNs+8TG5FoncsT
ahh8JaGGvcfLyBII2IPb5oWU4VBoZahucr862dodQCm79vE4w1Og3BgfITh5T/5F7NyByL6YJWBh
NFfIzjVCqeRo7aiPd2EZ3icq4bwh/DkSw6a1PQTbAt+hkHrJLw+DdorOZLB9KQfj/AIwlZ/FCb0z
XVax9gmQ0EjfyE6vKgbkk/kNMsXkvYamdfPObyGfAyjVlO5v58hgagdsnvFEjoHOL995GOjtkYOg
qnAEwvBp1izm9Em09d3bEZMVdz8f5dmcinQ0rhM22E5w9f7U5kVsNyO+SGl4TxlKlyRAvf4sAYRp
fHiHSczce2FGR/jR2lysDvI+FIYs+cg9jzdZNKS36k9ECVwLGibQZ1mXaJTkwxzrAzR/xlPmss/T
TwGwm3JJMg1wtOhLfwsaIhKx0+BxZV92T1hUtDWd9xly++gwFm1EYeTRwW+920jVDaNttoiyCqmm
67i7+IdgqldvFHTBHoA5XhFvVSSJGgb246LPMoCw4231cYgDTG3BldEdCwZ9WdpVqCkBtay9k96M
akl0aoN09v/ZwRrOd3P0bhRNhL7FtdhWldu8cc86gJm/eqLJGk8TZigeZWGfAhCHKHxIX6B5MfA9
3A2fxiWTtruNPk64lg0mXiV8BvHPG4Od/cy8u/oZ3fIOh4wpGqG3NOVjIMdcOZNsVzCN+bfZL7oI
bnQL4eWxOjqetSyhzkNZpjguEXpq2oeI/cAs1KHkSomnssWT+KQzdR9+2Gu0PGaXcwow6HqGsicK
UHqr7hgnqIAK5ORC+2tCUtA7asuag1evxG0Ukcv/dsjMFaCvrTEelgG7SZVhohHlKLiFTJVsNN0U
vZv6ZaFwKbkWu3RFMokCVr2voRxR+/xfVwqS/v8WGu6uKl8mPUpThPE/vQ6PwtDwiWkZAUVaVdn6
R8x2zzTdEm+DvPYdhh44U3sEoIDesESK47n9elg2gFVy7MAhPYcI0wbEX9ZgYKLqGJwnWr7r6Xb2
V5FeAOwjjUAnkObTbn3Ik+Iqy9CccN+ZI9yIXaNHe+zm42dWMibrdvBQfJEQ2iSqGRO+hoIE+Z+A
YeiYSBMOTO91Bn71qG8xvtsL+zPVAB/m99oEbCYS13gn3+rdY3umERYy/I4FJlKMiKJpuAK9LIdw
oH908ZFCngpAUWik63QX6E30pzLlkvSEZ2UJmj+VWOxIP9Mxjcg9twssIiBcy3UPCjznwqOeGU8l
a5U7GgKi/OJ6IBKKeN5h70luc6u0tW4GxaU25OdXFcw1fc1IGz3H8VC7miv8W6yrXd9OAlVSlADw
kFpWQSKQ8ZceRyxbzd/ms2TSDoNP2TTgmoG3SiIiIYWBih3WxplbckKOsA75oeNF3jWyhMtCxNgt
AWXmDnShK4HHpUhIo339uQ01WIEjJ3jJPfu4O+/g1S8DrXpQIFnUcMHwR5OK8gznwyW6YMwRL3Kc
YusumauaeBB7Oi3Iln/+dpqUMhR84bEwZH8yjbHE1AjpV3U5BkTmqVlF5roqVE8Ns6IWlvKhEunu
Om9xqr3c8cX3+wbh3tFu1J+hdfAzb5tE0tYJWUdv/16g1lLoWLf8H3Pr67hmaQVSoPbEAkQVq1wB
3G1AsFE01BTSxoc6uSn5JJeftm5ZXHvKI0Xb6VrRiZGhwDnx06vAToDvU9pF7/JJybaXo3dQtT9l
X3Vw/elzG0rgFV3EAbYbauuGNFDESyRlVL68dKAba/JdQn6Guw5z4DMdo0MwD1n6UgNgdCHocBNY
x1WOF0TDrtmz3fnyDtni9I/M66T1cVQXUiO8BzErUFJJBDm4KtFj/bIXRRGcZ5Zq+h7lxyiLCfUX
eqJYuL7KxcRCVpXfb0NenpPwIe22aOIdjAztZcskQp8h8pkQ80cLEH+JD/qaO9yXTtEpLZdgl93/
RyFxyAJMnjU7eij0YqakslOWfePE+WZn44SbRO8XABVztjjyCjVU4+pJuS551TMRPHAjAM40FyWH
WnT56tdUsVeQguICGmaNZkc8cMKZl9G01dH+peRAX+QvCypm0UEYuEaioMq/vxWYdGbzD0TIqaFC
D5Qznm7m4XFcLR3fworUluq8P7XJsqCyMaJBfcrQClt4CHnwLZMNu66o3yfkVGuo7sxhggvFUGDR
XvahY6wHUoQ1LnYjoAcgsZM61pCHnOXVs//zXwq/hYvGurFXYN/jPgw3qnxYF6DIqQPiDFTwWoY+
F1wlOxu1XjqQJhUXRZZ0WB01b9AE2zaXDU5E0iac/RQQZtS8oIgjS0uMN39UE9Io/1joyBVFSvFz
80V7WIbChr1Gozp2lE6kHpCmckEPSjXJm0JF+LSj+9pepRhOpAhDRiTwAl00YfWqiejdmftbay8m
TMh+JXaOLlQp8L1/mqEl7abwMvIQS7PriIkDKVpxzviSPX7ARfQDqHlvvc/eNfQlSCasUXEc542Y
eZLO8Koc8JoSA/1iSiKes/SVqxbZxzCxYB3FgIXcQMQWtahgl5gQGfXIVognA+l5kD9rPlieAOw0
vwRkyoEEpGnJLMWhyP9gfzlUScnsyu0y14cRhTKqKItB7mmG50K7H7u1jD4eLBvoNzqi62t3dPei
HqJ6CRUO8PTK4aoATF3DOzYoUmoavKHIU0jjKr3ZJzNUQtbSXEO5EX3GSn7BkABkoUtz3dK8hZ0t
yxtFtO+ZSUobebehNkbqb20n+VpIJUl7c/+2e5aIjcYJMo5dh+MP6ZvqnouX9vO65YOpBUyYVnjn
7rAJ4IOtT9Qee2Cii1b22Q9MK0CHlO9Dir7rHzp3d8f8YALLKHicnfiQ2RJZ+zjoTIFDwIK8KDc/
dbq3KVIhkNTPnGHSEuHaS/C5OrSF3pWmW74ae3z3bSlL1XdUu3x4wOcJDaAW1fzQjWqC4X1v7vwe
2x/oakED8KQzghdtjrcfHgwjxzmmeVBeAegjysbsnWRY5bYeO9Jg3LOCKDT03MP5cr+KZwVXgd8d
1kvQQUT52GJVOqwcV1YUSkX8xjlGAj3MvcowKVCXtBcgZb3NEiGBu+aJYO6ewK6Wai7kD6TcAM8b
tiSIt607FviHCYpK+lZ/6Y9Ym/OarJiqduP12Lr/Nu4QYyn39XNC6GvxtiwWvLsyrqn0WwduY+RV
+hpUW19pwZSqQFQhE+npsOh1DhTQ2nNfymC4vOtuBfiC4nKZXZNTuVBcGnOng+VdI9pxmq1yDy5c
MEmwbUDLabKDTiaZcLn8utP7Q8mZjsjyFJkwRWVZt6qT19WYjTxCM4sityW/S42g0K5/LhfGT2u5
SbMnH5dyblPvBDuWsxM9LMQCgPvdxKaECPwy81Ttupg2wF0DDwBBph4nDzIZkPjIS/0aY5lhUh/v
SRKi4+Nro9UjkQz1P98Wmr9Jf7aRgBssxc5oiZsvyiR9kwMyFfYQpyqrBMass1FrEJ0WJtdlo5VI
TZK3Ij98ASOU20WWZUo+UL1efI/jAbSrGG8Eel74uLzVll4suczbu6+k6muHjntO+pmkSiH42QvU
zoVx+m6tnpOa2WK03fd9y7dnfdsbDot5V0X7ZQ0DAjhf2Yl86FUml/ISkuGUfyXSIp2dFZahpMHD
+RoErpISwL3X++f/6TEQDNvMY4BoPS3KKRJDYTXsVJ6QLkf0/KFhIkZCgxte2O4+n+pF7e2/11lb
SQJB46An79yqmBgK927zhmiycB21kWWQ8VQom1bq+ExprmPcH312aS1+2RHHVVa9a2TYpbHugIOc
Zmn2bum2mzDjDIOjKsE4FZbfeaGtMt30fCh9F0hdcK9LTB6n5/0OOsvk+0KWRTo4zdlhlTkvFOgA
aXF32FDeusBJZigeZnACAcArXAfPXNIkhE0pbPgkCxteIbtkHRH46YI5MtGDHC6m517mzqEWY/sx
cXRGZ2W5uzE7FuFWoAketl0qAw3A43nfSVqx/YJmZQFmEX1AiyKwcl1Qwnekg6H22R9Nua/S9Ns9
NgJh2+CtAStBClHwGpsKWK1eOhh2jH3Yznp46ZZP2Xxi05/AmzLT4JMAyg4JLrZWeTzoa5vgz/sw
6ztutJvexdAvWII44wa4DQAryLXwSyJNpWp/B/iU7d4Pb7Ao4RoCgF2rBI5PvRGmTuD5SmLn5CCC
nbhriuvh2Bwb0JMaiD/7BqL95h9xjCal9qDnBBn65sUkVRfUTtmDxGuHvXd4pstTIeBc3w/EzJHx
YR24zARZWhN2Rmu2qbT601E+C4m/lOneFodBSXO8MGhb34V6fKnHwF2U1P5hlb7KkN0FUH2LBUo4
fZcImPtNFqlINy7MM6uJBuU+9SBgdZyn2xS1P85gMmvnDHDFWbaOVczgcfvRVBJeTp4Jq7HNvG4v
jeAPjsXnjLUUnbOf6zMSoVewX4HB/twadIlpGWy4mLBdS6Js1ynkP/Nl0icB/rTxyvHM8Kf2TWyZ
jJMjx1l77aqdMwo+1KAeHFK4XL+GxFcNTPFVor8sTcB9GHDP0Z52nfouUWgg2l17DBT46UVQzVTm
GijB9/wm41Lk4ME/V+lO88Bbz1BRkbuuV1Q1AEPvQCHWj2XrD2d9t8QrtQgh3Adpw9gHiNaDBCCw
4B06MNat2ikh1dcJdqaC//LWwUpSWMIaVMYNL46c6ZGYort8QzjRf8Ec8dYbI4C9zS/fKK3pEg/n
hsfy56YTx9aYLZ8ZldnEUIrgaPvtBKt68/U26hYbJ3wglyz3jD2mMbWmcidbgrWG/BZyY1Ytzq+q
PWVJ96stMbaicvTsxfFaLHoAlXbYKqUD15bSaLR7WTyNniDOJdJaYwZm/jtc+TYHDzwthkEooTah
UqaEpTQMrWLDUaNupwq/jK5lIIRXC0GcEk/WrZdddsSc+Dh5qCFBA6ywrmZI5fE7KxLIaB4S44Ua
sdNlneOtfIk8vGJyyY45ztBA6edj8R2RkgPllPYkwgk5nzmtLoua/zhjjg6hsFCrVoBnjn3u5aHc
42KvJxYjhU5Mnew+60aQ1vnCJXRaToA058K3f6KA9JFI472juJQtjXnmB9RcEvel4/hsRFwvkyG1
+0g4ocPsMq7sItIt1nj2KX5lnf87HtR16+hgkSBT3fwLScMFkYdtujb26yZ0xjMYAEfuIuSNkQjY
ZcT4PRE1HUJ3jQrME0V3lq8hS3J2n4nXR8WEkIILI332iGxfdmQwGH1MuJdCGc8By8yy+/749CVV
pnKWbHMHXOaJYOlwZEQt866wM5BH3hFcU0JPeY/1uSPEyayaOMW9ho32mDuwZclo2ikbMzXriyR5
TfC0FYWtIKqPQrHAkvKKJxZzmqU0AJNBe6cb49TrdwSHo8FKQKK5Yn4FhPB/OCm5YWkNHYYnrGjA
EZNFnEur/rhVLtV09ofjhZuIyZq19/e1Z6ptSA4HCypXQy61aGk77/XrKtgXUj9ru6rm8VGn3GcP
JkQvIXI3QfJeIO6lTNM932/GxLA+s261B+yjCpSrWCLN2Tvsnrkrpq/jOiJLr1O9nUNc83mBi/9o
Aj4AaFnS01VF34VLkRhasgY2nBSYzO1vgBb+moHOSNOAy8kNBw23SH51bnIWiya8L8INkli7Ff9a
kph5VCcD1oY+Rti/TKAJ1eACI3I6pwgHYtlZTihiXKb1WBH6CeXjGSVkVp7FHQgYkePckxhYXwnm
cu72EInA8yjmFrd2VgTrpS+bhq4FZx8zKlJGCk/vit/bCur1sbM/vucb68elMy+yKmnflthvWgvP
upt2+57rge9ZjNna0n6cZlcbhfRoRKvCTkbHoVuQKVozYDpTgm0ZWzXnQI6WQhvt7iuV6ht1cYv6
6uW2jX55icMIy8rfNa2rILJT/V5Yc6Q9c0r+CUevEuiHXP5tB8XIlK2K1ivEcLRIInVNr71rVGYM
b9QGF+BS9gP5oLB/9lP0OQcyG5NzRhnTszLm1je0b7OQLc1mfrVWDZ0LTQe8UO7UasvnPPLPy3UQ
z9OvUssypZj5Oyw/emAHl0HoL0BABGHmnnK0aUC+LT8pVahCFDJCmrOjh0F97j9D88hdSpt4MQtE
eKxdyyZtUwZygbZ7ADAfyr2J+iFQ+q2EE0QGrZ2+WjtJ6ipr1HM8DKcniM7qAJpFVJT2/7QBfdIT
4ZFGe6WXy4dhBgeY8BWdZL9zThJC0QSQi3JLpudvj5en4T3NFy27Cn+pRrrgLi9cJqnDcV9yRT1p
QJ9UAJLo+VEq1axWtqsdR1uhvPPVjwx951z+KudZVurQBIZUev1Ajv++j6GfnOdVciPOkqZFXifz
k3SXqxouo8CrEbwMpmDR1S3xmm0b7Q03HRMLoxt1lqPO8sck4LAaNPQQaWsVPO6joN8kvO4aBgXH
PL1WfwHEDUR7mCJgYMb4Rql7Rod10GzBVP7KLJx11V6C6KG2qE4XLSLStsFh3xhz/LBJ/dO/4++T
cHwJP1bDX4Qqw6OxNxFVvFyiPO+d/GsN2wOPGk2m/Ejk+hRACTJ/t7DkOgzEHMD2VU91MmxFbKy6
tvT70BK/lt9VTXemQjjOjua9LG346QTI/HUQmocw3Hf7OMW6kIBkEEHUDF7WB6AuehSa/zyQr9rA
3QQ7xA6dXMUeryfBIHqLzD+uRbfpp078LQGoyeeY+5cRwKQPE/WUARCQQUjkqK5P19+zQLRZH7gN
Jwi11JX0uYsMTp4DVHLBWofCPZL5xlyPcUjcTgyGtCVimbjX8MKnA8g79JnWyb5e6JYRYunN05iN
d+rNDnSz3o224XgHEYjy50Nmb/QTlfg4AHLIBMpLrHoMN9jilSC/2UJbLTaH3kO+i0i5bayh7NJy
cKyNkJaE0BiU4K1Wh3ap4d870D90xFUrrcH24rqDUNLCGndeYL1gyb9Q2Rz/Frej6C81wv+lCTWB
gQ0aN53KtW7spftn1CyrlTAbBiKU8i9Vl3bOEmLEEoZZXPm2yKkAEtaHGFfXrZ9KveCLle4hhsRl
mtkiLCm5mfYduGxOhYi22hexvtWMTHNgxseu1MkRhttSerdh0LKcvlm9Z9v2GCV8GSHIBLHtF1Dc
OL0mlmfC6wUBKoq8MWLotroxJ2c7PG9xvBSBIIvMEEnpZc8THAD8iUGK3V5hNxflSa+XNyVxwVeA
crH0PoiZJTAw6jg49bx4NIn5GRCoMD+hzduoZgUWm+S/67DtLAlwLWiju0HzZFVa3/IIvwflOsR6
0abfI0mWzsYrVv6OwaPWHkJab/tPLnabzY77yXeq3aQuoEtd0ipfLxS+a3U3piwcNrTrDUgaaHan
eS9x4iTBD+51FtXuiVZdWztkwsxv9COrpFlE5GIw8yaTqfpGa/3Covr5XP7HtRLBaNZ3HWGXc4nx
EWSgBEzABlPy4IQ0opvc68lT4neLTdxOEWDCQP4AmkTeMa2geKeiwjzQarGr9UaRALKWra3r0uG3
QbuWB+Pf0BbGXhGSlt1jDqRtEtLMDMNfg+BHHTBRQ5nN+tUEJAgkFWYgQoC1HiSFL9UNnOkFbRna
JRceC9UtieHs31RWADx3G/kf04n4RqMspnn8bCP4CPYUc0OyxKAjXitmyXoE4QHsvFcwiOPOaEkQ
lL/ApxsukfYofRjrEbX3ebhtGSQq+e4PfY8mDcRbbnSolwq5xHyzX7291jSjDhSz9laPkxcGJIh1
enoDKIVG7j+2IxbIGhK+9FoMSvcSZWf2MC2wFTEanBkHEmrxdJaNTwey7PEd0KFUKoMIUeMxC45d
+Vipb5Bvttmh0h0LHwS74fho1X+rI1LttbbOhKxc0vAjSJ9v5UFvLlCLvuCO/Pt/XVVP2KhEj7yK
GmQURPu84lygPV3P3J7nUiJ4m2xgr8jZ8hf6idRpTc25ejo2v9N+kMTQ0Q+XZ73ZR7es4qd0k4hx
u1D+RxxapwHgg+V2izoUz5FWX2QdAGEgOJzps13n7QUGV+aJ8lkUn8X1untCKpCMgZAmmbmciXzb
aM0i+e2GgYp+xO2asr22okFyr7qdl8wsI6bov2TbLg0vdOEgZAaE519hu6bSwPfgPnqbuE5h585Q
qo1WmbgibdSF6wl3Ic/qV7CMzJ/EE6rGQb/d34Cauut1iHjLvIaaKmCGE/oYh1q8XGJiApM/seGA
LStMfRvonWoRJgtQFuuWL/wIqWSknz3q+TwdzihazNRKJriAvvv2slxaO0niZENrRI2NNPv5QDvF
I3sfFaXbeSwJG2sDldFPCpmOnNRRruUFYGhJrFLOMsr50e9/9KXKjF3KADrGYMDhGdvKFnN0XBY+
YpWzQKD1uCKPx+WogSUWSWouq1k57CrYO1ERkvdCjVh321eSHMj3vwG6mtWz+lbbCSJg9WnB2wGD
sVayrpMe1ACDLaLBVaxVVR2eDePCM4kHEhE6qX1b+dq1vBX/+y+mxijH15qJzoNgFIT9rSeawUR3
GrbXSwXlQsHQK+hJFtjpPTHs166uzFCJ0bvudLR208z17IizAEv4X3HLe6De7rpoubtXlOfUhkkq
6iUH2qP9ph4JS1lEbNeUMCeGpqi1PdEOupY+mnkXMbDsLxMRfLn4907KDVona8H2xgvlKm0B7jBE
CH4Na+Td+XQX0NAg3hn2hlp7eP/D9z7slpukrNkWqUKkd5LYMlh+PxPo5CAS0p2WWUbukxrVTrwJ
LLGS53Zso7cILLWXBfeoQhKueNLlezyoxqXD8pZMvzhnvqWxC6eq8Y0OJT2fh0t5KBuge1wxg6Jh
fMlZflqG0KFhRx+5GWmzgHDbAdTKGawGIklUBCxfaj00ktkfWpgqVbbv9pbkfQVCj9V7XrPCRCL/
A7SO1fqL/nHBVvKm2jln728OtDFSUldgQh6bKWtK0uJ+beS/7jIirnBR8mMidKo4Tx5/GSgnB39e
X/ws4RovIBGBDF0akhc0+VMUKVUFL8fI/IRu6YjueempQQvdlrxkv6CS3vzDUE6b3ErBaFe74RJk
ug2F7/cHFo2Fcp+XNlU6wYG+6Gv9McZ9yoWiYcz+zmn1tXoHCVuFsGTg+1VYgYw/+A/M9+G1N/JB
WBpDHmBgjYGb5RvLOLWgQIpQl1smfeONkoEcYbLgU3Bchf64gCw2PmR1irjUMYUXKG0eS+KJr1FT
CEqZwnoZZheov4NL87Zvnn6qLGXZVGvnUmoEn031QpB07zKP8B83GVwaBai+6OYi/QWo2bgqGZl4
0NF1o0iAdzJPOj5+hthe/Ig0rbFgpQjSmLvi3Empx1x3kLk7b2srhq4Q8rGHbs9w9y+ruvLljve1
LBOAWhfxSRln5ndpX3SupGR825lInWCbOx8amoAOhwR/+l8k9l77Kchkbnrrgk5Ah7K5qx2lf0b9
U6kvC9KL6XykGgAO66FoVcWYuRjmjrLgqzok8tvGaEDXFvusnVYPLx3swBbrHERiafr5v6LZgETn
ItSNyehclosjTFuNPsaOMIeMwufFGRSohiAW2ry545L0x9opMR5wb/pT5zo9lxUIm67AP0OB05Kn
fMhQyo6jDsEPBlk6GKUO8JDsGCablJzJdlZzP37nC5by1TZKTlciqj0BDHcDR+mCIY1cTaBDUoJN
U1pzqZcquprUirIDXQQ8dlcfUzG55pjaY4+O/Yr9QXXaU3QLSA2k4Mn9vUIO6dlTPkfj2ehVYUO7
8rSZkHan1BbZNxz1qNmQRQTCRvWREUoOOm+G+Shbaz+eKPjUOk7KXwFCoA5u+uPfH4hRZNT+oVv4
1Yll2ayyCKDvvn9d2eIsBiOxyWSMmb/MvJSqIDaDH3s162bEjwloobqmuOlfFpqiovmclsx3vp16
KgjQoOYQ6wT69SAUOWkGqintuxGhvYMOTF+jxXgUNbWAdvS4wPSJIuo3zZsey3IwPhvb168N5AT4
jPqiLAvkrFFBKyxpptKUAop9HE1FRWDFB/54U5G25yrPTU4K6g2mkjUfwyRJDl9TYFRHO5cWOuIP
OcQi9jkxNreRtdi2etsvoGUvMvsQTj09wPbfs1Q+8QiblLgvCL2KIEJB89w3EbYG+cx/KfTW0qeF
tpzFtYJT89SyVe/zBOIYYnKG8aDi2JMleOUXjoY5683jNSCh7YPqpMK84bVdjc7cDboQogwHxPdR
OCoxOzx3YNqildKrDjXOC4HNMZj2j/oENmWyMmCloTBSqddMGBbicPuzbFZYwt2Ed2/vhrtvm22x
XlO92jZ32fdrEG2rMUEuFBtSemSCZOrYDqg3gEK0Yl0AF4NYDO7NV6sjmTEGuXO8GAgbU+2OIpp3
yjio7JtnJcE/qisHTGN+gcrFKXp0iFE7EIVVjJXkCiAf5PGS6GIctpktd/d8/QKKZbxnfD+ebzmD
3+BhekwXhLXSQEM5/uuvzOYe6YNQcBzXwsr/oNCxT5JvjA+0V/4mgoJHLw4XcnEJLG6vpN3NCMRC
Q+G+zyNWw4POXSNQlEJnTW/u9X/HypZzshjeIxcgUHJOKJObFxxjo0hITaJTvofvv6LV82ezYFtY
1hEO/iTx7EiPX4Zy5c0K+SuSXXQxoyuDg4Jy/60WYYEwMAYmbj9fHcbhGsL78/S4HtdWyHy/PqN0
zJ0AC8MWAKfq8SPqWOtNq3v/7VC9juOAjO4L8wdJ9P1+hC+bcSgvjHFWV+o1t8jIhsL6IzJ6g7bh
zrc66sBPyr/xC+Sq5PkANx26haQqkerr4kWgRIv89XLT726xGU3SF6tQpi2pYcT9LN/ebYKf99g3
oWWqFUvLrMk++Ptj4GphtkgAkSknEUnzLJKUCRXtqKt+HOTuAC4qm5stoY8uQnzW5mA3AeefPkoC
v5otpcT0I6aKJG1Coh81SJCAg3PhmNLLLvfQt62/GYS6StHVmJZhWFPZ1ZFMkTLnWUIELAy0zH3/
cTFF+Hf/awnN+8cfJLt2NY3OYRDGci5NOf8VPswngx8+zOncONs0i27+Xr1zrFvhWdwlhCM+FNuF
ohKbmZXvmBYhXd+d4sgdNBOtwDBabLAqMZsARO5E27ShYNaJbH9pk/6sgkWx8Rlk5xqvp+wCVn/L
Mfzli5LaX+0uamgpyVd/wxw9YvP3ymhF8OP4MbzBdwfAPUaoLFpDND2fAqDCfjI1klm2qWEK0tGs
gKAPUiVOliSQZrvtCnoXaFZOavAcORTlCSC255wPbYyO9zT+c1CeOAfTd2qPf0iL3IVBrT12T2pL
pBZxwfHzrO7r34VvW3pFInMEWRAqYFo002xHHBnU/4fFL+AZfaDURDCtooYj+gydzTIhIYJTmlww
EppMuxSPcaYbRwnwh/T7p+AKhtKpaIoRGSat0GqTKEMMymEYyXAMA0vH9LNbvCN9r8r7Sgd3HRaK
0L6Rp81P2YOuaVg0j/CMTCl3qCdM2uO4u0VocDPJCT4fHBbls1lLvqJ7AJYfDESSuMSzGeCtT/M3
IOuTJsgGGhZxnxU8KmGYRuCKIQ9vQSQqnFdTPqCwGAQv0vPhI/ZH2wtMl2nDt0csMV0XKNFjX+CE
MyUMJEYGIGI7qKl5R79VP8/rpu0CFUDQiLyp/NluY3Xm/4eTbuQArIf55tnpeWoPMGtt0ecFHLiA
k6I0T3aem8peaq5NX3Dmgc2O5PGmQNi8Gc4iV2FikNOGaxy4qwBUP0Gc2hlFqr9Rte/3LJfernes
pj5sIX2rn/q1VzBJGXJt62OgQZFMjRNP342DLsZw8QAWk09AJHJWFzpBVlsVKD40Ad/NYcw1naBI
OeCHU9gf9V5zkmM5hKTYF6KbQZ0ol/HcG6AQnpey2wfAVef5IO8Q+Tj1xu2tKp1FrvN9Ib65BNiY
jrPqI9IPEgdhCeZbwZx13+hjG64OrflVTDOxpl8nKKt5nC4Zrj/ntxMb8OrJirpdxopSOaVG1TvH
oCauH1bJAwUPEhSP7J9+L6LJqcpbM7ZroNIJjBHQxkcLCxe8fibwH3YWWuasxnDa0WgyqxZrYkor
9Av85wmXQURY7spSpJ7lNNJQA2CAuxuv3YcMsfUShEqRZBz5+xIBIj41FQ3Qh94w/Jb2xG5b3oCc
LN0CBlAbjKpcdNQsIiSehRPLW/9AILdqYiSXBcylbPO3g3SB/3HPQiHfIQSHx9C4os2bzkAm1x2v
pygolh+hKSN9VuGPhEEZYY1YcGqBMejvh9D7DKygsM39Fsa8sP2qbwDTNt1TqZqk3t5XC6yuLntg
tYPXRzX1nwUW6BxpQSlqrxVn0J01DF/CB1tq5w4KCfotNroVBMqlXTbgJkO7vSrbSKTVc+hIjNEl
vRMYIsC1CFPJeKy4NX/Y5i3DaXW+OozT2fiSDQgAvipoAHsybbQ0iOxwREnEtCjY7TO/Cd+YddN0
LrOBgeOOAJ3koGMd0GvCn2l/ZCUQxgHlkCBOgPRLblOTzx+GL/ggNEH6AdeOTElznZ+51Wl+NHdv
eJzKVKPD2TP5RISLeSXpIEW2/HjjtR9htUVswsd4epplgaN19psXDHq0lKi4+27pwuynqwU+BsR7
mpqEFWYHf1jdZ2OAxqoXb/XSxl/KpsVFOJGUCHNg33TjZBYS0OUPbo0HVm/GPhTGRzsw6LbzHTbQ
3ZzRH1rqi041+Fmi15GOZ5/PfvrBDLLFPgNOTQZunb9banBkfq/17fC5mOmKEr0j1dQi8vhwmo1a
N4n5lh47h9vUzqkWEJqj8dzM8731H+SM8isCadTi4kslzLI3ZjuJwHGp8mFf8X2BEvuUe3YLDfwb
54OzVUldETUyhtCLbYTjFZAcWgjbU0rF7mmaPgfaPkWG4i3ZbTnnGuXO5ZpeK+KjDhfEjAVpECnS
Oszp04DnZ9Qdu5CwjKfFv3v+ObatgibYgc5h57ld7O1/DXcguVyfQYn8BiwXkzuTBZlvwYg4MFex
ZjEk9dfRoe8UTc6+4z9KpbHKeWQUBp+UzBSY2lBP2cmldDJ5EWcb5IVJLgzDW/cq4G+S0si5z/cE
XUXW3WxdxKGksOymuvwavWZXcPjxbrwR6Pofl5mpDZfyxPGtKoa9B6zGAuEpZfP71YfjiQbhMleJ
f3CJ8sWFs/+RClVQ6zvpNT4vjT+6QMr9isQrf5IOzmzp23YHbUIgiVO0NPdo26pcxoPy9/A/JXSB
Tyh/4z8LVXM28rs7SKtMpoMOAHSrUK4PGPrVu1tP3pDWn/oX8rT4y61uJxzyjStT7HsSeKYxkah9
Dp9T09etMPAlLu6afJBVxzcgeFI3m513tQFWjuTj3c7vz06E0iGqOXpVLHLxm0EnYzQNMWlWSiOO
1dd3ZXMkEPADpB+XCuMuTm4tVGnJjHPXclzLIqcuKZ3lr11F3qsc9sOG8zeLmCHNJiZ3cd/oph9N
VNmq0JhDRppLUDxTdRoBDWKdKmhm/W70IHa1gwebRZZHtey4rYOshCmI8pzru5+qyWnVPjzS6djh
JPfW8MIpc889PQjhwVQ6L2Ew7Zh3YxIhsB2e/RWpOaSCIKHT3DBGK+/LXFL67if/DbHOwSrs8bqi
D7H1s8bATOAdEC9oTKG7co/0R6TjHTkaUgts6iT5MQVOcBOVAV7+b8p4uHlpUU4rWJJWP5j8sKiB
K8RqkvcMrIm20ul8R0/yCN7yBQLDhBCjkgchPA0f7AIgTMfKwrwMB1Vs1o8Y72AXFq5ctV9WNO9L
YbHVd6bYmTOwQXmFwNpGzN5fYleJ7ouUHJRlSpcPryaQdpf6u6wDgT9jsmu7Yo6fdLl25saZK4FF
BqOJWhX8ZsSEwtBb0QfduNmjPHCqo1xq3EErgijt8WYRj3AjClXpgO4g7e+mCyb/FOgqP3KDy6E3
DlqsdBlfyjUgigJRFSBf1pXh3LC9AIQgel0wafgVdSH/rNNFO0wsBLiOEioHne1cANCr+qbhbz4i
hUn56vHl4vIGvrrAM0gAzdNY/PXedi6ZtQCJqjjrHAmSAPs5aHW+u4pDacmYmgb7/AiIcGKdfDSR
wx8PkNX9paVrl/LMX36Owi+BtIyg1AMQsRBdXfeC5UHYDJO3mBF6BqXTqvNz2wFZtkC3ym+DKjBx
mGY9OBaWpsoc//HB31W8eKQcMvZg/4VJ2Dx2FZVnDja+pooZEqTU7tTgMxIcLLaO4zxD5fqK86In
Hx2+U0iT91pj+GKCaUIUumOhaDvpXME8B9ZFFpI5eerslo+6HPEnyI8OqfxxW4UGj219Yv2owlHg
34bN1Wq0+3PDiLos83HGWYMiJNAUhtRrdlVnKVdxoowO7POfh5w9hdSkoP/gfBf2prwMuSHONMqO
ljrbwhQjU9hqUndoWOzmdHImpScxbPJFGUWJRBRIYqoXvlVZp66DsmG3U9g5w3gMGGvheOGhpzQy
7rEZw9rbQGrq8I7ClJMWluMgi9etCyj10KE3Xs5BRth1zhcJLep49fNfSAhZHFVessW1DR65Nwll
VrWXJijjeCA2HaqcgRzHlgM0dV4IwcUbiMIHKBBjv1T7GNpFR92IClYj0M/bR+sIz59df1+Cedua
D6fmk27aKl+VDI7qJcms8CWW4dn6kQEJNTW/oLgmZtzYpeIx71rxOk2fGmrIJO/T9po7g1Etu+AA
S1i9PJCLXqiHacDzbYrW8VzmNhiyvCAeui8Ox5t0/RFjjg3Lnwc2AM/2IIUjRDjHtEfAnyjMbNKY
aZeU53vKgH9pZnGmbgZi4RpeOZxFEsTCLj1pABAClkvg8+zD9OwTTiwW6TgZ+LDfZUJl7SYf8p72
niSNFSU8BFknYCF/chb1VNKyi97MikYUtlp/TzA82uvfICCKrQpjShesyMxFbpwa9odIQoSNaGtx
LokN/sH4vcuWUEnVJEw2wDli8dWuXG8MGVbuR5bL4bFL53VtL63kGoB6O+t6JxuyIFKf3Ef/uBW9
+ec8uV+s8qs37GjZ6d/a5+8VVC9Dl6H/DJ6eXzGdSf8Uy3YSSJIQeoGYyG44VzVHl1MOSzbU4R/4
G866/gfMdymgyWG4BnC70KcHcB5XSCqGRuWiFITOrUW/L9m4sQSBeIVs+XHBNo7rEZGN4NGwlZem
38CXRApiGWBEdSXEqA2nhEuZMHpsUqUl3JpQBjIuzdGWaTOsALnQuYFsIhflQM2qvRLzu/aAjNW/
GQs/H+7d661eSvqo1+Y4h2aBQbm/ROua5GIAFnEEJOELmk6RGvLMc2SuKv34FYkDhCGgqaANty7R
chZ4PSKxx+Gn+/7N5Z1B6ljYwKRBrtYjeERx9mToagHWicWEdkPSd7cU4NcryfnJ+Uibx944CNFy
i/72dO/cogAaKjTSZb2Qbh07CxJEP/A9T97OMtxMK7+79UI/agYupzN3691+PDeFGgLe78U1WFmz
P8vVJ5Evf79FOEjAjq+ypWWvwkiVL1m4ncMTrbQlTfGgpHqVJNQrQnVVww99AcjCFUWa+bjvcEST
lvsxthT16ndPQlCOUpXD7L4I46TU/MwkcUNeGXrV7wYeXHI3P3/LuWetY3Y7duNICnAvZ7apBtfs
SqH5BUEdKrlcyPgBIUA39AZNo97XYAqgPA/7ogcYDWKhGPcIVM8vS8yehECf+TT5ua5Kxa0Cx0n5
nk4MQmNhl/r1d/VC4RXdRgxwDFvZ0+xzkSfCHqQXKyRkTvgNNm3Ce82s9jGAQ8RLGhvrWJcVS671
PkbSKwpM6hjfUWx8qbjgcexN9gEN6CrgJHbKavLodP09XO1ciVqOCF/OnCMoy4AckWFDyrhD3Tel
lYwl4pREN+AmRBoHHOONXaFu/uK1u+A9wCLk3D5r1J9Nt80KsZq40Hqm/11vhgFsUzW/q2GIF6Sn
/CaYgaPxOmucqLkF2br6OcD5a6ELdgodhD/rDbYXbqw/W5wwm3zRkbt0fGHlivASVTefPWTRyiYw
VGjvPi//dfD1Kx+zdt65nPH2X7VTA9j5ysbhodRPUMvRG3sgmtx9ftSnKjxBglGclkCnGLTh2nRj
TXo2XuRCR97k48iexpkNDNhEC7Of7stoYGVPslYVgHn/ZjgQu/jOLmMSmaIT9bzN3+tjoXqz8U83
vrqGUyNbXMdhCcq/BO1CJ6SgNFVCBZju5I7AYgI4UBZTqqDixUKsO3EGoCCDS7Gs/lwPkFP/hK8x
RZR1YGh6LbOWA8V2esaXu5CWC3+19f2gepnGXuCY+V8kc+Kk3zXxL7+fv4eBRHZgV2h4eBjeJtcX
joV1Z8Gg+wXQaqY92muRSfbH7UHLF8Ntim2J9K8XTlJy/EwhiGIL7VcgwNgcqNvmfpb1M+03hm+8
hyp76+YV4dZelxhH+/6vDgl+4nXGIYqU8wa5mZfYYbRafDin6ih9J4kgJK8wM5m0WaBY7Vl9RBHx
C4Egxk+U7nai2VjPyrN9geHe+QVu33+vapZMcQt427L7Wkrin4YMGe6ZQnd4XbIVxlS6b+ccykHo
f6tSlBuMOP7nPwM3Hu/O/3r1SO2FddJk3g3BtzjJe0M1xzF2FGPkLlocJF0XznUImXFT90dNk8T6
65f4GVc2Ad0/QQJoYmr9uatqJAYqlzRl8gV+cyfW0Lkhm0FJTtuXSYEDBVU+wh9U9IjKbi6TWvPk
V1rlVjoWCcK8yPoM6awPxO0JpNDtq8GYqVI0D0jRtU7hMqV0EAbQVjI2Ictj9/VBHdgMnH39k1YB
taxjvVI1QBgs5k0WNOtk6c7ll0InF0g94xTAWv9R7ijL0R4xYPALBkcjKAjDkhw7dRIgQLlBpzvR
IZlw8oaUaQPnO9MF8ZSw6ke0yB6IlVc3lD816JB6AVg9ngj2mafHU8MxPDXehmnotELRCZwUALdc
BbK+AW/Q/oOSl1HH7Lliyvg/jJzUB6vlS7gShD23bxitkvde+AEC/DpeDvqLRLbJovolWWboJcOw
REfH7QVtrrz/OoYCbmC8xhyL/CYxzBXCcSjdmJwDQAxLEU4mCNPKz6SLgkU3KMzgGxI69C58jBxz
DZcqCHP6rke9r7fdZub9B/q0B8s5xTkjdP5/HQG9/gWmXF5KUWk5BEuHG2yLybcN+QTggkPX4E4A
wY9EYqpLr4iloIbRsfuNNms4mDOPzWbFXsxtO+xGbOgxFdkJV2i+rr6TDiuIJ0pZ0tHKQ9Zb4MB1
RzbRztRFT166BdcsjoeYu4wnZTs/GCmCFdiKuT8n0Yxso7VYFoirQhsEt8iwalT/FwbYfkCGI+fc
434LL8zOw8oSYYs7BuXFXg7GUWD1ejMi4jrbwQx5zd2KwHa8mooG79ZPy9UUDvUUCE74sPPWGrcF
bufFBVskkqk7na12MDqiEnbbvxuhm9mOM5gDsq6cChsyF6VaiNreyZo+1HvoQRUXBtO30S0QSjEh
1FSTap55bgdpc7TXTs8Q4pgfYm/cu11jQUOZ1q94Ke123YwjKCnYTm2wAMo9QzkJMHr4YFb9U14W
r9gBWcWDi6C2kK/W1lRF5NF/aB2MJzYc+GqBd4Sc2puwNwv+sE1ahC/Ny0bKSePKC23z9kgW1DUP
MYp+OFOUpg3OgWHDl4zRaKRiXaJsPIjuLQITO9yCWqJ44EIw1l6uo04TRQIq5puHpALy9AZ/BQ2k
F0MKzY1ZjKFeqHRacCttdoTRZZxfsSdUBwsnMKqOJ2xI9nN7b+Lr6Vu3OANTPNHWzwM2z8AUqszG
zXpF/lxBZKY2vpSQ4M066LTEHnn4FhhT28mNL7N/cA/jmp/MV1ig0du+Bf7/HulKibl56p8Rj8Yk
eRqvoYKmGvfuV4pgY3X9xdqMovzk96Ushlt7vQVi6mj/EaETIjqWQ/Uqn0sAUyBQ9q0S5Uk0suwl
rooshtW3nv+JTJ62YuwSvieFHQ8rj7sfrwkDLZkRk/pY6+42bAyflKr3bXDJStQws3k4H1jzAG2a
ayMudjYLX+oF88mgecaF7xN3jFcoP49Gpd8/4GO21lvp+2jONXI2Z66pNENCbXe78ORmBTxzzjIG
/vqNnImNYGW+u/eeYUFPWUIiha9Qvx55unPJ2149TGgaeNnZq9zmy+sYkF3fhiuFM/qDJKcHatQO
ARYd/YgxLhLN2tTiOhYIIH+7QWmOPIcedDl/7yJ6muqpIr9TMtBeltYWW4iv9evhzZzQZdCTuHc5
df3whWxnvaHJfH8eMac6vbfQsmOPkEhhPcAxRFVxijsFFQkAF0TwMBUasTHzEVz8jQRCf2OSpCuj
jbXfUNt+ZbPPR/bjHNBl5fhXiOU5Cd0x740XHF9YUvCiY/vSZ+yJTt/biyRxHRtC+EYw40KR0dTH
fqYlvCr8Jj4xKhw9omE6uMitKG79itILGeM1ATlniTOL+pkV0cJ0txcfu7TTYohugwLG1klIyIp4
XI71tSV+hZ4yRy3nll/pOVZTZMKt6hlPXfYYP6sR8zI2duY1c3bSTl4ggheAYKRS7cRPdCKwia/i
yU0EML6BumIKFWYzkaEEMQtRlPRB6aX/yEItLPsFR8Nd9vYwozGHleymDbPsMBczbyFqsg2e5VmT
7L+fQzJ4k6N5cuMjA+qodzji5bX9l8ZIN3ohuBkBy7MmSWaIw0K1CAS1rrGqgs571mwqUCJj30de
r58ucPAB7je/D3dgvwE8DHQZmFQn7g0G8A8ppAdu1rKYOfNp7cLrR4P5siX9dTqu0+FsvWHU6mj5
3eudrGY28B6Qpcnz8XYR3TWUoi0VIvCDpWT8xrkj85l/XS2VJV4fTev/ReZ4ywq76oWJmFPgJ/z2
6eiGNKk2QybvYdLfpoAhcmrcm6P3iaH2eZF0lU507Pm9WHvtcA82cGiV6Prf+6QsKbrlJ3ZoK3a0
v8cpSgrMdxTwPVDJso4pkmEwlJMhr1HBg9cOaGgQyay45xIVf8q56L80w0KfQnodNvmQou63Ic4b
EzG4+ZHxqTAJkNUKy4YQeu5wB6m255FMLAX/Q16Bl6WsZ9PaYTgBCswHPdkNAk09eVaJvZvHaWdo
mPWrC5XXi6+IihmM2ltxWLT80Nwy/RG5YQDShFHU2GGB5+FQEglhDu15v6ILFcNbYjlIa5pz6zVa
RNH8ZlFBmVaxxJn0r9CcBea2vN7eRlJ4XR12eSVIQ/1uEXs/ecKAKqSzhPV84Md/4CTErMfUdyG8
tskcFMDIRQgKIlSimlidmh57k5DpGopBDMWihsDn8LNECyKJMpT6Lu+dW2UdEkwkoMLq5U+rel4i
S+MzC1+Or3p8BZk/sG1KRdqBby6Mky6R63E2ts/cFXqebAl/wegYgsrgTr/Ts/twM3qOHB3fGQqC
HI2arrKDG67e0KclVMYxGJvLw2DMPh6WPm1EIpNbjiO8AfwfxRabiybewcPv149j8WBkFPbPh9QD
oBcWVAi3PflTa7wL0koAlLtF7Y4gBTJSV4DmVxtBESKDgGr7KOIb9hTs7kIRVSg7aawuZ1Jpyy0B
FQeYRAMu1Ape392KqtAOZeyWjoSjuWSLs8oyR2NHp/RMDI0ji4BxnDHW2cN3W+ftvQC2t3mofIZW
c9vwDlS4ucfMbL5YAbuLY9ikRSb7A+EtTgoKc4emdkbY8tgGCL7TnCp2E74DBxTjOBCA7Vsi2L/D
gfojQr7P6ceGVbd7V6A6wragOw+SvqChdlKhD2eo1rG78wDc04Lamh7I5RtTDxfraAU8uzgXWAek
cyAV44/0od5bh3cJHkknCNeVrxLyTZ3VqqOUMV7lGYRM9GkfeT38iXiJQ6W7s7jHMeZpacWuqlvb
lhf+7ftclVOd2S6t5W+8koGKjoyJxhvP2h/Ua7vQA8SrGRdq1GVye5/ibnK5OHge4G+i5Q4Z3k1r
ebSjySFUHessWfqh68TTtV95eEoJeocdCcH9dtQ8gfhlW3gwpdGfuvvPrnvTp1n6NKYqEQKdM4ve
qDtfsk1sUY54u5iS1QdmYVI+gzuXaq39en8YqMzO1OqRN6BvZE7RQB/mtTdCJ4qavQLDhHVmHq5p
vKXbQWnAFRbIbMe3KBxQJ+oyTxWWv2DqKoLkDyVnokBLikPJUc/X4+wLpQFFnZ58Q1ixCvnQoyoC
cX0IS0xyrhWJA5/ezNUe/Oq6s+Qe0ig+RB/hro4s+iNhy63gwbUMfFQhEQHpokM/xxXd4zKiemOa
gSc/VtpxAaq10Sg/69V7mOSVXW2Tv8PWd1uKBSjD1eVnoT4ttY00lZX7G6v4oppv0I8xaF/d2UvV
htuCJ5PDZ+AgqDGGUnB5YByz/aj85xAn6xb+sf1GyhImS3VY6aYkU/jSM7chyuoMmKO1Q5Qdui8Q
XWhnBebVyNFQBWUZlriuDKUWcZRoA6uE2BKoAnm1PABilMfT/j/kdLR3o6PzwjRcio2X+i7ppp7L
YHFAyg1IFpg07shcKoZxhULFosi9S2Jqro4i8cbq009A/pGuNBAgsT3W+JW/bsCQl4AHF8cKt9hC
fxZbb//JDGiq2w8ZgvepYCPE3q54IyXA7fasVCPaw6+6ukfSg81lZiKlRUqcT6SmLP8pewNeV8hx
U6FEcMzTYcE4E1XCMiukUrY4qi5+BIZoSqYLI70t5Sjw9+iPRXHnz1C/mFdOxOHkeL64XxEhx1AU
mD/W5h2jAifIyDflQFkg+dm1hHB1lh9ySpHciCpHVeiPcVncLvfqe7hLCjRVazCYq2I9op6w/gBw
4wS/kP1NQhjXiM7ziGoxja/P54cPtE52SOoZCuaf9MGaSdcwS9Q2g1bGkaiZ7XgZhZjI3vEnuD6f
Wbie+hZ6xCSOHKuOdn8IuqBWXCkErmnOjG7IEnHQ0y1w4lDuCJ5Ci7pW4tAA38q+E9Giq3rATx1y
wIG4rEou1uf1Ig0wGi6Y1xzNKgC9iUSS6ds7xTV62PzGoXcHmMihXzSkmb+6nOpGk5AJyh3plOHT
iHx/AkRnqs2l8vftPP2QzmgmUM2X/hzsNgwkURYD/9MMfdcdO74I6ndrwYGSbIG80/reXDFq+qUn
SP1hZfaKAu+83CViKUo2fGvwEIiTHuyAYLJqIDYaloI9RjrTyS+bq8vz+r/NrLBOoNu478J8uWoa
fYnUV1MdEjsJORwit42JRSMOmewNlzGsgpDWdSzfUeniUp1l3cujIpU1iL7R6j7uC3t4h0UqDlp6
gEylfZguqPBUJcUgT8D7KL3askZ4i3A23oKWO2pIrkc8gF1cV6w+FkdX7gOUUH4uMcy//rTUw/DX
66UBG3gYHzVussjGpoxVu7VDkhkp1yYsiL0e66iWDXI4YVR8qIsGuTxvuBvS83hhNC3FVZKZnFaV
WQbodSKjcg17uwIsgpOmOZnJ/WYqIj6H2mc7CnV357yHqcU+OFqj7iasXKr0ikv6vo1lVnVLTrb6
1qnMJqsqTXN8QXCqkWT9C+QhW8HoRV0odm3XvgtxnrY62RNRGxbC3oDco1bBkRVJOC8L6Bh6UbHf
0r0j9jw9/wr2qCu38ZEuL3IkJOACuredV0LP2qo7s9iG0hgj6rr0F/hsIVzgIUCUE1GBHH+8NL4a
eBAzK1+rMjQjeWlfiW+LvImNcqH51Nfkyoqf1gT+pdppl1gQwZ409S/PAcJZOQ4+EYSEMjFrESN4
9DXwDK1tfOCE8pb6xRGrRKFuGWs/PnglLON83yNiKzgUTIZ6NwSZsasIEqPehbnBtHAOUCPjizdR
09xoH9/pWFUZwT7/vW5wrTsaLaEk5s7+0Fvy484YFjGbtHp5Rky6TNhv3ZJJ20E8aCMYOxGSj6Ao
OE0P98blP/5zH6awUQtMo++xCuaeSx0/OoEAjFuCoxGiMRN2YnU/CnTvbvtAbTi6Nxktpy/bQOU/
p5dPFV38APlkL8wARDdfqOYL0i01yOXjAHI/ZuVw4bmO0YNO0LLSYV2g+lyDwv0/5wOFngbE399d
Tpm52dntMskZUy7lL5GHGuoqE7+FQA44uybQRB0qaGAwO2etMmf8bJPl2n26m0O+xzlsuno3F5ND
dnCDi5NZnN8U3sMBEYIDFDoemulY+x0ndktVJ7LaegIeE5IjthAN48MXxoEsafn8ErSe01GvtnnA
LyJ26NRnck9YZYeNcSuMEiL6GGV/ZE++RqZ3F4XWDtkElu0ZnJzBzHFChisUYu/U+XAOX/ncj9K1
qxN1fw9qvCTRplPJFF3x+a1tVqImh6IG1fJZXN8lUPvU3Z1f3co0Fjj/jhZahNrDoVzu0CUs8GRx
GjO+yDPq+6LlVUz+SupToJ/LPiiTH47AI/HQQogIDTnFrgcnUFM0YtLzkSBaKauDua4lUYSngd3t
p0ndLuDOnZ5yuvekypgG5cMtU6nGy1thZbhPRyzhnIEAB8hH84AJtXU/TQNRxD/DIXb43tkT31PV
PHrIUxnXCNIuCEqxWXQSNFYJBYWL5fiwqwg91U1je3k4JxBvA6Xggr82aoofVqSQH24PB1+f8O2y
QzJFGz7JedysgWdeIoftLhsah/CgYGwndOl9KI4yOHaaY9xqeNQUZBx6h4pDdAeXm1ZmYXyp0Ymn
B0KiiZMuRrzh2Y1lONWkt++ce30LT2ZzGMZcd4o2JJyiY93wo1QaUSZO2LqunJFx/xff6TnIbVCi
67HQOfpzJ3yX9RHAWqt+lWTOe1/QGW1949YG+RSyoMF0l6WhDp65o8WiTksIt1hzumiEW0ClXS53
WnGk3Vups4RR8Zq0j6VY+jHCLDoJyK8+kd8VxRrPRMzTqKGEpA+gM9r2RdhdZlUUUVAEvWH8MAqN
3PMthO4uiWo8AEYDrnF4brXz0qsGUTlJVqjjipiWGz7Pq5YCGv551Pm9AchJPiHGeETvRstjvn1p
R7tdBEchBU6aL0/mpMnSJz94hJqr+iR/2FdcEI20dnGgLR4fiiukrNfq4iu1nc4E5DQ6GzTluin2
H7ADFgKI4ZIL5mKRzFCLmhuVXhigvNK63h3v6/Z9uWq9Oydqf3tF2oMhYyYAVRRRSGEvigILkXcF
MtD0GMaerbonlWLnx/n2CjWA9jIuAMcx2xpqZ33C4/OpIVzV/KeLNhQHAOvSi1VCoaWwXCuJKcRN
wz8x+zua/eynNXdRxSWb32FCD22EEEisteovCioiQoxKcmqg0gHO+4jrexZHc9MJCGkZNLoR7Ujg
KojEWidJUFc+szPP29jQ4Vn4UTJewAbS0EkhoXP8P0gtHtik3AsEPV67qe+dVo++N6rXZchmPE3T
7tEgwwcEYE5Vo7wWWsgrG+OnyWKlPwue/LI+2Z2ZEku0csThyH4/Ch3nx1QaLeIWhknh5lO9dc7c
dFZ2Q4jxrdz7fq1dnmV5cqPHfU1ZDZXssNOUKf5joe1DVmlitQpo3gHbgykJYP8xWZ5rqBucArMS
VmrzBHFdpCyy8TyZrcTaF2gcSohSr8wqc1UMz/VL4af3R5L+DV0ieBeSBd9fjqW7soKWseoFFx9H
AQ7+drUEWDlE5IwJpPDPzqmYlWPOLxp+AA8c24wc9FYvfgzryQ7bYjKMnIp4zDAhoWKe7aFXUSNj
5gZWn5gEVLXegOYD+D90paFwD5MII8l+Dju0kcCZ6uYu5diFAseNpyZxJJ3/92q0z8NiXj3Y5ujA
iciFLp5e3O1z5kZ0XZGGjJ3oN9R9jwbbHHXZT1Vh1uYrsiZ4b8ZSlenLvc+DCLhy2fKqv3Dcpd7Z
MUNJ/Sii2d35qoTHQUEFLU8tMMhv8geHCP2U8fceOSCXgXXnXnfmxuUojwyD7T1b6goqUCge0Otm
3cjQ8NW3B4n94/U+KjYrxkHcCfPQf07l4rZ4rTSzorMDncgvXK72HjRrNe/h4MzOt0KoXyLEfOgO
JwsqxsI4RvfOLRRQKlst/5BDQyGdnuJ9CFXp8IW2YkzHsyqxd3dboVJOGGwNXK/wnBOlXmlvHFuc
TC8JL87+Cl/16CVWchPhTaFK7kXTY/5aMRZc1VUzRIHaXD3qYUEcSyN1TF5ZDfEyoKaTr0l8jLdq
oVOJ8k2x9HWKD104DUNDLGDLId68A4Yq1NXhlB+IwH6/yrh21XIVxWaH4seUUlloZ5gWzrB22LZ8
boBPDrDjcipnbEjacr4XgAOAeRl0+lEiV5kjPZSJ6jwHss6D25FJQYwnt9f7D8q/9EO6s1jxCZHH
+WW4F0eWond1EBP/J3NTAXf+yZNsN53/VWF/RHESnrobqm03gLbtiuxi8TgnAQsHbjNpAFod5LTu
8ESbwMfSbuCPoDp/RZlWWv61UK4ZJvKuByVJFce/WS2cWkHm3LiG6bxP0efV2qewi34R0Dib1nJP
9Jm6VLtHC4dcbURwoCfBEfyd3bb4YypEYH76Nt+5Eiz84Rsv9RZjmGFoYVF5/h6lS9ze6q95HILP
tBo2gFzErM+Ad/vIqTX8+ppBBlrz8dQhQQ/wri2yeMnlqYyBBMagwCjukBsk7onlRKntuJdy/gdd
aFlbn5eYFLCC57cvTj0ixSCMFXw4QgbUWdywysNRT0D3siDYXU2wYRLILLPuUkd1bPqtP/z32LMC
A9uo1U8acOuMA5zIFPDQODtT2RSglgkruIaqpzAVQ5FHRIm3j/4zGtl74l4sfYA84aSmWFZl1AuU
ZdrHdrRsQdaJhpH+GKKVykojLQ2FPfmqmdbPdHqPjZoBn5enGvz5fAZ5Bfm184Q8AaWCMShjUxu+
i7rEYsiCMFLJvXr3f4UlKWYo1gEPFAfyZ9jIhYlM1A0w46K6f3ynoYaaCy3ofQsqv7IvcUy+Nb9u
XO5JpGWcuN3QNKZzg6zLU11SuWYIGo6hLnuqp9xFq4gQfO7Bien5s5U7zU3feEJwemn8JskWMSk6
9aim+ctvkaEUVi14n1CyzkS3KWYGmm/XkzDEh90dkFLIJ512KH8ok2RtWvDcf9U7m2cM4mA2MNh8
hX7lUvBLcmj2GHg8WMg9gJLknH1vp9DPZ7TrwovcK31Za4RQ74Zh92Uey8BhtAUadVkIvx80ZtZX
7wQSUWSMCvsIMdNPYM1BVvANj5gc1BzFlv/LLCl0bCJV8NJTUGJr+wWwy7+o1ECSGsG0iapxGpyx
Gvu60hiqNFakRY3GmcgNA+wvF/D3+LLVv7kCAC4PIVhlh4nU+JiLEz3wag25G9jEkK9JESdNNa1U
la1z37OCvgrYM5LUO5hUimdM2+dJ2bPN6j8ClA+GyN3nf76P5zK9PXquDzhxde+9V9W0jdkDxVL8
QTzLOfdRdfZibq/5pfyoWUnEM2rsOEiHA7S4N8VC+qW6mpaGfu64cbL63S7yq5hi+XYnhQ6IMm3k
fDR9h7LwdYHisobabiX2Nrdt3uRvcRd09HHaHhNtvr2lsUPjjYcPQW4jVgs//k0rJdoey8H04/X/
nDwSlzFFvA6iUITX2WgMgygcRmrG+qzk2DvFiERxQqXs55RiYRwy8dJa26XUWQY2DkiECVQgAChS
Aw6RSnESPmApxzVXLopSRbRbUy5A3itX/PmPDd0XoMsFCGWdG7P86JcJX86EHUq2Gj8tcDxSJDwm
Rl7MF3ETXbWfhCYPPTDGlmHqQRcQQBUzsXkCMEV+HxafhBR1sVpCj12wQDXrORxewXFUtDHWgtCg
zedDoeR6MA1Yr6LSj/QuEONHkqXZ524lUAQX+lgLiRJsEutvqX01ks948yNUufgW5U4LLTgQuC3b
s4YLJwWI3skNC5bTogfKvaBZ2wYDxsXY3XkNqXa9gN7fsjl39YWsomWrbXFTAj7dcpNwJczyCssx
H6wyZWnNeXgZmMA2lh/Pz1WvC5ARdM9EEDVeCFwo9ztS8tlkqGRCX6IPfAuLO/zTXvjhMYR4yazG
4krP/qz2wm3DhzpK5vY/qFH8wwNyr269igAMjiM/bLVN+ZjxmY2wGCUkFtdgsIy4nj/gUWgrSQjt
Pe2clMgqzq7ShYtYb9TPh8rOMRslao7NpJdsdp3sn/5JztUdl3N3ML03O2FZbgwTB4v6e/esDHnS
QXx3Q//Lnmy2hfWLMhtDhIAThxqnLNnY/NiykHgej7/VorIkvsaDXT1E1ARq0kTeiAtAZRM38JUF
Wg/0sMjPPrqWZKr2ffBmPYka6LLa/0nLJMks1YtFivdbqikQYoffu2GpqvjgibUdEjJ4zxRdTu4B
7F4LQDdSo0k+tb9czbaheOQBWREUJuWwfjTjVY/QrgNlOuJM0uxUxzfrtGw2WOPRLSJb6HJJ4+Es
7zS2KmYP6/AkkokGV6Mn0j3ekkaWaLqYx/nTBDnieoD4N259jy4lKqsUk83mVeB/bWiD+7hMcq0m
RpZ747lM2pe9zfjLVvph2ggs7Lcv24uFSGleSf9XZSWeiRSNA3nl5xqmjSo+G1P+oUZOeR/j13M3
oaLOWQMHshkihUuDHq5vhZMBom62Z2dKCCUFYlipCET2p5B9UBZGq3qP1vqu7n6ryIznCIXYDtih
lz0IB9E8g0S0+A3VYWlbd4BHxbQxKWrwcN4aVGzA7bypQTAM2+yLLP89/gX95SjYqM3/PbWNhMgD
Rt/eWlrW1t4oJXiXrrf5otuDne4LRArU63z4OCqHA9VKAgnc0eOlLSl7CbrrArverrHYUG9v+W1V
+1bvsPQcevn7BRn+l6X72vf7J2caNoiK9sLHiwtd4vvPA4Ns2+4l5Av4wyuMCVwKTP6qDVVmigGm
n6S6es4M+g1kmwfJPUjkktoE6/21HBRX2gaKwpcW3ePTQhHF7dkjudquSRZc+PY2+auDvSBq/Ig0
BezLe0i99fhFI0YfEY24UpoEfQfNoPYj9kafm68cMSQp2ZSgfEXECz22OPXJP5hKKlGf6bn39ZNs
ryAMvnIA1NPrwfWWAFNjKLAGSWFVoRBJVo5IGqoBJrk4axqxNQuA7qoG5kAh6b1sP5RbX9HUW1y4
fZME8J12QQKogTCEimsmNEB1DQ9WjQeTsTy3eswGKTm9Hg5lz/0HBHDgTRKS+mwjdR0ao6AOW0U8
5/6L1TOgNZT/UWvWgV4RzXc+fhSF3JProzgo/w9l4ltFr3rSYKYXlNForU6Yn/HJylrdUw0agGDr
J3WPOArRAtjgmsrpFvS9zFGQRKuH7HsDBabW7Y+XZHpmM75A0J06UxKaDcpfMzHrXEbir9XSf3Dx
eHmZZVO9UQkhSiHQnU+ZrNR3Dh/mc/dginPSK3DWimXelMEE5U4XCv/6Vt0TNd0I5noL7GKVqAW3
yne8M40zT+n2LlAHBxtxURwFpK7BD/PAYawH2QnWG9vf2F6mMYwVeTG/oSGxJqOJw5wTA/oYnjkH
HGmnFCAYO8mibZ2/zlIzouaKf0jkQMGr6lEWdyDgVPT0Hrgyqg2auVeA4Ap0T1CRcbX/WU5/XrKC
XplYMJ+WFrQwRG/Wthk3Q03ZXV/c/mfQvx4Y9FedizemDGLHp713b7I+N/VEyxjCiScJLaxeYUUF
onsGbIAj0xGyGG2xUSYiwDRxDrCZLbYbwqKVOo8sEpKcBCpPWRWb8dh9X7mtbvMb+cdqWthNmdt+
lWSPQnxoL3QYN1EUf9pVwG36umHRRHfAG/E//K80Kgfh1kYCLPNTVaFoCDN0T4vSRnxM5BWdzRxf
OOhuI8iDmCSMB25Tlfj3VQdxmZlxvCCiKDUIlPhbE6mYuCNSHVSeCyVBMWq2CrJo9BRDa4EKl8bm
l2QDPQ+yVBJJ6P0WJARFrige08QV3oWwPmHhALOWGW5USiecTj05SP1o0B98veyLJwfpna45vQy/
d+mKHrLCJVGPumRLIgUsGKyG/W1ldkv4iVlT8ECoX6HQtDQ5kqwq/mJ3cSB6kScSvdBkDsHOTeaV
rL82iZTP3Ot5oZrvUoH9uKMC0KN1uPAq9xjBt64vzOePE+vBS7BPL0+2cR15B7kgKIfACglVHiba
gVZE/PkPgLHC713wOF5UKVoVDTGifsDp0pqL1tMSgMrOly3gCfGOjhsy+DCpvILAYLuc3FMuMtDo
m6ZeJ37Dy94S4G83C4oNidPWxfLeisoXjbC+mdUoD/97AfdWNMy/pBFhjskAjxrAtNuYGGqXzQX+
SjeRb2z8WbYk94SUtlDt6B8MlrgidEgqKKFvOZkHnj5XaNgpmemlEuHh53GqaFMq9jCFixlzKVrX
SZuSfl9ZxkZ/TFlaFMvWq2+bWdgZ6HRJN02vkPCZ8bn0iWys+9wm7fnQjz395l1aZ4v7kIQnwBaQ
se0qsD5vNaIRc6LUhuTXtRJ3HRK7ZBbc64mUqFt5xbHFyJoUzIvqL5r4FKbLgs4sPkb9l0/bEEXD
L4fCxtsuL59dgBxd2GYBK3gwDzhumx3ZAmpx8vofH5a3ReYDq/vEi2gjOoc4zwfKmViNLt86VOQb
JL9zNkxC+aByBnZHxd7hhykGBMcqBFZoU/sznU2viJm/XSfKiHpkPpl3xRrx7YNYJSbNI93Gmdr7
2d6dHqL+4ZfdgzyLqqodZVVvsYEsXkTbLwMmIgat97mI6bkNrn11Ak3Piiw1QdrHNn/GVBKtiOJ5
B9sXY2v0keP52a0+gNs4XduxIAf9Ino1T6etF1UZ7tdu9hlL41H9+J2EPnpVfNStVwuYViyQxGLx
DWWIrFsbIrQDYKzRf9zuF+Qf4U/srYIfVrbUmeFLYLMNb5Qifj7QpRMt5wOsKYKZUFXQWxICQ94z
XwfxYUKpe3A/hpVxl67D17C9mZpfeFDfznRLAZQrFxsFXIK6vljOV343ACDmmL5+AMeF6tSuQjQT
Xkkk627SxYrRkK9yI+JFIMtVhUc6RBdu26S1vK65N923TlUMV+wglGMrEavfB0+x3ZlNBTwgCZ0b
hOKwqk0RDsCJEWHbqdBpokhj/cM1yrYgvBMZdAEDTLT1QDD9pwyxNh2FHclLbpj/LxF6RYWE/788
eVzV2yB5JsCmczH0HWlpra28mqE5yPePteyc4uE5bSbrpIuMGPX2sI0hdQo39tJI/D1O5NaL3hVe
3fZDSchy5RlsaSBgtMPiIE4uNNBdeQFTE1X0umtm+44LnJ/toiSgevIg9e8IqIP5JpUe7D/Vqpls
BGADB82BDFEBKEJNgG6mWanodpgF4MzztMXqSM/2hJCcnXYC6AjayqtXNHqyqy/itAaxYHEVMHu5
YgfYdU5/lGonqJOa+yhIZSlB9C9pWAPSrp+M/qN6bNdcUtA2ajEhfz9TnKGLr+0LZaOf4NFbaYFJ
dMXjMw9A0j1l1FdvItOpTHbEDy3lnxp4dHMNoXTqqCyiM/lc/Xn6/y1dUQGrGtTokMwEyxgXMNbZ
lt8l5M4Ilka2ardp+hxabtVSFqlSV3scCAHBioXqtWCC3eDZPgSBk61EkYrX78t7JGH9PMwiVIDv
Z34W+eJuKo80tdUoFEPhaoHAxZLHplF/xv3Knn8KiP/Z9EcKzoCP6D7QzEhhb7rh+XJatEfFlBW7
HAZ9dx6duQV9AQs5kzX29jxntp2fYyQrFGR9aZiPnQpeWKDEi/sN/mG90kJoqxhbra7HVNtGSlwT
F9Sx47markJ6eXr4ICatPyeuE3v2K+VzOS3PJM8hCKo8N2H7pqcP0XluB4sBXC7qaUYIwlNu+7dN
wP8hvbIFpg6KO3sawcZ+JvbQfjocmUKxIQsZxEKmpIR2TOPj0nd49bbNNvpPV1A1nX8BQrp4gypv
Mq1CFSa/kt3XPmc8mxiefP2eZmAJkir47BAbH5b7lJRloy2UREyRcmC2Ho2W2ISLgDzC4ztn9NaB
qZbLwpNFTyqSxbMSN14MtO5Yl+ncm+JiQyz/GhAlTbaWB50QCtHTYEVgWLlSIZ71yHPNQEqjUTe5
m6zE+7oXqtJtB62u8m/0o65zw5xZjm9ria2+wB/qeInSejTAc74Dmu9rMJ0w9jZlVdXWP5OtvsWK
u+utpozvBW1N1L2LvMQ+CHfQ8G2ggYua5fDgke1zq5yfXwKRGoHoT+2ZfZVt3axvAmxnHSQE670H
YTyv+kKHpGiENbiqvrnKBYCcOYMNGQtjeOCjesZ3UHs4tKZLKxN5yHLKm6oBg/UvOEUo/uf8oRJW
H0OwK8SYAGpwwyfQS+qTHb41PseEn2x3nBSv5VWotBtwZ5+x5QERrWujv8b5NvA/+mPw0zNnpiUi
6zCMXX07jo6T4EFhJGekaK457skz6bI7p/PofZa2B6JN0Rr5a4k8yYT5PjqU8lhIf3gW2beza6gg
XAnIAhjs7c/qA+aGwdZpoxBFB2CeE6WfRkYLt+vCzXLRckr0FRReEDFRzB8yt3lfvH+owTqQNPx5
+zR0b2F7K2VaUkEMRrdBMww4Mkl+EZOKKJ72ZCtFycBorKYVJvYwsnF3Wi4oQDTP6ttnfnxyUkTD
0rer+2B5B+VGJPfkfBMzZRXZNcuBjdmRWpnWvA/CNlRW45Pf8Tzx8x/RXywGpFgHBP/LGPbHJSmG
TgVcssWgzHGY7Nn45Ngssxk37esJLTsFAcOWZHxMeArwQP215+TeYzmeR9JgTT2HqNKdaLKD9cUB
SKkdJTsjEI1bQ6epKCoCSxLIrU8wTqDAb3VQxVFAtK2pkwHYdFVw4yN85xf2PpDruVo8W5oCfnCj
0qJYF5veal6XYh07/5UgunCdx9cE53wraeo9i3Wbe3OqoYyFlUd3i0tnBJJbmXzkXr64xHOz09PF
S2+0vTw2ots0p1eJ2RNiFNPl14tdLFXEAX3nqmIDOydvp2ZItcAvttFLxCZcY8+YxQV3pWxZb/mN
++F/8WnKquf406446RcMEnbP1z1NTzo4pqCSDaGzg8tAquO19VLgaprN0I4BXYDFllshfqku762T
rHRbzWkaUt7MGA5EgiKN6+L/CvxLFMYPXF6vLd0XqQQ1jyD4YZpepsDNf8Xxd1aKzA5jz8BYRVPq
TM4nziPEecyQTFj+OMn9S4Z5JD3FIPcPmHuDN6SLhdNQ2oVRB1vkAvl4mHwkdEmmdGV9EQioRE49
zjzbfhvKXWtA/7yArLgofbYGQAqYzaLSyYaS4Ic11HwZqMg7VCqfrB2TmQ/dCpX9pCsMJ8UFMX77
8nPnGAHptKwkXrlJiBKrl9sL2lE0RHCkwXzzDn5TTKMs/FA4wOpqblm33LyuyK6MWuQCIEYBqPNZ
Y/d1pQEblMqdIHn3YTGaKG4Gw9rg0DtToOUMVTSChGNb7uEIABQD/+Gz33r8+iuCtw/I+Rx4KEqT
6jYmGooCspJ6WmHwLs9NXeHUc/Fy/UT8mtkagC1KIrvenh3c2NmRDTKvhb3BspledsmkJeqW6URY
HgueFC/530w8iVO+DwNWixliQYxp9hUHFDhG1f1WRNYk7BX9fL/SESRvt+0Jcd6O7uEClYHTmxFn
cO+sPB2DKFjkJou5UEHIzfBf+/fafkJmeVl9erpzyesBYine++aHpz8Am9Qz05zb7YgcG1HIwAOW
X8M3v3AG8YafskwSYWIZ22W7aYoTfnTTKswtk64O+oqE2UfCXDzDIoWKz6yAIlr2TIvlhpiflqG+
kVESaqsqzlIM8K0jZhgZve2j6AjLVPwV0w5YhWCOw5wa+H4Se/9Jg2TeziI3HVwrcEVtHfskegaZ
72BiPZjZ13LijgzX6vsJfwNHMFSDC0mIMreFeo0mdkeNXZIjvT4YLSK4c2of6ULKMt0II31+GDJh
d60noyMBVmflIIBuagIaYmq/9eivzdqWahpllKXwC5AAS50lASwGhkh2bBPUWTssDsZJnufENdHO
u9nQL+bgPiCri2+3gACbvS4ShYOAkjmTsi6vzWuTXhO50Zn/muvG8Flb0ElUV51NeE3mi77YsW5x
v6Jt6zpmfuMJWMmWgHam963gqawMvyCDUoN7TSHd057YOS2mlJbibi/uhmxD2UA0TvqZYxJECgNA
qF1Yf42WCC3CKf/gVIIhr/VXS4sMZzvgZqWQWt0d0VvnUAeXf5vKUJ6zHa7vBuLrMyZasiWLezYM
PUDs8bl7w7OieX+khV07sSXa839qEuuZvdl/ICBnQnbQC9rv4O9C5mQoTJIBw/ac2pUMwYdQkc6C
Lk1MuC1d6Ej80HwliquXBHge6A5dWfLczPuNwNES3nbtSvWS8ElYIRg8HtvOX66ahBEkJsii15H/
EZLzXqUqwxTxDVCPSkkxfDRGF5iQ4RpafgRnaUZjWnnVKiLp1+5SHN5trTAL3LnMdzb6j12E0xqr
9UtGzx32y6E47UbWHoz0wmySXtvZx5i6KNzRwYibs28shCnB7j8YOnq0ast8ORU0AXvMVmIR3wdn
eQM/dRx7VlFdHoUzGNZT2mnF5ybDmtvpdxKiEySIGDujs9S/RiGzEQCDxdcF3wpiHBqDUjGIzK5q
j/WUJd9Lw9ktseYaPQPX6vGTp06Wbbd7bkHPdv4G54GwI5+JMP/hHMzquGqvvTko0KywKd5T+aYT
JFrksPyNFE75hVFP13H0xDf3R0pVHGWktUX81KgDdNGQt1vpl1j0GFmz4B0lS88S9TtEYZTbxCPe
Iis+LSVo+ayXzqbQovMcxyXGkDsRwu5EHqtvcNZ3HbTALLF6HH7dVpD5fUhFgHI7PcOvgMUatsbi
tABXTOrTOKGGUbxVVDqyrmXmN5xo9IzaRumaje9DsIWq6QKkhXBRGoHSFtOeGfvy2YRXrlokC8a7
Yinmspb1nbKwW8sy6NP4z/RD8e5rsY5r63Hle/y+UB7Qg8veLl64khWQpvOKGKJmTjPevya4JVCA
3cQYX3kxv5U8KFACInS/4D1D0/B/ZmOctpzl43VMHcBFFiILGimIbSiwLZ13Sreyx/pbIRcXT5R3
MnoKYbT5WhuWLREHPLZ2PxAHsY19hHg/TVDQdCxwPqDdNUPIfRjKAzk+GFcwZ9OHA1RVXQBB2y1d
iPddBRf0mHO7Ic8oZpGtA/6WbyknJ2JHHjTGKKthg3Hge7urWUZtvIE4MNPF4Gk8g0ZBJDAOyL94
fJS1SpsOM5CZxBjpXvEZiMQDFqT70r7x5VwMyLS/xXbSQ4uinu8ORILO//M5iDZOuMTdksnfjN7t
EXq0p/ugnYTKq2SNhGmdlwkn6ZLQxx+aPSAuZKbvSY7VSEWjg1UYl6J7M9pjp8Kk98vZhiT12qEt
r7XKKbrmOAiiQaDKOAQBz4cFwSUztIBdOPzuhTsEqx+wflN69NINoEue6/Yqd3sTadVJw5Ju27Qt
vfIt4q2TzPH17xYhEMZ4xVdYFZKBC2g980q8PHgRDVpZ+L//coWZc/l3yFa+nY88EikXkwS3BoeU
DWBPfLKDJnrCPXmBZPMDEJMdmvKJ+QERDy6nbiSFeb1xtmvhjg22a6gkvlyfl0EjpbgHkPUrcZCw
Sv3OZQyZtIsm1yAmo56VhRB6cJhKPIJ+F73q7IANVrDpqEnpbTt27HlQ2iccXGRmGnurztG2pyR9
8ShJlVRBmDXEiD7c3Y1ry8E38YZzMF4Ar9sTcqmbKFkkxkGpFUF0JKC/GoD37R/m7BHE7PbKvbSb
0/5NMje5BzhO+9/S72gBdgDxCy3VlXqkmokZ3S4XLGkOrZlA4izP7zgwXaTgA2Pty7o2ul0snqly
02MLRtekuneKA5mOkWDUcdW4f8qLsO1sr21L6HhTeDk3wO4m3rShS9VJUSWe5oWxKj3Vz3AZG3au
iXHdJIDNkUCiGChXDYWgJH+bkcq91DcqT40OS+tEGpLmIMK8jV+19Z1wG2WkVJEGMkdfFpaFc8jg
FMZ53ONmilXgbH07xa9NaooTC5qLC56TKjWy0yPT2U6mvcWqzvTYSfJJA3cH7MOLP84UQ9QrGSar
KfERP4lAoVWIv8a6TghCOhUTbuM+bAv7OpB82kXfwydnuWlWSMxKUPgni+CUG9GYrVvTmf/uf2c/
61ydT43fWrgX2fDQA0vxl2JcfmCmRmyCurQvXFBQ+bbihIHFTOEf81cnkWE6Jlpk4ubbQlZADvJO
saE0n5Iv3H/57D3MUaxVLAHFJ1RtS1LYrT9ryteNp7rG5HRNh40xlUW86cjti0NDJNxoPAxOIIwY
/ZJ6aShhOuU9SZt/GT8x/9My4x2D5RQNRbinmPStOMsR3u3Far/VpVFwWD0RQ0WGK6kjU+h2e+1X
HSwzhBFufKQpIAP9vehLhbWuTkk2WFT4Sn9yA798sFic3NUTvw2LJWFgvdwXMGT8Ap9/KgiUDhTN
1n77+XLszhcDGb/CSWELHDti+X221X9kyDwQLh3f8ATU0EAXY2L2NUYOHmhVV9ibdA2eWnGjucBn
jCJgpwKLpiTjlLpCKwhZg5wkQpHlGJUDEky6dH8JJUegaRNHoHfIoScoKYo90Pav+COQxac33lD7
+fYYmN2+vB3ogw+PU0Vm1muO+Q93y9eYrublHR16PQyxg4/e/Q3wpgcZWWsGCCYjs2DNG4PLCbMn
FgxDPGnLf2QxqePwkmtpfuXZWHuUBKFXxoTXYiUbElXu+DW6kCIDjiSaplRFMqmrvZOLXbpsxOz3
gX5kduWuT97jR3HxZi8mrMrOldPbtzuW8O3Z+puC2vAwZNn1Eoe03VXlUrfYxd7HsH9aItiFUtzn
gkjm6VH5O6UbCrSKXpJXjKSap7okNZo6hVOU4S8ZXNi28JGnR/8gDohNRosYYkmh+ctNm0/P3v34
fPypr+pCk/GLZfhTyS/sJUjiRaWaXv5Nmayhuq4Jr5JNHo/03QzO90VBNRQxJn58+K6r/Nk1C2hJ
YlfsxoLxXHk3KxJwcr0dK2cuQvqavPjkLcZGedUarpjNtlsONxCjZpH31ZaXNgEDelqQT1L8ym8I
eXs776CLrbFNlQkvBpjyjmeeCEaPPNs8hrM24JM8nPYwEBSJBCUqFhemBHJH+x4opH2LGp+mhRXi
azT/Tyw5hHAjJKFFLk1IifXJqynUcBG0kh0FGgSm8AwwSE93Dfalcf7J1FkFYh8Gxl9Pgkl6YnGL
+i75WpuC3d2mXM6Vku2zOoQuaEfGL6Oy+EM69PD1ClAzmwBaDTYxGRekUYetdnPUeBJ/1tw/GoTN
KrEVDnkFUo+1jzgFm0KKuaXjrYY5t5jYj4Jilzbr31O7PDFeiKcRCXnW1i/EKY4f35p6nFvIgnKa
amKjl9UNm2n47eve2UsaGkqxZlKoxwglxy4XSKi/zsWxipo6hdX2CYmIQ9qLdXqz04oK00Mbbj6j
Qfh/zlh51DMaFHjxWK9gO6wJ8HMkN2WpFzl9XmaA+3bftAZSt5gQZ87AT9EIflmD6Qnm6WrvK8zI
y/vbAg7owN31l/divl7GRIAKyeoHq2nzJtGeQfDAvvK4rp0H3oTfDXeAOzDILQrGOgA51+S3pMCm
AmqmKG3SHXAFrvdFjNLWOaZdFz1RqcIeD7Ck7ZEM2TBvujqZDNMgSOwxWGfrZPEi1g3+XMk6fV7X
UjPoDoj7NJo5t+pkNGj9cZUn3HSxSbfEwdKUyXf5MekqxFlVp5gsdw0AUVqe7iCFmssFYe4w6+kE
LF1ooWDurtrU1ZpY8rcXClzixIfkofVdijIRIhu4fsIeJ8cAaXtWWE8KZt6c6DfM+08a8W5iZz3y
J+VT6QfgI/IBa6fHSL40Dtzah5oG1rsbwlxgmsMBJkVU7cFmP9VvHCV4jT1u8Mmq9lZWQc/3L3gw
ozMNtahF7mjdFdMbOBJJQRPAd/ZSkM61AhSa0cx8oD3N3oT+9KL8CyQ6drWj/y2s68W4ysfh9td0
gRTim9PEwPtGL4CM/qqOpjM9LWlQcffR+rp/XkudWgdWCARe3APg7+N4s0qAYzwN2vo4kvMuJeSn
EYEacEHivXqtM8v1C3JzPFXo8QSVvUc4aD6UnYSeB0VZjGqizKG9TGxpKNK3FtcRL0TgRYYPYSnm
XYQsBR+dsN3uFkoh7Y/buvCY+J7DR2G0ll3H3UJVBRea2KyTZKpE9L9XY4NeKK0WOxgfX//IUSM9
I1sdMVDbxn40mMpopVNscIsV0AtSMMYoc+B7NxaYEvx4iNgVlRMJL753UbUQm2ZEOvtal/wPIeRo
Fylj11Lmxwa3Zyj2i8hSJPVyfzrWYGm+AiVqs1yx+9zgtzUvawt60fgR9NTfvttOzQZ5PWRy0mxY
NEadElhoRNEzwzGY+MHjPOczy8V/4VlOAmCCj8I6kKbZIV9o5ZRkdV4gATar2FuBrrs+lUilFXlJ
563U66ro4SUNJM7md6EnaUk1graeOBqlrDizFfb2REWoePagQTp/ex+S9tJzzBrGNBC8mZ1nPZOa
oMTl0PhMvPw2oHpCwlawI6tr3mAPez3eNO4T89f6z+07cxva42VFh8n8/SGv+dM0G9/taZ7IB6MA
MK6adsi3vYKhk/JvU1ioiWJh0dAnzTEl+5z/werBfjLBH64TPh1CM4FbmhApCoL/5/mBbLEXC4hA
wJk2+i8t10+l/9xNrQWJ7JPD5pDVtDQ88j4ZQwwNMlw/+hsc8skRrFHp9NWA5LfVq5+2ST7dp+5b
xUsSEQFjIuFgJnpbn9QsXCc2iHoadZeulewwywMw3+6Qhye/ctSe5oYPfApM4Y2WNPIf8Gt5rV9+
2dd2w368dj9BPb3FVqw20cpyk+Vn3j61Yq3z6Y2+d4WZYF5wIqW9WAmyUkosPeVwnae9MlBmVfPp
WEaV8Gm7h78TRNgr6QTcYCGHA2uc1wR+xCa5wt1MLDLY5CE2RAoVzJYxQtsjExDg4eAdSGGaBzR7
uh717WEgv23zbl5uRnkmrPEZLHz2l0UTQnVK8y06ATvdm6as2VWTVMbTYmEXsx1rewEz2Fd1UBHw
QQZBdgLmLwbuB7/dE1Z9+5t9fsBCXqNqE+lWbyytDep4rfEr0ysi3gU8eUc1k5qqLeJVWJqbaOoS
hz1WM7lTx5zlY5QuKc+844DBcb23dcsHbxTJJnO3W2N8d3nIvPJ1ZQ0lBtgTlkQc0O8PchCkQBvb
V7Tesm5kH2pamVZidHT317Ykrw3tqnT78S07S5I5Y+PDRhtA7DtcBTMZ+MpQNNIJY0qJ30eKAng8
3ozbQTWb/GBNNNGv5dnE8B6qVMW9bo1jTlvmI+jWwf75O1ma5/dH1LLYcOrdw779I7JELJV8xpS5
Zj6oqeGf9AYlTPeTjZCwzuiUTMmrZWn11lmzGX6BdhrcR3SmASIYLS12gRUnmnKvZBjxyj2GQcbc
j7F/6corPLPzaVxKOgBYJqOCFb11Bs43k46fNOscwGyXvXcJ8RumSm8bg3PN0RJgsC2HtNpmHstq
xTNSbZxN8k17HqkMkWWJjbs5/blrjnzMq0TBsHLulzikUVpd4g6D5wP0W7eUmL37r70Qi+0I787W
lX5WUjbdclRciDMC6e6Zn86HEs7lKMPC9aJ/LeFoOaULvwuGHUoChX5yG5GBX2Wncpqekq7ayeBB
I7vIfIXNarppI7u64EFsHXHXgC/aYrlKDXDGXLrXwrygx2AaMF5REE+N2vraWtvNKhmdn+N6hCdu
OKXB7mTS8QPfpdPTX+g0atLbf22TGewut48h7SEGLsKnTDZJf8yD7zIq2OuNzIcvBRUwAdk60INj
LnnD/wBsrWuszFkc4JqyJDQpfwumzAKbctnRUF11YmzIwauJXREi72K7FC13CYwuK7IIjayTGxxD
aF6sDxz6kC2V18HE10JVsIxWMNDYWioYj6iW5TTXqVjaoeDGVhjO0s+Ic6j5l+aB+skjNKTbEkd5
r/9Yo0ueWWNLM3RTqp9hhngrOTSFMFcdNxGwWAjiufnj///pGNsSHQlu+Lv1c3KCWvTRVxWTJmPP
FdUXfxKCidaRTXl9yNQUgF3owFLUDhvTmBqULIOviWOrRkjfHrDHq2LLvSlIaUauiPVYA05iUokD
uKB4GuxPxN5dCg/9fBRJzydAFtAvl5CKsaTEbRic4KvufJNhxS77gz2Yj7+MmoACuc1z69h2LJra
PUlOl49blba8CBAdmy3xyFMdCHOiNlTjo5IYTBMlZtWSv8S3nH3B8z03sxJZgn875sychy/wZWTR
WA086EbXxFnP7mLhWO1jiqnOVXD6wOyR+KaLMVw8TbHVHqi05N+q9C2eaOM2ak/zXqgusbYYTO/Q
af7a/2aOuAdm6+6BM86/yBhOjlZ8X/yDB60+AwmwJ4LjsnmGpbTCt52SXzxrCMZASn0p57F3jPu2
Ven2nWbYYX41GTEXQiWuqeCzxt3gMLcP/Gdm3bufdAkoyPsaf0MiQJBA6qeKoD9+wWcqkK14H82T
mgYfPQYpDTWzkoYgqMBmAfYGPn2ngYAuInnCs/+iy8+6OfBx/zc6newtJPVbm2DTO/jw3cen4rEU
X3UUJpawCHwlyZfGQYfKWPF6T0+1b0esMiwNFyHYZxunhzqTqtMyy9kz8znvlKtvb4s9XOmFn3PS
KZUDmwALgCSnljhqkAczi1M9k4sMjSnYcu3ipQ/Ja0KJYmpl7AmGxMkk4HbvXXr6nmAWNb1kq+GO
UtOFrhlXatJMYNXuMQj4ooLwd4dZe9APNCPJTlKH2DKsuhefNNj/wypLwq4OVlAlpLjOTL5+taoj
W/2utUgt+QdIFlwRTYlF9oHZ7iGKKqhNhLMh8rjag34WjCtxn+Jmv7iuy2rBEHAv/0ovu9iMZ+3W
lTOaUMdeGCJVDs2GRtVQ+AiAjhqkKt3La11VdotHxJmZ4YHA/5He1RCva/feaAlU1Apv8Swiizt+
wry8SvASn6SGQnke/e9XLlYL9K/NWKEu09VFuidtGsimgNVyDa7AYc+8mUqMK25coR7wGZUiKIxC
/UX4E37kGyZuBqB77kuXBlt2IwOgeFIiXDFbuZQfvdmFhbUQ65Xd8tYZPoqQwT8e5VZWREsXbdNE
Wy0/2zynSTdoL//beQ9Tfy1s/eDOBGpyyaGtDZo821kS2S4kVomIoeKoZxqvN579oHp/B5TGZqKe
LSjY8qLhdgx/WlRM5XYNCEFA6NKYp778lQnMLefO8UfbtMoC7/0PALpAq/xeXhg4gT9G/afjUCCw
vP9zKDQpYsiKYgQsTf308SYJSvBjTQIgoP9eKopTLptoX6eNMfHq9H2qcAToSiJNKw883n60hxXK
p91FzFGsop/SceLkvSxrgEDXvn2PCA8/XvDTm/B7wllXBpkfBzubp/UbdutMQ5vAynUgQcE3gdtW
MUMhs/+0+sG4MCsTuwjLRmIhATjPZzqpBPGCVzrcu/p9VgUuI2eP9Fq+v2BMGmTmJOaxQ6xNb9JP
/LJlVNJNvq9RbKehdgy4uEjhj8NcLpPnBivGWtMLxAe+5DezO6ycfUn90qaaAvxn3QxxAPMybZ3x
4a7LV5uJIDeHgFZwtpR70Eqz0REUoXCKXh/3A8VJCkLTYio8PWYbmmSRJ9hE0WoMJqDG0R2hcyl1
UZco9Hmdlev177Z+Rdxw57UBPzYB1zFr4Hk9fVmpffh3AczVMU0sy0dKoCxYVlOQTu2Wu1mkxYWK
dgG6ZuC+WIgfdsPhTctvTNDyDJVSAvKLA0U+6lWY2eSoOZPKa3zzsDdWaeYAk0ZOtgI7njm6cdp2
AFutoKQcgiDIlPaVJx93MfUvbuvErjx0MB2I6QuKB8yZvuiL5yci01SzptOtkry8c+YnRlZVGoZZ
20Duaec5CcaRF0WSGwxuRJ0iL81pQFGVzh4CJd3e10tg/bFb+k3mTjUeeJZo3OjBosq1scOdyLe/
PN3XMrjrRXksDEK7/LR1SAzDIgX6T2OpR8pfMnbnCrO9eEGRgvAhPAJyQt/+kBwS2ZyhE8ZphxV+
oDAZKH3O4xZQfjHExzIciXHP4PTq1y3+8+QRdI4SNy6Iogq85VWEZf26TQTP2jQk/c1W2eUV9HGR
BvV4pubjvpdizw237H33tuHPc0q78+Y5z+X6n06R/IMdGKYsczW/bK/j0ELlpmyRy8ePk7j74zcV
ieZA34Tkdp/pqeLNqXa2Wd4KRISfTRttvzE44FSy3OaJgo0K9u1GOGipdpPnj7gIZySkdE/i109q
ZXpxX+khf6Lxgsshy/9ZukmY3JEwIxNFlRPMdzYrPtAWmNcnwXLURTLKOGv1fIvLahRAMmlnfviV
X3KaMw52O0oO9nWi7gDbQFisw/wCBy+lT7JI3E4TDEdhR4DxSi9pQCE6CcfAuAKxr8KoS++D8Lg1
M+s/SzcAtxlg/V+NfREfLtU3SSOPwP2DMf0xeopCEST/ZGqSNT1q+UIEL+6rDk+HdGaDchuExVsH
1+xscLQknot4k83TX02KFH1Rf47xDNHYTMgdqybnnvlKzdgLIVF2KFQCIf1N9T/OUfhoGNYvBvTH
FUeduYmxs16ZRj5Lp272kA8ErBzRyUWrHJHIz5NIfpIC6ihB7wpTb5bUkg2cUZ93awsXQKmhY+K0
EvGUNODBkTVxVMgsbZ5lz1ZvuPYAW4GrSBHDHEUZ2sd8a1kLw37/B65txrdD1hOy2/dXziivoFmJ
BQ0fJij1erM2HRAu5p5au/mMduaqEIw/HJ5yZPh9tlvfsjJ0ovFI49DNzm+UQhCznb0sPc6kz5YD
90TapxSIr8kuQNHrihIOuhlCv9e6n4Ufn1R5t2iVc69TVvrrvIGZ9mV1W0OoPSzw75Lo7VBzPKPQ
nwUJJBRYB5bNNyD2cynIl7vKTSUCzpQatKf7OurFQ0S7GoAFFEAYiP0LiiqecP/jbSumyqGoIWNz
0onSdwdTYZawcUSyY6lI3SzG8ZGYuUM4JbIF6K4rCIWJoN8Nph22A4dPc5diG3RG0SuFqlohR/U6
pE7p1K8A10HxE4yGZrShBdmZQQFYwF5fSI3xoQ2vB0xt+vWHMsg97JZq4mC3N+OdUIxyAoGG1jSj
YgHXVcI6wDgna3sxgu8PDUDgkF8TfjtD+pSItETugNJMUA817nhdm+20oyfLHsknCKiyDvdI7iwW
S4oopKfYhUKfsK5W6ocdmYR9lN3+rx0+pVNWDp7x60lXKMO1A6aH6ta/qDMRyfkddQi63/ItmYcU
2od8ApYe/l2uTz+2DxaQH9olq7kuyBjEilVbIEy99Ha3mif4SSLBq1DKPuP3VEf17qgsn1yDiAt7
UVSdYc2MScfus2sfsK9wvEbwn3l6vq0iqxZ+oouVq60IzF9TCC+6RjkfV/53gvVevvwwOc2VBTkY
9ApURDzPR9Pf7CosI26O64G+lmKp3Bxe1j6B5TkmpdpfhPpcPT7qmNbi5YfJGz8b/5v6A1F2x2z4
utLRz9/ogi4vjWy07fK4QEsFMFAvPSl1dNYSDr6A2Jcq3DRNDGTADF4I25dqz9/IMdS+RiELaHzh
82DUebAdtHuH6Wbb5y+5/yvYnKyTMrgfu67rc4UomPwg6JlwU90zoJJXar7CNNogw2qUjSJZ5b2c
2RlKivT+NUXcpVxGH98NNeuh3WJ0teQjR8rgA2Iy1OAhC3sJkCSN5FpvyerSrOooygaSYGasrXEc
R/YPMsS/zYgDzLExFtVMAhCSIg4frbp29BD8Yf50aJJ356axd3CAOyG26OIHYlG68WKsLxx87ocU
OniJiLOXD5Twexq35CA5tTbFIKiXG5bHCVZAFlq6oMhu6HUS00fuFSaYSAToVwjYpbPuGwiqJ3zP
g5l2g4qD+rAphR7csEPsNLisPx5qcd57oWxJ1LimXbId3+pjNmW7rwH+GELPFCbt7GsxqGqCUGKE
0xKaI9PBbkuw7nOudqmM+O762EWKB4vVZvlI2EuXftGcBSxigNC9Hi0AuzwDlqevi1jLEdC//2YO
Zv1SLj1M6AtK4CjEr2zV/H8CpCBCPlePO4YQQNeiVIBqVHzD949lx8peuX4RWltmrImbgnRvBwKJ
YxAAcP6wfvMOuwH0MsyzzUD+8YBjeMwdacl83EC0jwuwDSJZSkeQ4Kjgxh0NiRxY8Ft6Mpdun1zE
OGJzBwOoaNTB/73ocXqanGfWUhMl/Gznjixv8jeF/DGA/O5sV1DfFcx9hwoHh7EfPE7ZWxxiLxMP
PDuQoj4sGhZ11lcR8mUuqNawjxpTc6rj/brXBYTjepbcvifVGGohB1HNRaS0i2OksAgbNBtJKooz
tatmEpHYd92yQ0LBnxad6ufFb/wZWKMs3r8GUvu4VviL3YwQafqQZqhwdoq8OOmL8yFEF3sR8aLK
wpL0gtJAhLZSgwQhpjnLQ+DAqjuLT4BaBbBOdBd1pA8SdiM6+0JOAAYIaUlI/b9LUKVI+mj2m7Eh
HYNNk0Qc3oxS7qLFpRLSm5phMBi/lYGgk+mPnDPFDospaFEdhRFZJ7yMzfpRCZe7yuDCAF/CSfif
xgprbI+NX19g2qQ1HiPRdsKmBg5KXAoSbJmBMifMuRsLvXjJsCoKh5Wc2zLjN/9c8n+/Uf60tuVf
3Z+9JY4NQKvgl4vqvRPTh7dlsJU7IfWezzh9rY/7nt1GAPFBFaONg1gtwUyHDGcuSmskB3lsJyWm
gUPXFKGbGIXE3m8XZQDJtZTkG3U+jjKGPEku4m2TMLHxv3tBWxXj9Q6yzezV4+EL77I/d43tfBJp
bxXhDx8rQvHhs/rV47IMozliiCi/fcMNIvLpRofOQm3OkqLZ1xTonK3qhLi1WetDbwf5ZsJiXeAi
hI17bmW1SKwDEzi4gQjDpMLyN3k39TKlx/Vx9VkvrD21yJp1+NUDQosKmlS/cACgjktahap7Jmo5
M002Ghct6IiT9218568LdyVdWP/dgjaXy6xzSoP7rgQyAM6iLPdB3O6My4+bL09b2ILRBV4i5dds
8TJRSy16J/TnS7rbg/2nR5jnbz1lY8z9Rqc4GzJA5/kVMdoHHIUMuBc3VqL09NblbQ81gCr6DN/0
V3OUD+pxNbUNSGPp4cEruuhwzdc59qxw7gp8panCOwNQaZnz6kNzb/xbeP9gwuV/R9I5ttv24qIb
A0l6WxjaUOz7geyfYTV2WmVamLdFpsoiYAXTRbPbQWAzHDsUBnTO/QQKUj+zGESJnQVTkfhzBigj
UT+q6Yfz1xe9GqLAJyCFVDr5LYMBwWRLL9CFT4UM2UajwOLua5n1AB7HFPzXalU0qgigmL3Y/Z0M
gheVZNq2uExMH3Deg7Dl+TwIntxzOl35TijRQApqAsSbX+pGHI23SjenOOYRbaHM9oenqZtetDQ8
hhaNm+4qXmyh0igEjav8R3i2bu1lKCHXlS9RG6MflOjDBmK2idfgiwGnxFSHn0L/DCNtgdR26m6w
CCW9sQFIkEw8U0sTP0RcZKHBxg0KvYSYizo7e/9pZADKOw/0PiKVNDy5AxclGyxhMQ+0cvGHSJD8
hxfMEeOL2Uod2gn5ZtBvx86WbDiP9j1VIs+MR+N8zXc7UaKqQcYGsIVmhvVNFFTqqPwNH1+jXQFY
PlFFnNIXTN0/LycJFzXn4rv1MbATfb9iXwqY1+Mo9OfXC0q8iRhAx7xFRmCkSziHmc+EYdk0dgi6
w7g0wawmYHvjIej74xhGezkIndJfxoGBS1ff7yQ2ANYWycHlfUKNw+T0ZqFrW8dWc647+6x5ZUEC
hKAlH4/9swdejeptY+umSGohdAp610T+osDSAsERf169GFuNbPu5JH9hZho2/3kjQLdotI78Op8n
HNX59ftavw/IHdegdSpjJhHkYzEbNsn0vaAZypWtgtZ6Zbb9qsX6OEn9B1w2U/32zWVqK4OGadqw
Gi/M9pV4V5VYqumJzaj46l83wkQcgSdbxLuQBQ5b0ksm2o3otVGOc7Qu0tfpubeR4qwpF45Qz6O7
AZknhfcpHy8o96tTC+u1WIBkRv46/MyvFXUQKjHgd1dznnqEG89Zgn/rsmsgozJAuxor8WVe0Y8R
rFhhrZlVKEjv+sSpqrcfBwOH+X5aWtln7NVNW+uM0x7bMOetmYenhXlkFXE1DZz3bBz/WhjthGgY
75glJcMKX9MHD7MXrB2pS/QgfbzDsU2ZKTrw/5N6S6Oz6a30M+IlDDWXkXTI0vE1j5ToMzv5gKT6
B+XAu7JfORWvReySjeOAFo/RpgHbYRRxjNlj68J0wuaot1XfWh/9oIFLuZD8lH23axzM2O61HzJr
IXQcLn8MfVsHM0QdtN16H2L4WRCDjUdeVrnxGkrKNZdPK8mPNY/WXBIPGKBjmFzbkxNFai4bTDK6
niMLoarheetIg4hYpGpippxxukut54XHq38UYkvbM8O0qnqaR50paiVM2Qz9OQekFNwCToOwEufV
HQ4g7rLZG5J4qQoyHINvTJSgqW5UiZlTk6SvEXuD6A3YAFowc4y8GlQT7WtkpHRl9Q+E166HjGOg
TIWpWIN1t0qlyNGlEcLw8PXqxf8tfoaXP18hoEGFhDpl0ie+1g2wf+XMBJ36mXvbsJo/ARdpsOD7
rkyll9mB6g8zrwXNihb08GnIBeJTx+pQWITXIf02kP7cEh8AbhEr/RfgOvDnXOYJf2CCXpCZMT4Z
TZbqKKEy5m6SgC8SBEebSM9knnPVgYOlRZ7GiD6eWn2E38RSOTk0ODXIeqlNcjjCIt/oH5HMJ1Md
91y/54gDsk5lIXS69XEE4Wt4YXjx7yKOemdVhOgEVjSYpHWvH2GXJTAKwtJABHrpeDI+SGm1cHYu
L2eFXPe/35ldtc7FIrpStUYrqZQPF35NZghSYJt8hpfc/RRVrQm0KJDmP8MDFVCIQLavMl3XySBe
H06V3Pzu82XolPAL6AExDJg7U8D5y4SSsnvWV1xFPZsi/7JqKUnnrMF0Zjwm5zlUtvkeQa9qY6bO
mk7BitHa2PQciltFY4+LVlEp18l+yRfXxnWNXystDXStccmc5Tf3ynuZta+/afJw0CX6cq+nXDo2
PM6T4D9a2Rmt0iuPE+PKzZHRQh6jZO+0+DXDKcdsMQjUbvjZkZuiPVh/hddWNBHl1UHHIZYfCha4
UYnsFUdPmBAD7ftojPoRgoDTVFSlmL8wge4Pj2MUfnjkfIXxBEu4WkOqJ/tIabFBcptsefx6RPcI
/dayXu7VkotHJgsXU3CKeeNuemvRR3Iaw7I870JwmZK5f0evZlESrXLVE8XpefRlsPHnlABb7xzA
/ujBbdQC1yPH7LKxd6aECwsVvcIhiFfwXpOuf3EERapMr/HC9IaPEXbapf31J/h7JqiBVepeB1/z
pkleBUccJep1XqvHO+ErfWOL12txEZEtmd2C+6BcB17sg8Z7Yj2+3qP21C0LfVXD6VZ5iukqpIOa
PUUPZPVvT3EnZBca89J2B4BhwPWf5IEzw4XEK1k2rgO3xmxdF4aT3Va6Pe6h+KnR9YVX2apP8WcX
oDxHfh3kCI9YoKkqnKQlaS/8bKNZ255nrXaBrZT9ZWC1QMw3xzC8LEiwDFZbqfiNu5EA+HoyKqyH
/HLLs0ePfzXhPtaNX5+mboxhYaXkgUQpNKQhx6EEsIGfzAddHfBkXbmJyX8rtBcguslzQyAxDLl+
OlB4DP9w6P6q9bGe86T7DPPHywTl/RF03d73YLXov2GwpMAHTrpa1jEw7Jq59mThOeMxgeaan9XI
95FlCBGJ0pbxfs9TNvr7AbAx7aAcPexO/TnXjaziVXM861QCb7cqj4udM5+NilegPRi3TdpW7mNh
cYR9jB1Xprb5s/RZQ0Ho6rR4/23pR/q1zFrpJ/q7M3JvkOW+oX70uEkiprR+HB/Z04/XfGul/5fz
Jj0JWg13To4ki0LMcFJj8eMolFSX+V8zid7h2bQ/R+SbGpsmgw+IAQ3Upa43VVp+ETZ7eC4QOTo1
aEWccCRTlnndBLcGe0fsbRTD2YzmdDITZ+w4k2/DgEwy0fxtFqdAcOqU5P/GJgl1J/qI46V7YZTP
hKdDPbkKQRMXfcVWH0K7EK8Pjs2w1mxdz+K4Io0i4iF3CXDpwB9FWBtA9SyyfYZdrm4ksTgvuZXr
zcBAgeZmYkcX1fy6yA/QMW+0DzufPS3Bl8met4IhdpGuMGj9fZdSt2cC9K37RlY7/TcSTshIZByy
4zEI75oF8Po6fulFmIz1pU6EzYUW34Pd3gRUqqXxotsv5xiaFwylYIsYoFco2aZuJvSLaxajksZc
HnhFTp/hF9e3lakdBMwlgUnVBo4bzmpXHJ+WwVkzwDKEiJFh8IrbO1ynbLhtIU8YkH7ySEOXL8dt
9xMzWlSsymvPv80c6VzyDBfKkFylsLVLdVnPJsFk8cSVHzRAZzT441fWj+HjTxRDoan/snUYraqg
sJnZDlkq48GXmJjGO3FzOpov1k2b1CiOhdssh5/O7SzAjhycb2DvKtY6RbmTuUEHLvou6fQn7oXM
os4XYO8IVSQ4jj95/xOQ9M4KjU7DDSwGm/ILthi9WJDxV4JXjRhDA6BUQSgl5uKJhf1Z5L4Xmthr
+SDFxGXF733somPMNyLZ5z/MfOwaBuxTjk8exFTc7DBRMg+2m1UaZaB4ZbEb1rUiAK0CSOHbsYCX
o4q5RHguFJfIGUMGpLISb004LC/8jT6OibJaZf9IM6+wLwMqyN9CzqfbSuJx/dVmCZW/UhKoAYV3
eu14esg2C7yifPxBYNxtggYyt2tSPXkyFZ2MdUWKDEOr6zVjSIYjQ/jREIf/AXDGpqsXnDpwd6Mw
eyFHusSWEv5UdPJEUap8mburke+/jtIlCmdXnyFG4gIdGICMahU4v+ZhXzxuRhsjrTV5GrSBlYIX
oKbW7jm8V0K4bLePFAYyKvKveiuDYrYuOhBgQf5au7SoE0geglEJkX3kWs4wwLSlBDmfN5q8lWUo
QT42NCMWqM9eUIpkPVj/klR5F1MtnTY0Y085NrfK1jS67ER2AYndDN7taDuSkKlc8+JKhiynPY1y
1ni8wpE/F3rL6WCs0deBzz2osY9wx9BfLesEM7Emz0ooCkX1IKXwDVNyOJ7wACabHrXZv/PA3HLb
tX6GN1jT0yoxCYSu8Ub+AuPhbbZN+SoGXTB2e5SLZ8AfuwdY92qMgLQeN/LC00twe8OyLr8COsoR
f4d/ycHI+/K4Orh1bWgMFwuyNRe1gnwXy3PzZL4JSjehtDGx/jLEIB9khdlviZhGF2bGILtRHvqF
17vE4qqqFenmMKWOIB2dxa1QXt1kavTYNT1r3RyGT/pFwGo/Pvclq7y85irS7rYiSIJcodSUXn/4
FRG25bEYZN4NxWCpBsy44G5pdAAbcRM/sG8u0W199EpNAXVSOIYyRzvEFDEWuPdA0a7g8j5Pn3k5
xOJ7DUyTp+GuovbfyDWMU7kC0wHh7tQwa4s2DZLkpTs4iZ1zi7EIF/QYrSfoZVDzH+9m/zsXB6vy
Pnc72Et5p/7qxbDXvgsTGly70gmWNl9fI0pzydTuhtjm3UwJy7yGDtzZo1/kkaKkrnHEGSUX7wTJ
bTZVxNW4VDOCG1Wd5lvDXWESOw0K08+KD98scGpkzzjZgHkvN/eeumNdCYC04ZjywF+roDTH2Bl8
+0DJtkk/2F+rX6QYFuPXrMqardeLoQw7qzipKxyHubIJZZsJtySUNtbK0DUB1oFl95jPaROWkIv2
/ze2dmp/ll8P3gqVzj85jTtSEAa0beee0Z5rj13d8SDuDeQLTrhPfVx+cIrKgjozBuP2NaOmQCOd
i9AXjZpBlhdaOtLkPSTGM/x2RAwAj7KnvjcSe97GXwIP84GJz172SASZPBmV7cck/qmIbfDo2ULv
FvWuYG4Y8Bmx1qJOQAIG4LBGyyJ/nrqECxSLJ+ZWtA3HfKzzKZYIGFWjZZa5Fbpr10WQ8RUamhn5
yHWvpAE0ChjLSauanf4HGwk6OzQDwo7I4K++kjqDAEyP78ZU32qSO+bGvvqXDNE9KmOtHkXTN3Fj
xKWduU8PGB7cGQjY2+i8Bor3m34kIYfl19nK5nSdWgp6cWG8ulsT7SngxxOjVbE9yW1Qcp4amFe3
WDeBvR13cLjb7jR/aIt8GW19elgm0TEhzWTdhLK1cE3gLYJkDnMXuu/+UAV44aXKDOYZCZGZ1JsA
vcWIvm+iqPgYa0UNG+DYq0TBiT9tiNnQOzNhfR8JQEpgO+YISop/99Hv9i0DboPhS+JNnF8gP9ff
Rh7Sikv+q45YynBSrrzU4YKShMoTZurgH02P/Ix+DR8tRwmUGJRaqGhZeNfFWhivRPDvzz/J+kxH
6vg+j2FoJCS1rgi75FdlaeA3nSsIgbbHLUPw/ly1i0KyY5qtY55QzAaXkur2CBYZ2fAsUG64HvQ/
FmBRkdlK3Ee09oQdpVp0q/gbgLyp/ix0HcjlezXOPqlg5tbR7SsPAsynq9G/ppShzy5Xbp/vdAhG
piuHq0cEHDO/X3PSPGgGzevJajgREpR0UwgJ4ihynCIEVXOiO8NP0DAw4Wgtf/9PfVinIFjfKMvq
8lJDuLqCwq17Z4xwAYp16EHokXYgGf3hym+Z3ZS1ExLs1icwGy2JNxpzFoBPbNjsSKxzE5J2BOPv
03zqdvigYM185vy5gtgWIxdDc81sYu+na6yuYQddanJB/nJcoyIAGHvQmsOWprtHHPrCl8I2yIeS
aPPftOuW8Vd49mAx5HSgfQL1iqglHGUv6y7mksYE6Y8BEiZWYKAYwUf5PcPPvWdcqq7tRa79KYuK
4Ihj72eqch4DFH5uCLxXRSI5JCg21WLUWoRbh4x22cIEjdZMcHODHXlT6mAulIk2JjJtBoTyG9R5
q+BORuTzZEfm7+8TrZJ2ZaKkwQahvdPSjS80OclvP76IIFAEv5b6WldBlEIFWdUjKeoSL93387tG
8uyx81uVfhaN+NvBeT3kQXJxALYWqxxTUyjxU9uW4KfVxasu7ISXn26GFztczCOxDge5RErQDmjd
/U1leLGiBGLHoUumgFg8ALaImOEWaxpQ2kUo3Zj5O7QXIxfeMs49x6s7e5vD6lLduNDofqfSVTlj
X6fLr0amFCViaGvstJNjLVpQ0QbZA+1wybl3FB42w0MIsCBFxnJLg8DFjM08/zM+Dv1s59E4dB41
INGb1mnfEqBwsOeZ1cPrvXMWnzUn9UBX6AMpS/J2uirPMRCncHl3qcojLzHTMBVYhmvNY5VZ30vb
WusIp+X7y/XZ64LGN3a1R6IxDRMv90o/Fm6CqxunE9FM9/qsD7kH8y4Sr1etNDIuXSdeZqIfQ/G6
L5MNcz1+IWQ4JImx2WnmB5KY/ith8mib6FaK5VU5Vr/Mx113NV1JijeHEZLWLME7x1ZI2uAnrYvL
KwlOpBMaOYxqYwtjqYT2JLM0ZUzfhcqEruiKAn/n1XkekGOuzO/+cRutdHoPPfhQ2UWQmjb7QGzg
V+bT/sPyNzf7C9Us0xynhFQusJNfW5gU07tOw+agl3IUR6NrzJ9M5Xbz2pscbbbK7stsrO8YlhiZ
Hsjxs3wxQXmgnGaxa3cobhC4ebMjyATzYkwSR0povw03P+pLteVf8wi2EO2XwQh3a8MBJNRl5CgE
oVT33mLRYBgr2/1e4cvJYI7eZ/8WvMIJTMQuVQrDJr7pcUnrfZhcCotkeTJ9MD/P4xRf8nKy3FTW
V7DGHd2+9AWvUkFkDAHMp8ow5Tcfe397iTE0Wg+K95OzoU7R3y6WzkT+GFVCaNlFc5FYXn2a0X1e
FfuRJjsvnkTAl3xCuxEFoYOk3nl3nYgVoNTBnxaVxe01RfckfUsLU//yjsZu3n7lQCW4voZcSW1O
GXmNAZ/V6T3PqRq1zeCrt/qYVAl62fbbOgLT0eTs/8QmaTfd3GuWcB++CmD+QwqFbw0WoAkNlt7E
LkLOLWxqnB3l/4czblZhbqwqTnSG5b2gKPabslbf6rFsRPlSinjc1eml5z0gz7m/JQQ3qeJfnHaP
LnGBCZdsQlJGYxTSNJVLuPj6YpMHDNI8oKBnIsTtCS4j70iUK+1vwl/Y1KNrGbtXgPIxiLgmLNs+
6ebbfBlGcewjXFj7Y2McYBihZGvHlKgXLSQz3PyXk9X0feDoZm8z6OC5Fz90d1YoQC5tOBWYLVfE
NpHHiItWmGOpYPEkCFot7Szm3cMXnHUL6RpDwTgj37Ok5jLDDYUya1Ob7nJCGCYWY2raDH2nJ9pq
0DLgPaEUYQBtoEgSds77jFJ/0XLB9lbV9+ay2syJh7EqIDSaxdfEnOshes/S1E4Pb3b5u17xWJXQ
eDZOvjZVfATKD4AaWDhFT50WupToq7ShYpEeUC0TKsWs4acHonkHkE5vSdaBt0TyikBJFcApCMQD
9L3ywZSTS3hKOK6Z2Hnq2GVeNm5H26OzzPZKLAHtF/w6gWHWRv0F1xJqZWzqrV+4QYhGDkapdviT
qE6l6PNIq8COpjqsgHsb6oYvsGpPLf85vZydFKokAQPYJJuhKP8lqN0F7nTmwVE3UE/yBWIkgS2r
RTLg5fuQ2sY8FafOpyQ96TQlWrUx9qX51W7Owv1Dz4d58lEbLVcNesvj1prFP+fSZloeaxcj70gP
q4htyAHZyfTG+WawzB8zmOkEbqkNcn58xntozWF8Ith8bPm+y9Cw+jWrMSqAj4/MzahJzNdcDvn0
bPImCp7CVjBZoKCyCVRsh91lr/EQnptUvo19Xwbaq5g0S3u/9V03WNNtfabMW3c34H0BOelRKqkQ
Oy9iOF2M6MRrkoZ4kce5SKjPSkNt8HAcKQQ6N3iI8BoA465QtA9T94j+M7t5LH8Wz0KeKA0YBeOI
B9psCuDWliPC5diwdPkYclzoeLlXta/R15nfx5BO7UrVAfHJhbbod2knEx0kWvuXO2NnG3zZ8qqJ
4UWsrRdyGNmirfLY45/zMpxZEOXFlMhIck/5ym39Ml4qgvA6wja7hetSVOpfxrHB+3tGY6jUC7A/
fP/T5R6/ZfGVC8Jl2DLw5jsN0aw2CW2QeBNghNn6EMe2j7cj/f5FagkQmk9EvQUs8x6MasDG05Bz
PT1rCawPpDab05jW9crPfXQi4MtdGocn8TwDiWxRCSFd9p7E+sG+kxHBOzDe1r8E19/9MLJMGoHb
x+yNBU3+LeImfrlKsn4aC8nopDbYPcsEkIyAKsAzXnyn4iNE3xTt0oD6m4quGXgkp1gpL/deqK0R
SRnl1exiMkckMRMrs/3KkEb1a2p/6iTv4hUr7fcVJRxiiws2Uk5noHbjTkwEVJbNSMEAD7Aqw1SW
LAu/gHSYHT2kse47Jewdi7Q5frG28/2wBAldaBpAt/PZmne9pairiiJCxJwDEWEiFEYCURnOYZII
+Pum+bmo+eWO5VXco6GW+TdJBRyvZne9aF48iwd/aYrciORwMXunMEXf2xsq8ECLG48gTOZtQ7hU
TfIKCFhvkdZ05XngNCF3fkErRpjqv7kk5Rwi+c6GUZntx3j1ebHspOkcOnH0+AQbNbSNMPnT3N3b
po3g86Cy8i78+qIjsL3x+055Yrq+K/MAI6+7QR0HXKAvmmIeWYGCM6FtSpyfHAsuUmqv7l/9A/rG
Z6hjZHaz6nQOyFPpoELeTUafbySvM3G9C84n13yU8l08G+VhHqg+WmBF/8ruNNQ4F5QQdxbt/d8q
op66znImz4VGJB/Bc7lN6sZ876h8cUCfrjJh7L8vopkeglw8wclF0gwJpBc3QBQ37oO1NpSftyc3
o8u6w6Q93j+LUO5UBOgFPJ7PwAAJ4fxTTSr0fDqGylcludO4dBUgvQonTX5fyObKO3wdP/NQ1/xL
FC7Jj+Bi729Yy2MwIvuNmIY+z0Dz0Tp5KiPcIUhaRlvcaVs70x3Tnfna+fRVc2fKRX6ZCzBGkdmz
MTOqzgVJqk4dP5zBeAupoN0GhjQgsMG5NA4y/3AE5rX8dv/BYoxXcHpQK9TvctV3gd+yNXag5Hno
rsp4FYCzg7j0+0I15njV3FblJChR3JysndnmlOcHUJSDkZ3x6rj8un5rHP8RtpG0dekX0aZtXQeI
IU8ENNo3sAMaWvGuxybLWThRZ9phqqzmAykDG/vAgdeK1bC7fKtNgx2JQewG5AHgStkkDai1esAk
vsyBR3X9r71WQ5FuTs1NVZSGsAMUgx3klN2S2NfjTiz8x+i338/MLyoPm25ZToAGwDXg28zQ1TGI
X1QpJfN+19uykPMJQNSxUDn1e3RsZwan1deG2i5XJ55u29t9iRIjtiqwyuJhhrvePOoZsurjAIKU
JuiQWEYJuuGJonHfqI5lfAwmZE5gQg7tlxqlj6wMALTzfQeq4td619oc0ZNtjdyttB0j78eT2psc
klW1WUpUJWPM7fZ5aOtOUTVQWsHprqyf6gwx+bOt2af7lQPBmhtyvFDiNRL5vPyUwYvS8LrJRPrK
6DUU539xjKDpNOVxTSTzcyuuQ05nckcE7Ln1fFA4fiyHys2d/VTO6rdboDrr/S9BylNtu1EtUH5A
N/lsEmzQzELXnAIAJb+Xl1yOFHmgxzDsypCshajLnse3KkD0UFSh/hcNqP3Gn3bMfkYo5UBvWUsR
4rKbleQU/2WGO1agkqCJLjKA0Ov81E3iXU2j6tnX/YImjq132bjGmXaVhuqAG8XL9NZmq1kaihrW
0PlSZZ5h6YmsU1bQpVDu2eIWOXR+U/vv/2G3wAC0mJw1xcbnXzJlOUn5D+bqpG4X3kMcahc42cr0
tLJhlExZ6cKshnF+g0nijuR+00hlXiMSWvO3oHE7vSMlUOZRVuE/JhOyRT+x/VIFtWNtQnt7rDDK
SrCq1RgKOjDORYTkdODZnYt3lDw/8H6mVnMT9gdsgM1EkgE5apkIaLnH+oaqyG7HW1TQE9LIAgu3
es+Gp39l4Z8CWZRMwZs43zPLTlsxjMsfnVDPgMVJcTDQBYDUltymNuMeOdv2VNQ7MXVluz5U/R0w
DeV8SQ1mb2kk57ue7Mp8D71h1jdNbGb5AbMEAw99lS/2e2K3C5BZ02g2ZjYCGOSRAxSPBOUeQyH1
N/CRvO4vMIxWLPjP4WPF8xO9hqQQXQL2oRzJfXZvKtLh6AhskNRzKMUfhXYkUkq9I2+BtSeCQXKe
tK+Hr3XKFcDmPAzIVA/WmBdz3yojm2C0m4RK5c1eFKh9Ckm6+mcDix4YRiHRHJ8SHnv+bHRzZHm9
vYcWwUh4G/FlSWK4OLIF4/2+zxrKLXi9Vx7KmZaCUaeQsv90ycUv9wenysntgxFzmDyay139z0l6
7V7QtCX8x3W+0FZi+Z316hP0ADVnUWmHBxP1pGIZpigGVzyRhhECgooN48lIgWFMkWWp1HvueeR7
we6CAyEpojS5ymUSCl7wYKjYA0HXFeNi0BMPwK+tlDC8I/6PlSGtUEvJmtyXTRUHzHyky+aJc8H5
Y85Qmq46LMZVVv10L+raAOMPhqPvKGtdpEC10xToTkzQeHECNifFBZCZXZrl/dECTXgi6vTbVmsc
iiHo2OFzs+ZXuU6P7q6K/qXbRJNWZ0nUmjpS5nJmpslpdKno3QhaJvPKFraL757fK4B9LnI4WkCj
S10KLrtaV89fYyvxO24GDh1zo+UqvrDXT+Et56SbYlfwhtyJEWlcTOcQ+j7+os0+KyWgkCw272A9
XSwpY5Z/jAeq+yqGZo1SbTXCa7mLK2u16Iv199QVE+hPNST5BhLWOiozfxJisa18YpjNP/HDVi3H
LOTiAcofg9aYv8tBU14SST8Ttd2YF4whOdWOb+kEdnveTr0WAOi/Dq80gnT5UN1L5R/8YGFpC+ZD
X+vGgJIatpdtxPzVSVwWD7CV+y2K1lFRfpB/CCVRVbzhtJHCDCRrPPqxcCnJUBX50PmN5C2uak3W
mCWFEzvolfJAQgKXYQvjIeXbSNxP42msZizOtnv4Uq1lk1epoTqTrRkCOGnymltYQqeVArb0k8nf
o7aVbX5mwne/rsr1eMW5NbE1vaFMHuSr7CLEOCIZitTgEepNOMCuej0+NkqlMWwXo3xDFEsN6Ily
cKVbr8iDY/aEYUJDZfoY710mneKmZmxK27bHhUCl4YO0LUYCBqWGiOJ65pFWey5Lv9QKKhebH4Ug
/16dPwovolHnpf410Yxb22jcwgPgHGgyIB1ad+Vd4ZIZ5Vw6M8oriQbuv4/3TOnH2b+5tjGx3Jcc
vwJ8FlWNQNWvF549/r+wZCYj9OTE+aVXh3iFLCkuyJWtLBAKZxzMnXMPWwqL4gbX83MjqXn+qhkL
2H3tza7cu0idSSg2nl42spCIYMerFuYpR8CDNM0jpS9pypKCXfcJca6L+EGtUZCFN0l80f+Tthe8
+T9823m7Y0Ldf+sHI7y/+RzfVATGc/VYH/B5IA9vkddgQ2zqKNdiEsALHHV4b/GcW9JkuE9kupWM
HcrQfmCsm8oysYNWnJfycg4FHmTpdWkRGltgrbdaTvinJY0C0BRsTIVXb611OjgR5ZywBUX+sfOc
JDSILWwK0FxTr4UbFKT4WyggJmqzR6l5OwfNFoSO5/oxP4XcMbS0n+W4PRW3gTWgyPV7Z+YFM+w7
rVf+7tU0Io3Mbyx1mjG+Kie/ozTSPcueMzh0PfR8F0De3kaBkzD/SAR4izJ3ljWbBwhE+L3NTmah
lvl+PFDYpqe9XaGrBEKGz2hLDcsqgRPugO4Vb76kcVy/VteIObSQw65UQXthkXkXXeqrnH8mSH0n
yvE3CWyhhGZe5kQRJdeGDzOnmx/VFluEMiQcPbS8POVl1XfPhn4IK3yHgpsUVPEnYdOjyWhNq11k
1hcTZ7/XXqJVy8Y0WY19tyAwbUNpYS25+e6vuql3+v2VPce1Pdf5g6Y/Li5DBFe/HFky4sM5q3Oa
k/SHUCyiZ5qbD73+NkeNR0FYkC4KmyaIKdF3G2Mb0HC02yL5FEF7uKKGU9psWlUAVX2vvkq6hAbM
4doIkzbJWQ/rawUqzkm8I0ycXNXx2xWj++BJTRScpECr1v297eYSeEj+Z++TXzUUQr3f3PGO66Do
WD+mopcG3L/rxMV12l2/e+1+hAyLR0ymzhDyJcBeMJXzGv+l4aAoEsraN3z25So/d8HA75mmsPtP
ry8+cMWPZh/0SiZDZuqbrWn8J/ObzBCWG7CNdEC5yb0EjJMaweZvJgMSBxPXn8tChdPwnXdmJGlX
gvnrbX65PZBmykL90YrLf3WvlKFpqQdOaXl7fU5MVFlt1KtZo8Pl+9I/6BZ9pFQhVoqspcXoHq45
9g+9LDX6UA/1Ku1I/VVVuoeyUv9DwBp6FVxtEv76IMRav8o9te0X2iH2l8K40YZmhBXYH4LPCoQh
L1HD7PCM8YcNM0VG8F/egvfkjCXeHLIElYTAwO8rTQK21bAzK4UWPbh1fxotC0p3Yf5o232aRbLg
amLJsq3Ce7uW5yQHER0ALQyMv9rbaBnHKqPdbnsKZH2LQiUVywdJP0hBYWlsI3xhVDtIWbGsxGhe
CCIri1KtLGP0kvFdso3cnghCtaFViW2YXs89QC6NMWo2MwlgdPUvo0/9Ks3POisOD9wn1lOQpBsU
MaXYAro64xWY/eneLPrnH4sNVOwCX3lLnXmzUu4sl2JxjIWkJnwgx7z9lOzikPbmaGY3UMkamK1E
HQcofvi141cXIxlRs5E8s3/dci4gPmMgaO/v7ZJ+MT/xco04EYMrF5yUeQHJrMJsauDMRBmhxvmW
PQZbuMEf3BjX8CAdxRKytGK8D07A7Ble/Ks0K1K2+M+5VJHJaopkl4puDn9P1zkGs/WdrINjjzVk
o/giFnQoVN0S4BBqaHfUmYz7NKiGS4kaiOkqk4r8l7nL0r5fS2Pwys1G1oDdkoG078opAgyXhPP4
uVgRjb/zPVOLcshgElfxywlQh/HJf/+2ZXWlcRi9OoNbXW6xo45j7j/q3OsEDzVwxw4LFdPLHBTM
L+dZHieH8smO+PgMBRbh2hpMEs/XYP7vfN2hwESqFp3m/YV8hqVr6OgP1zBryCwKVibrnLGn0nzs
G7PexeAv0RR/0J+YVOXIegluZOqSAOhkEU1D+OirIFceJGG0YmLyL3P22HmdqWeLB51/QJZR8I+4
0TDya5prq44DBlMTj2lPT7Xu2SqCiYsfILwCksNaJ1OwqhS6U3Eq9aTm+65pbHpW+Yh7O8epN+2i
uTa4O90teazZV/uQ9mU6rsKfzikOLDxJdJ6+rA1Sp9zfvbhLethmH90nYDnwfIxuVZfPLBR3ty2j
Xe9En9DG0dYc2bx5ElEj3PY/wzAkFk1SRUGnkE/tk5gVJvNnhU3gjGefwwvXP7BdYuqW3oddrGhI
nBA4cfn9cpg9oy1xShsyq25DpPyPHgy9U8iwdHEP5JGnOag5LK7pVtVjEkl2srB/cxe7p+37zJlv
vghBPYWZXjLy/KVC9xQdJ1YdHwxbTwZWybpn9kEf1m3di5CBnqxsMW62YYO3FCmcEvLA8YkmWecT
PwQZDgtxr9WNiXOc40+yyZH0tovs0k8ajWPoDitgCVUwhR25W1R95Kj5RBJkJkP+q6kl6HGNQrkN
qZDZfEWGVhxQhL/BkPrJNPkgX2TWrbAti1t1tPV2yYfBozmDcSOxpnz53JPTSZBPrg0y47r/jOlE
8dc/ApRNP8dLtwQym9BPHTB9fvc6wr0/AhokKpZh6tsomLQxmIj7YkCOBwXR0qIqXeAGbCY+Adt4
O9ASf7YiqvaiuGPcJXSsFeF3vDxjGMSs3juxaM61AsYakLNRuqeU9yikRpRJNwXyn7QB5lRC2nBi
X+CEiK7BdGCbpLfjLVAImaI6OSMpOt03fhVY0Xhl4Wp+lH7MJN1bXpGML4xh4AG97Wu2FvTJslFG
5LDhmT2bPZ4VNmbbfvXS29Z1bYbBXpQplMv6knFJmgoPVHg/QuqDup4s5I2uhOQhH3oj5veaLu+d
WuajgG1eNekK7EnzjizRySpc7M/YbRnNkxc82Qe0Jbc+rpCppZbzW0R26uCQt6HhktWyBsAQE4k1
wgTwz9bYVc3u4y7MVq4zumN7r9IeBYdykotYiOBxCFe37HPiRlK5r5UT849LHl40SGXd8esK9jWg
hqh0BxIvB14QdbFhNsteSUTYktvdOZFf0ACxLxp8YgO+7aDTexF9iFFLvHhIPIUVZN151d7lYfXw
dQ9wdGaN6O0bmxwvEfrOYR3+pddXGsvDXMLqltVFD8a7v3aJqidAzkQiCWLw/UlC2G0sfjA0o0zf
Y43tkAO4w9Ex7ADyfWWmUtAzRK9Wy+f5DjDiLb4OKXdCdXl+Xfkxd0WRB9sQYiKfaqV6kTyIl9aQ
Ymss6tY2SG00N8+39VHppPehucrXFqcWHczKkfu3QiXLqrjVT4rFJEmubBH0NquuMtXUL3h0jCbL
QcMtjzOwW4lAHyMM77wuxDdgnG7YTW97XUqCuvDDfdHwtHqPfFQPotH+wAEqOcRnbYQUNTGA5QP7
84CRzlQYmeaUNv1qHDsJtXt1JNB8tboL5xfvE8sj8ZBlXMUqBoJJGKxJmND3itbsH4iQJidr3Gsy
mSt2EU02MRIVByISfrvmVXSUdIIStqZLExF1VNwrLiYgjfdmbdv6g+gBlnrkE2cGu9C9LJnJVTVS
fWhVxf4UY2bUonzp5VB7fT8nNH+i140T+iIZ/urXwbq/L/7ytRpqKR/ShVoj35v+jYMVen5r2jAW
sXirC4gv4jhSZB/a9VuHT70dn/GP4YQaLIYtwmT6jr2z2ixLqJRWBWrj35tN3Dw9LJr467iYuMk6
9udAWwO7ReJj0prDkMyLAT2dV6JloY7G67juWe1rl4/0prJCR+hy7biFimjptUbBsqwUIxF32CxD
cFgCtqHkkdJJWyRTVlmHGzYko8m78CX+od9IniiIqda2JJRGHfuY8c/keur5DfXTaGPRv6UgTxmg
yzius3WivJ8SXkWkyH4DfmEaDgPFcPmLUW1jRw911HiYlCm+7+u1rdl8JkSpYNBYVxIOGNm1C7QI
Zcx96c/60FUGVt5YhbOdvfI0guRlRJAhhOLXCIvrdASwoXidP/5MzcTl95N6zqUoGJXci+HOu79v
+1RlEfV7zrM5DIbS87QYCBG6c9TbNqRfTjB8lc2s4ydwJ8v+RWzShjXDoaCtfqHi724adOMuejde
dcYcE4XfuZS2FAXxONawpdx10BYNfXAcPPyXlSF8f/jNZrWOazRZZAeZ7h5bMvDFr4k9sEviQ0Q2
u5CgBHZNpcT4s+Q+nrql7SEgaemVj8RKlpW+ps8Cy0hW0BEjOVHYS01jRgyICwDsR+22Dr2bvFFu
ITZUjVjIf/hiAJvlgQLuau9c5n2KGedcy51cgoPkcXvTAxtkZ3l2kPtdf31O7tU70v4Lvj1r04RB
8b+eCZXCqOzJ4djQeGhJzA5TPg4wikkCbT9suhtp2Lv1Lo8FkN6rnyS+HjvumP/GUBCAk6Fdb47f
PRslKJF2MxO2y+eo/HRzl3Z9ds1fimsOAUY/deBLodfzbALyI/NB21t7jdKBX+iGZkAN5CD8wKsT
mIEuZrh22qq14ih7XRinMBfAIK5L3kxiwk+hwJI8FLktr72eZ5o7xhDYPx9r1C3LwU1VPFzQVEY6
OBjXX3GPrbZgEdS4sXVDrvnB7qsPl3dGcL//StvHFAjyQyq6NZgXy9ujPaFu0Aq/HCeiXF2kcCqo
M8vZlTNwoWlgJHeTchKCbqckTzy80jiyyu+gKtHRNU3NaA41P47+lcfjOaNGdXWBHuxnFO1d1dEz
J6bRXhGfcabvWrOpAbhOLGAC8Acu2VjvlXGZz6Axngvpm8ZqC+tUYpUmboFkTKsgVpzhIVVUs0Np
6oPwmceGM7fSljcH1YfKiUZtsnHFokjymcJtReMJl4WCZXb1R395YMSQN7PdqmyR/3WDVok7BzbA
hKZ+Iy9f3sFuCRWes+2eilUHbUmeuvKD3IM6mGgSpxp4GAWuVEkDZVXk2KY7f6f2lZ6NxKAB+kLu
A978fM5DZrSwoxyH9+bAWuXdNik+QO+rrfKqDT2CKPLn0AJfXBxVkETLjj7awnRS+NefhhMlD8wZ
7gzixIsClCz30CzP5sx3YJDi85LNl8R3vwJ3ioSYZczPDKpDe0qjZNynYh6Osm9lVegZan0gwPhv
Sj7jZJMQ6muGR+CP4enIEvbWP685Qt6m+M3GByQM/CuD/TNk4U+2eqVdTkHhHatu7XRx/W4h+IKV
nXELW2Tw2O3ZmbglUbZFIcuoh01eRXFbkR9T/OFuSgSLkg2PrnFhHZgWurx3fsAAuswaDWx68Anz
LztiL2QVINiswVOMkyQ5TX80xbYZviIrsN5zLLCEcfyY8l8ZH4H3kfgTLCk3N8Hd8XNKiv8gZaZ7
WCzbrSdFm0oY+bhOsaNyhHY1HI8HkDyjvAyoQ2jjqdzwDaXNNkB25sqWmm1/RzEj5l+R68FJYf23
HNgFUJWDPh3rW0PFTRx1LYrGbVVL6Lvr535SBmHpkCQUzdZA3gS36O0YTIzHKPEUKewiXEddVj8u
lt1gDaN2H4dCIFlT3QvIbcHd+273HeSbOa3TYFT/eOr6I/gH1BIYIUDfNSuBlQcBZdVXbLqylSNG
pZ/jIK+vCSmNcc9uZJ7B3MGt4z2vgwG4//qMNmzD+Izmh4QO194gmDacIIfM51k7glmYIwpRRNE7
kxcmvKc4dkauq83AD8QzKgje54Qos1XqNsx3N3UlVX1XEhnZMhSjE1NOZxbUPNSxkVMy+yUeHfXV
Cc1WpKEdOEFyeLGpPaqIM+haFn1W/im3xEdp412hPYdOH31Rm90gGAd7FZ+8Q9WEUXUn3QsB/Yuk
EpH7eO21xKgzLjcblpUxJsSFcKLB2B71uzVJal5LduHkVMJJmK/StqAmmwRud1KTKdKQ88I46Ipc
Dqx0EKmbIWDWbwp4zurvU5hhymM1yXMnuk37LNUtc/aKIKmtYTJ5NiwWfO88jcZ4UK9EekYNbj1y
HWd/f8bNG2S/LZzTkK3Nnt85g6PHfOIRBICBwb+i+IlCzp4GGNfy171NZ5M7kf5XboSL5MewxPdz
VsTRX2z9v3Y1Se+/JBbWbXE/hRm1rmoDnKvZop0IrAxkDwmfQ6qL6+epuF1RAthgD5GzFPCg2ZP6
1IVUkk8rkyktE6EDLFjC2sFPM+b0TadS/okToY1CZgxR0gm+7/IpHhjuwygL17rjrBnwvJqUwEv5
z1o3KHFOfPZ6oormhRvDS8kFot4Frp8mOoy5M5sVc0HYKdDKWwhaTW99fKwE21kPnjztZENRSHrl
REipjT4JvKXvbXHuRyAjwkb9HlKgXKy8ATJmFe4n6/ZPYYnIeRFSPv2oECLpnR7ge3w6yvlpBmqR
CJbcB/8ncV/AzDzWPDDrde9lLQfO/KxIPMsDSQ6XHv35ZnieXGn5ZPFquG/UYCceklaGudwpefz3
kDwDVDQhCbNnWU/EWGDvfBhKfg4qwcR9jgi6jw/jcuYy8yqodhbSa/j9XDiu+2eX/kzzVb6X9SVA
RFwTYuoKw0bPb/Uhncy2K+YWiTfjD48SEj4I3ILf8o9tj3T1LDNrjYqffYIKo/gKtWoNuxHNf3TS
I/lqRS0jlnkV0fqP7WDRY3z/+I+fdaqCqqkfcx035W+lqxvVOetn1GgthmmA/btuw01WoWkdV1Xe
VRIw2wIlbUON0H3X6gqL4ODAiW5RTWj2g4I8cO86aXWJzeprZzNmBuB+Q9adGKzeLYHDeggHy5Bj
2imLGHNrzgJrXOVEsDYJ9pTfskNgrifxNp1sJmSchbtRhmyBGTfAxdLup2B6DC6/vkxtdgiGeatN
jqI9nsazoRWPH6YMd35ZSxEh7skXMfZnCc4en1Dx99Bof4Wqmq9plCq1sb3aCzgx6SLR6MkOYFKP
e7C3r60rdL7L15Nrz6REXfkOd2UBYCMskWFipy+r8IPbOFI/iUPjazXC272CSIJWXFZQ+MvRfYvB
3hmwcl2UVbUPfYPT/zS74z88bK4dsjbgCE9S5gHRuvVje0KfgIUirH45AEUrTx6+ZdNh4mZBLXHG
8rl2XgxfwXbtlKzhh1MXHELBkf4bYSsQ8NB38GTeStmCbD28aR/zEgJSIHZhZIU56ICWQhqAq0Xj
vbrFEKSJSuGGiCVAfPzWAQZUj5I/+RS+DvMultgTsG2QeP8I2ESp4V949SK0gCARb0pSFZi6LD4c
AjPUcrTZfWxPDbzZcXffYeEuqTzM7ewMSWUR5beg0lhS8O+uOH7IOROfwy4cj7UNIczT+FBd0VMb
dzXVu2JMnDWXdaY9vC2OniQoTZlXaClOBsXN11e4VV85FyV8ftGQXX3PXpdfzWAluLPdo/2ShJFC
OdkECMnrZonbx9ygCGPIIQXbvaLxGnRfsdSbkCGLQAxRuTaWJy98LhWSUKpKn2R3+FoQ9Fev/pNm
F7YwCmtQFZIvo0cY1F/bgIDnGOdzLGO/roxYqDkAv5+OkTnBeU2APWgL6kUbw1vC4IJkLPoC0pUD
IS3zAxaAY2oKe5P6YNQgdghDX5DUyk7+80wyw+P8/PeOZdzA5S/WH5zKOHmDAyBxiFWU2Uffkwz5
dbaF+Si381f6qPJWYbkeiP+4LqOA/NL5k7gj359dsKKeCpPartD1LLLC2gcm88mIdhDQh7FYlbE4
mEraZuhEYsLYGQjUkeTE+jmDeMuHW7s1SjC2XqzrtE5HH8STXqJ3yJO+praBptINlrMNJ1ih7cuv
TYZVr3aJWiYyMYgqjhs8EevXyPlF6j2EVJ9fhWYUlGZQcEKW7qLJ6Ns71HwVvxWwnEoLqArTXR14
+cYewDMUca6VEhMyXIo2zSs9Sj+7JL/KGxkpEOtUwLHRKkHCPar/okUjmaIwbOE1VhJ/XXVcgn+K
Kbd9zJwxHD+/Z19WNRBq6zIuFxzBZY/KgzxrULfVo9BgCMpH5PYBsOtR8WmKmF3zAKT+9tRWLKkA
yu6rdUyFw0/QdB1bPHS6ClK8W7xpnatdwu5YBahUXSLE5nrKpm3LZLaq5mQXKx3/yRkvCHr0IvJX
9qRztuRtPZe35w/nh1AODDCb/f/D2TiFXd0tU8eiJfMhHJUISZN68xMdKavWw+qMuAYza+L2V0NC
oBZ2wWpSuvHG3f1TUIGP6FJdhnJ1WIdpGKuzYhLWtP67TUqpYWThjtW78G8UtLy6De5BhUeDszSn
RJIn4ChPQJLxwQ3jMmpDxai9s9XuCjzKgzbIXECklNV0/k53Q1R64Y8tCCDxlmA6AJSAMDZUlXxq
s9Qzs1/WsCGmQc+DJy91uc8OojhOnvlxkmewumrZKRezRvrVYiAi94Vza7JFnmEQeLFI1lZEG3ft
Z1LnliJgUV+Vb7c4GL8YMGTX9yu5xg5pBOleRJDsRyrHvpaR0qf67kQIoBSn+qGuUyT1cT96bPm0
Q8rrJ8tjIqy18qinVAC5wHeT190RfMrQLLzGaTlh+cGm8JgsxDjLGNylLOX6TFh+oAT4v1S6eBzJ
1p1Pl+e0kvHmV0uGABJzQPxTwExm4n6Sgs80pg2Xz77nyPZSsbVLDE5LRZKLYtX87oAryfhTLb62
Wn8SYZ5Qc/FJMXYZWrV35ftJQZAeL0LVY13edcHTF+D1DxQvVmafU/en8ebrhVdHIfjRZnILIAMb
Ks8g/eVUhgo4fyG1fySGICUFb0prw8N4hg0unCSHpZsCE4FSNgoheQcSc+vKuBqr4aeD/vUsyUqT
lWNq0F0OX7ENgp6Nt8DyNVFmUKt5BXVgAgVIkOu0SxCHAfQ/G3+ZjCzP7h5gqxMsQiDnnxrF21hv
yhtlPPQyZo5V3rg5TYmjKhexIQ0aIAEKBbSaIRI6/E8d92bKCqB13Z+KwoaWpZOUjB0mVYPMWE7I
nAM2cazLOtzvJUGpruA2YTW6L/hOxlfklb9zsZaO/jmGBBzBt2hBwOJGhi2eUFCfHj/JR0/MvmeP
y3VKIFEkXSOtE5qDHpWz/cFHJ1zHO1zqMbn3MYwCw/EmZRH+dcvd6zWbtMFT7rpzTszfU/ufjXxP
+ZMBGxG2n3GQX6zTm06aX+WDWGgyahsqlyo7ABZTjsR8tIaDMqziHNqpTXn4UlHIMLK+XoKICJeN
jOTf2LUp/gB4Mj2KKtAUIoMCD/pmS227v1SWNVhCJG0hwUlPMJ5Y8PUrqU2FTn+hd7gjCOtsFJc6
EZJz8rdgy35RGrpZM0ILVORdgAHHZdedCQJgMkPgkFL5MUVb+kVPPCTDJUv5HLXH3QIL4arhP+M/
f/jf7fdwUgNPVf9JwMmXkENII5cHWcFPuHu84lsoNdEvMti2vY6cnd+hyoiQiT2DUhIH2DkM1jFm
+eomBqtbvRWUW/38BEt6xzesUh8oNayQhEiXpSs9gfYB82cgpdx6fOzgylsPv1tyU8IJ8eAlbsOw
vcvqe2RDej3k4tOaD1O5QjLk1hBlXzMWP1FX0Xr+kNkt4rtewR0L7G5PYdZEI9e4LMyiv2xdDGvN
BwBBbuUYqiZ5fvj6QMUIyuiF0j9AU90YIGH6732x8WJ7q5SUa/KLU68tOaC4WPCTIIQrCOOxtnRr
yJpS0iu+s1jlH97H5GlBgnYZztdSsZU/8r2f2cwVEKn/dlTNIG5zBGNn8MXrph1Zd6uFYyp5/zU4
98QQWHyxpPX8r+rDMch7nKub28+uGe8uHvsyMVnZ7eeyyWRrj8ZKUixZozq5J3j8d2eKOaFhJNfa
5e7j16fEVYYnAkVoZlmy2Y16NkrJVW5ZmRrZK+q2mFTOD9SmGHaQ+biKeMn80Bj2uVdra0aiExmn
0ztGE0eGhGu9ifGn5eTcSvaftvrxMFuLehjwCHa7GbI6k2VEkW65+1x6Drcrk9JcpV1qr1Yx6pyM
J6lsGBaykID7t0F3/ZeBrlvssIHAeGoYgo+0KoeAokX5YQ4APFHf1ujFG581Pox4irJ7LTDC/8yu
MOvMSnjLkOmukyRAyDiXiCzxzkE6eVQpkftGyv9EIzVmqCw6TGAwpQaA653AFveM0a1LsHFMQHku
IEy8vEZNJOQ0ny/WsEIplALDU67MdY39HY9fQHMDB+spRjpZxGduyp3o48+5PUGqsf4RdWR7E6Gi
UoFZlMJBn1HAvlyc3oJrxg3tUYEosvznaxsoIBfUjz6kaMAqh/i2sIFIouOg2WQyqIlXZWhLXVye
GNv6QW1zsk16e6ik5O+XUTZ0PNfC8+LrQiw1oUlg9cZpSJGW0ruoNifUoGveZt7RtNZf2PEYBJFS
apuEJs6m8ZWYC0VICsCS03MsS8RW61d6DOBADD/QCqlUDVGSqLz2WWhx/P+96Xyh+oAM7hj7x0eb
f5k3ohgIUvcSYyQfZK92pNGdxI0dtLt8agYbtvKxmL0EtxaTAOuY5jYe3hFOp8OsFqcjpoSTJ0J3
qWDmIEVu7lg4CzF+jMoW546C9VVOzwjpKawkxXTY46BeN5aPt/pRgzRp+dfhwlYtVlLoHJCHevSm
uksFH6rvTwTvySDFndKuSokH3Wb06KEIZJOyG20glfAg7yccy6HzHQqywbZpQZRn+z9NiuQ+UWvA
LIOM06E0gpSH58EQQikKxDlgbpZethrY/Ietul5L0b6kA3E9ucEof8swoiaABP4LDYP6UijtQDNI
iiU5KrI4c7HUQAwTlPVbUq0g+2vROAQ4pIgy3Ngz840wUiIaasmtxsODbNGvn2SAUJQxFOloNw05
g+Aa7JsrtoSamn03n8RLlgzD+K7qP6w1jng0QnlyEtJ9pzzP2TCarOStXM/FmKmc9xFCXiWzk26c
VgUjZTUWhAwP2CZZRxWQUg0NVhOppWWtmr2I2/NZBZarw52gbpd3Bu20peosGvUGZVkApo54GkPS
WB71ur1DiEWEk8OntH1vcindZLSf+MpEsaVXEGER2ia9nyQMQfSLQ+fQxN+TmkAMhdD3p+6rNWkJ
eXnYr6zZ8rlbte7Lg6eOD2kr0RdjxmLhi/bZtrdMHq+chaAmUzzJa4Y23VGmcZ80zsAe88R0vC4a
zBU1oEYmzo1YeZ4pXRRABQRgVGV4xRu6F8xwYNC3pw+1Ifzh6xEvISoWvokGknzJRNlgXuXEnbY7
iYt/jSazm0c5c8rn7jQY7MN8Kxw7Cm+PGJKFRoBo+C4x82WpaqmzEFyse28RMjUfIdLXygwrXEcD
CSUYaA9yIBdLKCmACCnRdi8aRmGpYWKTSJWFNNdiFtGthObqhiGl94UXhmeEz2TIsCr2SaEVqkeO
L77yWfjNckaTjAoup1JlwZP2fnMqIRh29IsFQ08fZQJ66dylhbys+zuE0El6k7IM3Hjd0QQuuYC3
HjwD31cb0wj+tkaC+c/dpRkBOoMqFioLhCpJJqrbUAKtqD8T500mDR/FQzFVvsKoa0unVzZFy1C8
7W4PldLtrayPbofeNQ31nWtr3UBUHm4kBCbqbI6dxgx9a18wkXE+WBZ8wLaZYCAJy4kgbTO8N9RT
es31qQUWgGHJ6YlOuMUVcILdWQ0E88TPqhxAKZwzTSh1Zc7MyZplTEmE6MkwpYdq98DJBEo7MeAK
cfqdblsb3f3XzwzoWcqxj68BYhfTlhJAReovzSHyiqnNQEe/ZLJb9occaNL6BrJFFpEAHG/Lr6FG
qITglGVb3kRg5yh+2Na4DTSFXk48wMi9BidB+YSSO0k+FX+eKLg9bog46smxLlfu/ZqopaZ3u0eW
/Z1LNi6yvi1tcNXQmFgfCKXG8tyFatygmbB7PZRLzFow6Ng4rxmTspbdBoFAFrbDytZkhi7EuGFi
qkFNT39+4X8NwGQuYoq689dAvHOkGrHr8idlWV3q+SVfGuiyW/pQpINJkQ7IYZd3sITNqarJnELu
h01uH5Qc4ZES8PaDWdKJFlgTqQvjNRZ1l8eGZ9/D1juUBMF3GEdNyJOn3K5gwJJt1XQZfQRsTDQZ
tjfNWH+Y8M5dzV1jsWZ7ozZL3i3RkJyi4dQR7D8ddACVTrgyF6TUHcmOTWeUEB3lZ/vrzYGy40Fc
I7qIYNnX0v/9Wa89+V17VlWol9WQn3h8H4VQuMZrh9OrFPeFsVPV+hWR5VJs1RTyu89x7JSOD8xq
9IaqTejRsQVtOVRHGFMBRdAkRH6pfHkGdYzTS52QPg2111Kwumzg6BmqoxWXR0oFKNHHKEKEMj91
RyaRBtFHqbiNmYYeY8ziEnRVvZ9+mkjru2E+R0brhCHn9NpAL5wfCXNPxL0bSesgqgjtp0+lHbv3
iARxC01jBP0iNLkHBGFFm2X8STgoIVU73GoVj5+XSPLH2a+dHSfS5fLOp2WXSeC05mxTp99PYyRr
6nk4TDiAzpJih31Hf276lRrhs3WPnT+099SiqLRwp3h8mPA2aSqHrf7jm1fgoM1oklnjedRegGFI
05iHqksqSIDCplCsqQdgvW99K2GJ70hHw4acESNtVf8dwt+X1D/2CF6CvJx1w30sthCQPuE9/bMt
GZfgjnpSkrosLrkY2GCjBUdXkbafal4XkcY42DRAN7lJGyJ4icgveVW4Dxibcn/baBEvGM7yGUeY
DHK0+6IDnMeCpFzKnFnwuA8RqgpXMc16omZzoLC2JHgCg/xblyuwwR87ujoc+CISgkCdVoZHlLrc
jxcrqeklz6BhTICjrMWYdLG/vkT6ej3SDKz3sBBA6ioA66gIeTREys6eQTBH6evzbO9cGlKn1+Vf
TAGX7/xgsnlFnlSSGbtp1u+Doj5wQ9ze6CEYyQfCcED41N1sk752/ao/fhVGXcqw7tuukwpOWHue
rCtP8fTxuqZvcCSVDgWL9KdXXY3UTdJqlDZ/pf9dgVDuuPZ0Nf79LoEBsHxHKzhC1FxzrKKOOp6C
ifR7bF7a3horCNuSwmsMadKRySP1QbQTgWnf9d+nSn+SYlQ6TM34+3TGw2wqGH6efukF3IhtsV9y
7YRG1coZ1BxNKspQl/cKEpIoUIMYEfk3JvjLZTXOjcZQ8aGewHLkpu/U/PoGpHLUw7voypZFrhHm
7E1mj2dKBy406lyNwioJa5/8aJupO1MMF+TqfApOUGIaxLHOfqbuDRFJGY6rIJHI38f8aCI9of2+
1uhzUsb7bEN2PmQgoq1XikbW69F+MIP+5XLQSK2nDazc063o1Uu0Rr6roJAB6xa1+B2otmuMMuwz
5GT7XRI9Pn/3udWop4xP4VA+hpTG053AUcxSeR3YWe/JWIEymawWRF2yXxCU7hB+UtWQJlASBW1E
ovV5rNN8SQRV1JJkNDiGAzNOBTbw71kYxMKyTWzPPwDxLVjm9N7YmUDEv1TQ7hAxY6e6aQPQFkRU
ShE5Mgu1tkOYynxTC4zxVBp46R4W18gN6qY7iCFwkJitfyt4AMuPH7KPW8G8HMSL6ofe6QybUIHB
M0yGdHi51e7h8K9MIG5FSE3O2m66gj+Ath7iolJs+ar71l1pp4O560u5mu2REImMrcpAtwJ7IIva
+n4ehn4ONBMQkkRD43xWUeuB3iC3ZJAZ50R/0s7myVRbmucfXJnFaGibywhmtW5lZdXaquY+fAWz
/KG1DpYDbDosg86KdoJKSjk5s96cb1nxAn1BEe4jedPakoAqxIDZrHcmPMj1If1PLnB9cOduXPEw
5a7E/Pufym0GCn9fAgmGOhBZV4H95+0iDqC2cRxSt+C/ioA5h7twyHIFDJp0cSU4A2LuAK83qyv3
mn9Je7MTRfawRx5eObRx9GVVfJH1/iK4Hr7yC/KbVN5vAaaKP3vGpp+ddyiQFK1NHOE/cG41taVv
D6KZEUt0DvTTDyi9m2dkw3wRiMqDZ5m/FRiReuAGp5mjIPSMpcVA3EcMxI8hxacMDzOY9SX48DFl
+dSGrsbY5Uy9LAkDgNpDvWA2hFGDXVVKf3x9k2PpS+Xir+sruT/8HMYs0IA9T0u9+WEset4wnyqg
mJ2tTOabe8PcIGbnLBxjyuQeFfLSHmTsgFHHbfYUmYJRBrABcxVjKuVr4R4aCdj0pJ06TD1cAK3s
BHWgjdpSfNXGzM5gzSFPnNxjR3h+td/hAcWcrofzqqd7g6CnQajr49RG9WBGbyowHUCs0aFxH1b6
1CPXYWq+jAROw/wvl7HzisjDQUCLeTeT59adVcND2rIQf3Bh7lBy2sGwRiET6s3pMuuicjHE1hzO
8s4rlX2FKfgSqg/b12HJMtQBoMq/Mk5onClq2dMBD9/zFO/NjBDt1zyT9vgUqeP2o4kpIFIe5bfs
MmDjGsPO2/vg//FrJzOTszvGOgzZsnxM81Larb6CqD1u7jzkH9Sp1vbMmTdW+lm1h0mu54EvrIFJ
lYmp4LGeXHzIsFqlnWPdLvD8lPKOCDK282HchoSSDGXaNoYuPWvNWluincGFxIiSAD8trdUAk1qa
lsgE4UYlsDgofZz6eImzS9jIDppxcjyKNNj4cWIttcJsUVB4ztuiFkhVbSBt5y9e6GgT27YsJ6Zg
m4TkrsVVW8uxIHI0758cMK7EdKre2Tps1WM3Vo17SeAYD6GOnWOXpAFS3cEodfBA+Lp6OlPV5mKV
hhW17X2G4cxzBuDSX2tKx9Rb5jXRD1WNFmHrxb+DwzHqZD/ydDW660RPJ6xTDkaVdG+nFWrHwWdV
/RCn+zbS9NjQaF8jlUMNuSzt93AwNhZLsWimOH8hSGcnHVcQpHzwesWogkFHZJF9ooCESNVo1Y9W
5y8ZRliGDaScALpykANOw+JhNLZiE4hVuI9qN+oVVuvuiUBGZSyFG3F75Ac1bCZKyRfoNa2Kq7dG
OqoHjOoxb8QAiIElzcUGLDjHXc8GBi0O7u1/x7EoXEp6pcU+L/+3b+aLZ4bDx1DzhKUh8swk11hV
EXjek7q4fCWJhHvsxEZJNUzD0OxmCyTyaWvuBG5IrTaPI/t4m3dbZ5T9MRgK1tC8crbNYXkB7rGN
K8C3qebs+KUZ6de3sfsmqQ5ese0kuacOW3ZKh4xabMA8UY9KsTtGKVTD99s/K5qJMRR7Dyl8skap
+UIcTLRxBPUkX8THZ1TXr/Ttz2xbgL4TpCXv1hZE6Ky20j5G+cn8TqnRiL697tbEqepqs6V/kYZZ
GyO2LK/0gAyV8r3XJ9AnIjY0yblWWUg6jj6VM5hmsOXTMEYv5rZu0DCg6bxyZiFu/iidG62tj85b
NHbsex5c+9V7lxwHXe1tEbL4VPrdFVFASsB377u4sGXnwTPhOISn/nt65znAcWn7AvcdvoH4tYJz
YiO2aFaO3L55Qo5r1XcdIJ0duSw7qb8BOtaLsUNeDOzD/3oUhnwcwVcdorXa/2ujVlBNfobQfR1S
Dd2Ex1ePXlFMxsf+gtyOGeU9j5bMZVLiCRmoQU8v5BISe7UA7+j5Zk5Qut4FmGVe325vrg01Z4M3
zGRpd9ccUJw03034i7LYgVnFYCtHGuX5SJ+lyVaeFXgVxPdjTcVnUtcjHxN/NxlFCHqqOUZX8Aiq
fPNfF0KVCWebUHUgSV9VSW9DboAlF2gdjVn7H7QBLhOOqCVWLSVXXX3O76ORj5rJQPf4ADXP3q9w
U2BAp0DYXvvzJBSldaadUdMFt/air08nMoFQBiW2lluk9k0gMfysSSfH1dcySQacN9i8WlzXrpKF
gQ5iUpVTFC4zCOPcU4/C0jn7MQDftuTl6svUEq+03Y8HqxX5hzqM3RH0xYIoyT/A6n3ioJhawDsV
TCslKoCzsZ7RZavzUcNDY6gaXibd8iKy/2SxpuZixP3+9XMA1IrNUUXYEyJ2PibAAqS0mZY+cUBf
vOHaRJyVfsH2Xb+TawQJsnlun8o1bjXevh+kaP9gBaXwEw5Kf6jhAKIRUBRgLgx3Gb3l4389BzEu
mrl8N3XkQ3BVr5ypajaWKFoxISKC8KblmapYZP/dwqPBQqfdY3uzQi1+7lNvBcK2xKeAVF0UOYb3
Yzrw65Ehs+PCM2yL+zqgvqSRjumXih0NuBkLGW5mTW91x/CBhpUuFaEOI/Jhq8V7ZpDiv2pN73FI
Yk6auruU3nnSCgJetCRGKEJjzRB4RCYdsgTwsKeJPPlWXvL01npuVNy57e9gdrRZqAjbpprM7Svp
cW+tqKBd3yA/yYRWdD1TnrOvUxsT3wMwIrCDsR1MoO5jcrfo7O184eqLgMKQ16EiHqwhglPY3HhJ
thpTs2RtyNwuDF6ojCAA4TzOklGRTK56+bnSZCqfijRMeZ96FfSj0tTiC8JxWYrcOC24kCcGXF0U
uITrCLtz6JHZGT5S5XONTX48kE6DdmMW0QmDgHmoIWHpNiLZsNkZIpVZ92UxtrS5OaniokhZOin4
HDNnczwXzM7s3uqyjBHxg2dgTxcwNazLyQbx/EgTmTcevv43X4lvUytnPnrtBP/tgJy4sCef1vpm
rENyCgVMBo+BqZIIxVfEQCXC8bY3HU8t41pNm4xlXma9TurRCjlgYQ9Uzd2tKRyuvzpTmCvpUT7T
yUuxHmiuqCHtBq43AIQZ1WU6p8ZNij0DEeRB7RkcyGX/56tw5frcnBKVHjHoHH2iRzA+1XOXaHyL
2ryLGemmriADTjSxTt6C3RjN+h+wwjYP/xShYBtfAzJfPmzUUKkp1sQbR/qE/md1w+xzuPSkDiqy
QlHlNLhaDNjgNGYCd1LnBvTdpork4vnxHHOKTQld7M+HOe0l2U6oPVaJIbnv+KVcQ++i8elFNSIT
JPAHgTRgwIAu59dO+mN+eWUGRVlHqc6QVvlglPXmcF8AHAbGbEYRPGVvFrh685uBRQBGZJRmp2OB
ww4q53BOK85/FvcV7Bryf45BA77T5GILcdIUv5HlwV/9SuLKrIVnZaJde86IyeCRP6JXlALy2p3N
hL3wCf64tmZ1o+Vg1aYaBSPzJDNvyE1cKBVt8K+40zvOJrdi96uu5LZGXXi6I7lkdnh1l0+M3fCP
ufaaV6KY0G7hoXgzE5bXgV936hfB+6D0BoaNLN42aE48GXCFlGTBn71OGj2/UMYKL4z3Cih0l5dJ
G/dRID/YLw3LmXEt852lBdU+EBTR73vStbDxYtAJUMdaaEpgLwXBJxErJo4BSkIvfprQ0LNs9XTx
vU914JYjW+M5wzWhn0K3nHVAFRN9jCIV2lIcqF8I0lCnvTfC8+A4uY2INXbCIoWDyfcrHLcfvIHg
eeA8oUE4Vly6dvj65JuoYN/MB5RZGGXFhGINEvSCJ3j74ugK2mWVrs7xbmObOXQ3A+paz8KRCepA
j1jmaLvaLfbAiNyZNU5f64gWBUcJwgT2j//QOs+uf941IbTrYqTrSR/PldiT3tkn8WYPRRzWbkyy
DjVbVU8X7XId3KYg/1XNhHJbGWjqKVUAR1dXj6HNs59qQcXsvHxjjCCexvaSSOZPlCsSZ9xSnpCE
LVU+R6IpAY6H/1GrtbeyPQDgBY3xVxl0G9/l1Q4LbtdJHYiTT0UbbVOjq2OSGMESd7qWkUzes2qC
iicvs0ITfUQgq+OwuceRuuUks9ejOMHxc3mkyGWZapQVQtCWkwxXbZioGlicJp178lT16yy5QO9Z
wLz/06bxAK1xfdypxHugCK6mLsTQ2ESNkvlszha/ygBCbmpSox39GijsKmonyt0NOKDUxMnMnEdU
C8OEKwX1HEBgz2wr2tRMWjRQnAPptHWuzZQxUfW7C01PRVHp/wHqOq/CUvfxyHe0goUzL/pFKPD2
qL/7rCgPl0FVnt1FohbI/AeRId+0h5vRENGKMSd7P0tRYMZdk0ewQ1AMZnnUuxLL2Owg+TDcL9L7
9shuwPcMDz04/Hx5/Yu+RzZlHpdale4R6lAg85RtTWG8TjJVYRVrOstEQahKuBafcnYktqa4MocG
LaZ0h6n7BmoMjsLXmIDJZycN2AL4ihSpX6rpnoTlIFPzk3y9FLQVrI8reNon0CtMLYF7HEqNTqQL
30h48h0Qe01ErhKp2WQi7jFz8eRmX9h9oodWBdD49MmkztYInL2S36XrwaaWXjVvBzWsteYmaujG
PM0GURMOQD5IwmNvvgOT4rasmd8OrbfdhU78Lggz8IZR6YL5AT06m8sKJKQntHthUXM8uu7wKFMA
raKuRrsPqTVg0PfhDcuBd38/+8sqvFyBuk/uld22HFoFVeIeBBIdpV8OPn05rz29L8Roq84hRMeN
EDB3CyXqzMTA9WVLgoRBffUsFE5foqq4mi21T3GEbOBdm+BrzfSP9SbPyLzg7pvITa0erwtjd7sI
VTkw9bp8zwTM2916mRHgHB1yFeAGUj2O2zStjaqgFRfFz4o4aACzbDCATC2iZOGdFXLMG7TnoGeb
gznnKddgmMK6bfHCQnjIKc88sfyDJv+pEPunOspEELo9bYDA8QEwGLu7ZGzA87GxIKIfAC4asaVc
xs537hXJdTbo60iaFbL+MCtk5ljoAlXx3vugirece6/vQ63mJDJWrEPPEq60VEDBSfyZkFFqP1pm
dNHAooq22TJx25vvqcVZXH5UdIh8tXfibHPC6azfxL/vLOTzgol15C6R7tkO4Sr3xJV935L4oEkz
0CKDS9W74CBX1du5xGfFRKQvGgLbQp6xNXioF3CZRIBeykhpl3HMEg82B7kiKZrnoOBo0+127NeJ
9QCDo7gwdZkjGn1gVkuJLVBkiVo7NNXbAq9owdTOLkECNRhPOG7fIZkgVeh21qx9NUdsehN4frWx
uNp/7aWLDcr7TSkGMQVbERvwxm6tgm7O5SLudL7pQbzTT6DGe7nhG1cHCzQvFadXajYRl9+9peN7
U2ttefe9MNEMJXQfnJQpN9jpWprVmBFcky6ao0jIwSljzNK3arUtyxZ0dT8buAtrEporS4QEpm1c
UAxFfkvljfEaIxWoJbGwHJg1mH/K6tuMHLZnLFUtv6P+35E2hG7SPSBwGIoH7hhASyQ3SJ4GZlyA
oxhf8Y2+pUvNFJRFhI18twZ/oanw/2r1M/aWAZ8eOo9M2xbSgYB7j8ybnZoFjbYOaWjQro11CmFb
VY13ZTyvlPpwYlDeV8zPlLGkP9Fv7DcnQK6oF4kmuv8p4GngPulMyZo8gdqPXqyiwg+JlisQ2WKy
jkWb5remiQJQtG7s/syKYfA7WDH18wKkkRLMUF4xEFGHhKKCCllDnAhhaHw5HGTFS0oWEDSm0P/0
NI1FRGNruG75ycndDw0xWrGOlpovsoJZm54nKyPO2jbe6G6Rz8Kme9U2BDyQJMwKcRyNBkRaUwTf
kRbZDO2LyCjJIRqgC13iqXDQ86e8LAJzYVqUvzw4zteErk2dsHzZ3+oEjQiViYu8voG+o4yceCci
hj9zeshAyDNTlf1TaCh+ZyYm0s9wiM+jCT3wY5k8567OWy9BWSGvWk/6Eb/6657RwahsrTp2IgWo
fl6M7PPqG81iS6odNtSHzNs6nF008vtqnIDkK0XkOvtQGfCCMjdtGFn22xKO0qtVfJpMlL2OjI2x
hnosV3zGAH5CI6I1l1vl9Bh/gsDJtxO0WFXTYesJcYxULSZKUbCn70wPc8DMyG7E/Z/iNVjBojtM
Q1TINizCzkwHMd7w6ZFlrQgB5M2oGCdu+qqk2MDKw2z43zKTQJcI8MGgz3KCRqyRPlUo7ijv7foa
QcHGMfoFfFyUgM9wOqRsxWCu37bh/3VP3u8kxgkT1fRHLEHPUQZHdV9NaqDckvRGG/iD30MV/FOn
6Z9Biw/0v+P2kIpDa/2pvrV/R88MPQrf72o/aiGfRjR4XNUhYV2b4WSRJwtLW6hmVkXPWJKTjPSI
zxwQzCBGYxVBOo529aWKAsuZW0mC0a1pOsoWv/jXm1OW1X5RybEDGoIPcsGI5K0gFWTZp/FIUCl9
q2w6t1IXpXfa9CWAA70z67SDhl/5/O3exNpqLVH0ccvBiipL0/6cPzbvz1qkK9CoIyAAiJjytJUv
xgvxiADClN+gjgh3+ExdXGck5Qy/kf3wix4ftrAWnI241Q61sMtVFzGQMwis5MBTd/jISDR2+JJv
xfxzxdWcC8eM0fR4sS0kWKF3/6rJyD/Fyy+ytygwQ7guMOQKQips5c4U+sJe2F10VMm2H8K/t7Xa
8TB2gwImCUdoD96KUYzVVN9AX2RgCfGS3bhulv91q2u8HvnW52TZuVlaWNS6HBJbnFdeEP3aIZ5q
mu85tdvfjXNxImH4o9TYXRzPO+UZmhc+hCb9GSihB6EQ8QxxbmxfZSlw7dJLkroPIVjS1uhVmFYL
fCZIz2m/txx5UQs+YF/6QduoRhnyd5NCP9Mj+s/68BGo3GbaJm7xYzVpFC/WS838nqAdXuCOy49n
fCuIDb4FOgV4MEE7Wscu0CeMd3/QZK/8sVo2XhgGI5klpJvZgxp5Gs/Y+rblmrWW0zPdjHda7h/n
2NF+nLmhwPdMU9aDL6RQjpUYHBeYuUi0bHhJoYxT7fzw/tZtohQm/ftU6XvgHHsU6MuTMjQzxEp4
wpOO8goGdP4cNffHvib+w9dfYyPWusFvxMQHDVg3TmiL8cLyXOJvm0Ok4LWuEwQqLwLCDSVXM3b0
G/j6Qwx8JkM34H1eCxbpL3r4eNJsuagRuew5KfyRZmgKyD6RkToH0NZvFlaTp2uAHTcwx8t0Xw42
2Z/NXHMgTRxYyFrdN0bMcDeMV7wXFAf8EflOt6wGEqkZR6wv0ugJ++r33av1m6qFzAZzL8RhDlHj
/W81JWUt4WlEPr1pqDdtOk+faDo/oHBTvgNPbbKl2P1dlOmuLm7U2k/LYAuMJPkAEiTrDZ/ecf2S
t0UfYqgBtPM5g+TMI7erwwooZBQHyHKTDHsm4CfeVV5xoqFpGQm2JzyTMdOUizNDP5OW0HaaOHwc
NKv+QCradDY2nbtYsNYw9oKXc4Pbhw1eCPRy98kjt5akNGBH7zUKgfGeeF+7o10zxqEcUP3jAhSC
DO/dHGQMhqNFZ/ECr/TFFHyJ4RnPLH0LlhGxgnNqDwgKMg0+obzWyr4fnO61qiH5cSGgMVa2vvYa
gtJiM9lGoLd4C47A32IWOnekAh9qPpGeu1k/rRL1WrDlutUxp0F4uOHKn4+RtnUe/KDoPrObTn80
TEe5gRcBo1wtsY/lPYsvnpdKZybEdM4DStidlE3jkru6cBSMW/aITKIs5tiroZz+GHUOg1bbcbU9
eGPifxoqzGWENI8uqyP4oGb8pYrfL6u7Q4h7Oo4t6UJIo3FLNXpkcrCZ9y/S/l2L9yiZuRC3/s9z
h3DHUaSUmQdg0txOvaGIifNeJfSTopeGNO06z4NT2NNaYLLHy8nOV/L+dZVRzm74CeEKuZG2oCiJ
uIxdBbz+tDW5haO0NK1mqjuKDBJzyW4jkLl+G3LZkXJ8Yz1iWCIRpjEXfmWEEO0eie67jZB1c6W1
onW1gXGRNKD5n2f1YiyN4Hrs45EUyVfb/Aw/saS9vfdQ/wphmvPhdWP++Ru8pPmU7Y+I3ySYk6m7
PTQiG2W1Jz0EEVhl1fxPJNMoohT0dQHHkAfiAQ/Y3ATp6beh6rrf+sEB8XHWFcw+D0jiqX8zz+CY
/bf7bGfLSrj6zKj+Z0BMTOQ3rjztBwKtgqbVcHQ9HA/XUdfcaTOjRV09x3qzVHdqNz4UXEUT9V0j
4Ulqj29YPI42IwRejfrpEKQrumm9H0t+F/ESaIOBoLAFSGUI54SbF+EEpR7+tFwDqKHHISrzKtVy
QXiqKJx9njaxY44FdMGOGzL6gO0PIgRgd3U1Blx8XXKKtioQK7a0KP5crUv7xn+DuUabsphbtZC9
s1WpEnkAiP2fRZSKJUiKswwn/oCHjJ1vYSRPr+vrzM8xf+zy1ctNGDBwgHjzGRJqXROX2qV/L7z1
QA4vW9YR2zIpCt3PAFDiUslgNBn+2r96IQ9HeRAxZ/UHYZ4MwKoegMew3Xv56UstXlYVFtjrZA2u
2jscrZC9lRDFsU5SAUgps4IiW4MEtwgaaiYb9dEjO8Oz9rIHdsa1HxSnKL0iOgumtP+636D4Ba6z
IJz8OK3dWwBcv9m1q8p7HeD+no9NTYu+SgI7eI/drGlKGeeXLBcOZftHt/BM1d5gCQrTssnKWdg9
Cca0xzCELY6cZsECAkHZLcNd69M8r6qMq9WUfpdnbQXovreIXF83XYM+f19pS0OGkqEZ3LLxJ8sn
BQHObw/F3FJMT/POuopfVKfgnON4O1/6g8RHuAonTFYgu7ypbABQXh9SivT4cb6yhBFwZiekGx+h
qm2p50ZJUc5URK/ZRwCZ6aI713+YkM5kExUIu3kMu8r86z48V9G2xPoUn9RwoZhv4nJyaVbLUlwT
eE2Z5fF9AVRzicgRrJzNboUtFVLdXQvPBUbUj1VcE7RBBZuFmiTKOpKmEkPVb1dg+NBRSC6GnSO/
ieUYPColzmTfJ68mHOb7kotpyV7ZI7QboPC3QKH0Y0LU+MBG9jh9E8wXxSNg5auaXS4aRLC3ANrU
pFDbp2073MkX1cWkT5vL67Tyms7DbMK5h80qRLkplYp7BvjRqhhwFWCa62tmt5SgttTUrcEN6/sp
/QT6vKfNcc1LUGYMxA5Mehdo1nw3SOIQLrWaORpstZoR44kmjM8GUruDciGBNN6W2+HehJy6puT6
Y7Oev+1KqRiRjIshDgGLMlmH0w/gl5sotK5oDhOcssX2ZPAxma9VzZ1CLBrmaJumaVdI8EyP3/uf
OZZfV4L9c9GPfc12ATR3T/fzAYKLRTU/Xo32vHqhnzqJDpWOEPHyopyPaDKRlfCds8TjJqHVQ6YI
E5dts9yvKg1v5rclIeUE2aLuxkMAf8ZswqXED6eSoZDEZYozQF7Ptgtqkc3ipi3IqlNAN4VOqyTy
uXUIW6q3I4Q/9dZbO9LkL5Q2RLUFZ18nNbzCyBPmGIb9LNrMBHO/gnAhafAd2x5F0/tqYfPi1or7
so1MyXUInxhAPC0LB5SCrlVAEuC90cxkeYUwSf3xj58jmG2XNAaYGIF00OCWySQX1a49YAePQQgF
uzKXrH6Jp9GPyQhuctXsTeeOWI44m6AbVm8xYtNs1/0pHqdZ/NNM8l44tinqu7VdiqLeFljXU1WP
mqbfPj9NPz8z5ZyDtecPPiJdIqFKWFX8HqEhYhHo9iYPqpqWQ88KY1+X3HUkAAwQibMIlwEKD0Mx
oPuDwB/n7K4J8b9TwBTL3JeMlwjOkG0kfp6PqYloRmwUkgGTfgTEuXEqugtD5Pt6ARj+H3XXsLFf
5ZGx9lOzKUrCt4/KP+8CuJcoa3HVAyrNL8OCFss2OtQWnoNwRCk0AneLGkBddsjVpjsXhEmCdoSB
KN0HTjoKLwAHbdtf+TZIU7fWa6vNOgH6pj7C/ZSfBPHNQp+ew7iLGwkO4lYLJ4PHkgXE678XWha5
9KGz8VwsPrpgHY2Nl0am3c3NpUWPmjXtM1/86UxQfFrx2s/3SSOl78diQkbUC5tpZuUWZ4TvdG/B
ScC7PiB/nLI2ll8e7OAu2VWsdUUwjQuRrag72XQWNS/F5WEab/wVtHpI210S+A/Ph0GsGDApDxqY
aBlL2AoOlRioH8t3Cr8zi3KDArVEjajExOBDjge+aRuhArAV9+/qMbtJQbKVJRxtwdm82EN5vi3o
uYh8rWNli37OoZk/+tDDAITiugi4j7O/s4zZT8NadvnDFHI3zhUavoYd5r6W/qv82tWIw4HTXxN1
HrP50hllvVT2xjMNXqtFrNgjX6olCp7y4gfti8SIP4o+nUPz52OApis/kU6Piz2im3XFclXOkCpB
uj61Pa7VgnlvaqRSCIukW+tHBmBgRSwEz9ntW0+7MjlAQWq9SUT2Fhp25B4VzHdzzoeYEBKKbjQ8
FCoAEvbK28zE3NYh0ak+4mHWT85rdaT98CD/hAKvJdGF/+hrAzM++Mbpm2Utn2Tmtt6g1nGVRN/0
tWX4kgUF3EYHUp5pRCjD56EeHPalngvyppiqrpa9i/cIZyftYpKooVN1t346jcaJM+bagfgrmjUP
lnLf8NDYCnzl9JjmhETTVXS8vlKjqLH8eUHlh2omtkwT9owPShihF1IJwI7Fgq64vTnNEVWkyics
dhhfLE4q7qCtXW88aTVUsu0fP6cao7OLdZFJRMbZaCw/4oztAeKjVQvrvzne/7fT0UB25J6cVZu6
AvvxSVLDKyZTvoIyFeJLgkT3RYisl5axU/RPfG0MknNWtjqJamG5/UU+anCYZh5Iiagj44/9+q8D
kwVKka1Czo2iKyFgK3ahEw11C6PzLaK6nz9OeWQeMI+GgaNlDByjOy5+JnKfIWDLdj8FTRya7+o6
TizXL+48257zwLANClXyswpjA0V+jDJbtIv+sPybbGBZSfdTfaT+cfbgibaleXiusSZfrh7gfwxr
Sf+Gw6U1/d3cugDm2jwVmnlxVF8PpofaAXCb/K2zmOdV03jwqNjMBbmfS5SBDlmp1zQBX3qZAkSf
MjYaeM4wLZV0wjSwebOwWP0ZeuxUwkoSPOdpmADonm0UUEsg7Q/FUDQuGsAULs/saueqkAMpZdjy
DSZmHzQgbmM/dJVFNGOSlUrlTpIE0mQoTpTJHi1U/VpZjvkU+Yiy48xLkVNHUoNxQPtl/RjLfTqR
3xqCqrCRmdjvkNGQnJD/jQQswMRt4hIkg92ls4ZzqYYgAq36zzzakmVe2dw9dIyRKn8gC1CsjjW0
ulrYlJZqASYZoRSSzqfwrMipDu0NhbDmARTn/HaZxS4cYidHBAch+qaqYZrl5TBIgAInkZygQdmH
a7XuQUywy6SWhAP4omP+Oki+crdrKD7BMZ2iJ+godOCWk+WK1IlpwWjaLF8mghHZuQA95jfaEvHO
9pR64xz2al5nNcCtMXfveY0bNzsSQ0+JIoaA1dmquoiQuQy1xdqnClnX2KnFBfvvlEGccwnF7PGK
46LFh/Qt2uLnbnSAcUXAKDdF6OAKWq/7bRpN7DDWwy2dKWe0lRNeDP50erwZvQkVyo6mbpfSQFPL
Ug5F4/Lgtotp0WfrnnSkttgH1drQWP+BNkLqe6UHOAplTYWyswxKUmKT9PoygJEKyHfR7ANpDEsm
J/Zh9fh4d4fQInfioPd7LbHXj2QQsOWz+GPLQlHxJSy9MYRNpV4SlLpwhd4kmmwjYqtSbfN/s7zp
F81UAk/OzGRjA+IKogjcae/W9qSdoqQhk5sEQPxm/Rx5oYgZLF4hZZHivZHGb/Yvb1t3THIYzbtP
mLMHNfwrlBR1WU/PY8z4UNTDvpD/EcB5joEJQ+uMMltCBWM0xTnoeEeUp7sgn874J7HbrJdeoB7g
k49ULGYo49G/OaOVNlDOiUBPuVCo6YYTDvP2Ev6NAzJJlrirMrafK8bOcK+MrP7hhCFsb0LzJ5kG
LdOtmakvmu5V4VA8UBMjmiOjSAXLuxEjE79E/BTsjsoGAghzk+JTqHQVlZZxc9QYChLMGhLQDXSg
OByyjEvJ2TYzcmBpg03MbfE2GbdR4Llq1eI6hXbtLbCD+UK4abD4Hj4IDzFX53PKPbEBtoPQ7eUV
PB/0cTy5qzH+DQ/1TBIom83zinyWwXgB9b1S6cxuP1hX179ypJfmFjKNMAs32vkLh1O6cQEZeyMw
Z0hppaKD5lBhu+MZa54laIPHWyosiT1HfzIcSQgelBHsOhuEJBvPKu6QxGl7sTOLOYi/uPpuYIRl
OJ6G7ZwK+cFXoOHj2MgsGW4HL/EXNVOlcvWiD2WijyqKomXRgrDbxGipoQ3497m++jmBpUDF/R51
aWIlodDjlzZWbaCg5CXe97TwoXnuIw+4yewtJPwmKFhwoIi86Sge12LUKo1ROBOnhQ2wl6hU3tzZ
a5enD2Uy5nxYgwpiOMqc7CUJUhTGBWMUn80YM1T7pLaUZcM1SA6/tMBe43D9lvtfwRfBlge2p1gp
odeM806uEFLkykuw1xjDFSmV2Kd44mq1wOZvZxKyQ5YsozU/94xyWuIgfml/zpbokRndE88olHPC
LbAVaGYih837iX9D4C8EwgBAbVX/C6m/E/1zMP41OjEjisNOWzkeUYkHl7msFg4Tnn3yIi93IEuW
iJtxjbZ6uBOok3BmC2WbwsgZ/L9gfGogZjGvS7AhpnmnzRUBIhs8cRRt3hoHSI7IolTpvWiQ/BVR
BOmbVaNqVApNDWNvVT9fe0wTvHEGhWZQq0r8AOIfyRGq7+cLRu2kH10mqwCHWdDSO9Z0Jp4fvQqn
S7LBamOxp/76GgwpqOVimZJuQENBR9M8kAZ+KPxhId7L+3lJqWiaXNJCxHO1OieCLsMFUNnSPyfo
+0mSmk5+jdhvrDg6OAKSgvtY89+i7zA8tnXiASjNGMJsC1Gr6nM060AGqM8Dv5vTFt2EQhqGfqMc
IYV37xSGskqEG3N6EZ+BnF5yPzTq3gRiB29Z2YPYW7/QRx40ekuSSZIG+nAYCtK9NCJwmcTbTz1F
E05MK4crV512KCs/RcY6OwNg0XB5gvuWkI6gZ8ZxSowfvcOhbnT938NxsgWsoZqE5claUYZ4+A20
OQ1ttTS8wqW0YOc65ibwq7yf11wY91JoQn9txYGMZa2K/RbI5Pn2L3HjrXbctIfWq3KHhZZ5ikXM
0hwRfij4wmS+qZr4gb49Sg9SwlgQQEQWfj9t50YkwNAvvNW27rtSf0kHQCWCCP97gCDDvP4nzPJC
H1ztwTDN0PZQBTLjlPaMO8RCsV+/2Euu8yqskYv73owTdINqyqXcbQXCX+tHYlJUF1uUWm2Fwc0v
6M4QLJ/99k1BtG4oBKKxcoOxIZje+U4Tr1IsI+y/Woe0FwVRCRvqK5/wtYt5iBaNs+HuJjTP5GZf
vGEMYt1bdI8JAwxg5lmulw+XKyP7yqWoLYHQxmGGQrwNo4AV6/f/BYyfaW6mRS/VRVDv038196mW
x/92+IR2lIc2hOd/drzq30H+JKZUDzeWVXYvzlF9Rqte2Ch0NEZWUAXwj2mXfwRg0rnaNSj+VFZ6
lQoKG0Q8BPDo5ibN60LDcoW4OwQsW4nJJBaob9Zp15da4QyX6gSRfMrlMdLybbRud2VydqiwGnAF
UvBNql/WBfKrdR2J5ao95nLSrMYvlTZ1PXKYPWYVhEa/9feuqk2K4nHgePS+Mth4E8leNIt78+NZ
Zv0HyJmaVQaCLLg4iSisjC7u0h5OViazxBNG0tr3Nh1H4CzXmeDCIcgap05bsKGIZ/2Z29Zxlyjb
jZsReI/Exb7IYVYjtd/zwLA8vL5YqxrRyl9cs31BCJs943bLw4TwF3mlPtSn4QNvBEvk2XohjkL/
SbaBpsBi0HjPvYjERz4zHNT4/MjklpM+dYOXjXkwXqyQjaq4UsiI1kemJw8yQ+AUOHhyEj7qZrF0
sDldmAUcLDutsqa9eh0SN089MyKwWoZe4/2Z1iqRkjSV2MnEaNF9+T7PgJcZfNLXEd8tnQPQvZEL
OCU3oJKviT5rLGWTifFKgkBKTK3WJlxcapxZQq0lHWJIxoB14scV1uM0dGyla3PhYlhacau7uXNg
FamOkSiNnq3FA28D9wMW+R9LjrrS232s9s0Rxu7JXJUXu5o7d3sew66gBg40OAeYeVKzPyIoUZfx
mmpKw1+1ZpJ7s0ryD2rPHdhcBkIsP0HlCuu80jmKLoSfaSA9SsjCLTCl7ZiwKl9JsJUboPwi7w2n
5ntTufDBl+OF71KfXy8Bu0gZBgzBQQ6+DhJr8G4JcxaN/FxHNIoOTrZ6LyD0esUt1sgvdVOefuZJ
jNmhf+zqbWbd1hkPDN7hQJtO5mpRjz8fDc3hzpeE5tloMRkpUohP/6tbyARMKKcwFWObbvjZhp5Z
pKwbRNG280V1VV18uYDfdbMbcO/vazgisLUqJrkCPoHACZjSY7dr/1k/gOTNO00GBCf53Xg3bxl0
SzNNIEjtrqo/i2sZ/pk2CRzl35ne02YeG8mHnAlpLC17zMVNAwVtzs4d+9c+8asBL/PSho0dRjJ8
xm1MGjwVgxVF5c56mugINoPW0caeYSO85jna3EoGUbwWaI5CBZWHT084fQcVAuwydGzvoFrh3+Oc
XXHKGnsDMqSLfjiZabZxVT3vCTNti1Zofg8C/xTUqIhj6V4ZmZBmhKZr212VQTXPMR5ldly7k3xH
Ub9lg69QhteZzCVhoxh3r4YvEIcNjDO+qkvxDXIx6jJxLBoCbM/OZTWa2YxPiPdX4uVF4BdZxvqr
oPEcRKcCowzVDyke0NiDOeKrQ0hxWiR7hbMUnD678chSa9G5NEL9gMzT+mp2Gc/JExJOevulE/VC
lBvXwAUHhc5Jm9WBW7Zzr6kRVIwf+KXGsN2qCqC2o5ed4QG8MsWh5Tj7AecT7qCChji1IlHl944F
ouVP6oOpk9rB6pOHEg6XJmnLtZqnR9QipvG8XFJbAq6j/LDUudOZzCh+wC5auH64bkHkN1vUr+9Q
DIGirIdDn0rk62yXxTd1qH+czFLuNSSIKi5wxgXqhmi/F496y1C3KiBdAxCSK8J2PcXzdpCFVIIu
XAJbMOG7VcAPjcztpPpnh4LnTOfp4FMokCnBsshb4kwq5eeF9qyEWzbs7UuVWgnLHU7TZSe2MZIi
CUy8t6dh5d7PXlH53jjRJnW3Dsxvkj1+CtCu1ca4HBti2lD9y+lUOC0uF0xdJOSXJgoKF9Brzln0
u42y0NymPKRKLe2tq3CYdx6fR7Zz+vYDp5wWtPMeAcg6dYzAgCrCCkKM6oLHEGsh8qtr98K+xraq
MSEPOyRr9lUICTYXLwphw8p6/lmlsedwiYGvz0vJPN2of89PymN4vDkbuMpox8j7xlzWJjmrOKwT
PsgSummX90llDxE1vNWXwLsRrXBnOFgFeqbQ+F2CaZk6PH4RUDgNGkPhNUm5pEX1yMhvtcS8TNTx
AxQ0anuLPTYosKWffLYinyRDN8UN+H/A2vYsh+hr1KvAKNtG82X28491QAQ0TVff2lvPczJqEjvl
HlnbjXXbFkeC0YwZ3mniMe8M0zdciD1ocEzltFDcip4PA8Li/GjINbnvL8H5Ekzi2HPdLbbpD1SA
uV8Q52OywyJRhzKOhyFhOIbFAuTZyxnoqatUzv/XicfLpQZnS6fdMs1RSu2dF7e5ndyA6O7uAIZM
2SiVlQHkSJfHJsSbxvEvhEvt5C+nlGG0Wq4RWZfZ8vCRYkpgo9Fp2q5I154XC1CUdCkOHuXKZmLM
Uph5tm7SYVIuvBvpFQVkiJyh8vVjKHKOFw5WZUKAlnLuX2DGuQjBMcP5U/Yuld02ITXDAK2DrViR
YwzZFeZw6IUjc1V8tv/oXA+i93YU3BIiOqrRqzQjezD4iTLrCbemsmyZJYlFlQwMxnbUlcrzHtdE
01CsMdf2TXnVCJkVv1vgmBrBbhO0K5Pt6ihJ6jhmQYm8GKJ/Q1qy3hPpZg43K8IU86F8yhAA63G3
YACwGd1hgfgYfWd8UUpXFBDAOa+exss+j0SoXbya2D4EejmQS6pYmD0U46YVPak5qYnijFEMxOvN
rOPFt+5USM55QeQYxj2EeMKRXus09ii/jWBYXXSwJdqmy6V6n7uJhFyXD269RFso6x7K7sez4TRj
WX1uA76YN/JkRLmj+iQFIF3Gzfa/TEC6L6RZ/IJXJ7E1w8Ydm8CMiXB0DAs6UMMcOwIWZkKC6cz0
qd7RKpXaiaoiKSzfvbGB+lgWrOgP+A+s17HooP4Sgv4cFrlsmaEdE4IHC0qjicfVwyh4ehIIFUJo
z9HJdChbC2p+yzs0Jfso8UXxmo8trMKu0bjaoHpqL0eY6d+dBlo2kwtDB4CURfeFOzY87UOHXNKW
PxAVWStjQ+aL6pyYLP1AfDBIIbSR5XwciPvMtZTkr5WO0O2yZK7p8Z9zUUyHNqI1tH0JIa1BzPdc
rTGtJf/0xNWfRKh9TK4nk3tm+VponcxCSkH3LvfXwVYIBYLjvmZPAmniajMuA/Pbho7ef3mlfegO
xMxNloQx229HRfIrC8kd4y3LEJlXfppGrt0cjQKRe2HwWO5U4XylDiqLjpZt2wRtj74ZYfrb6QaS
grS04Tydi507Oaf8+1nNs8zsUhdpfrVMpfqtDj0m0Ny2LLkAGidEJGUej8xfC+ADJWJAs2xUHi/V
p3bIeR5dI5wRios76zSv+ZTYfizm7bCbaI7N1Gw22PtaIRUaHhfdEex5d+/wX2jlIo8TwBimFP0Z
TNQgfHwzRnx8ejQ3750Y2cTu1KT1hX9t6Al2wqqIoJ2snWqE1gp4ZJFXcblrCwPwSXjCiCFEpzM1
Agz14y8Jg4f8nu0DVCrJPPhc2PdP+XaV3yMEEWVFoMCBs4L+Zel6QCRtzRMos9BwV+XmGc/i9LKV
ope95oDVBwUatvx1oSvznI/wEFOeCNYIgbKzbm63DmDZmnzMo8BDkC2jpXM6qnOeruWs7wq5WIq7
OEcTUfKMva7xwpiJq7NaPFpNJDN/wFa9s8OJ9sGShDh/bY7Ms0lhwAtQL7NcbKaViT6tnTAVbio2
UqmD84afz1p23CXSrdJoq/rwA0zcymcDmtSMYnk49Z7pjvMJXRMhmqwO2ynZ0TxSLUyb5OafVwuu
JOzsPxPkkp2l1PqTViVosSPayMvSKiRyUF1UcidY6zIS/aL3vYGl63JBXU0vnrZroCvQIbD6G2my
WMcRnZjmSFr6IiGaokYV+DBYmrl6aHbMRI7VW/G28iCP/8Mmvq4D5AFVlRPvAuHK17mHNN1/rBHs
AZZhFKiFXnwTQQCX1N7V7jp2H22vQKdySlnmHiw+IWKknW74SppzZ9SROdMnzkd0jvGG7jvEGxB8
QCAvV0lDOcO1fe99F6UETPT1Tg84YOdiMB4R6YlYXmeYcRuPHS0tH5LTkAgdko+vZkzPG19wsjlF
K5TiqkSl8TnvAJBjuiXE8WOIKm8EXKfT4UigTVB8mt2gtmr5kDiKGykNevPJRy07nhn0tsCWr+YA
9yN2Pvk+jpeQdKe4fPhQRvBUcjxUtHJVAVkbWCKLDme2wkUknK0aUZ6itsUfBhWby9zxcoNlhw8m
ffGT9BCcW+iBuExkHb7OdLDYNJqlWq94ueq5SIOCd+Bkl8l5Zb9OF/wPqcy7nL4U7GecNc7awrRD
Djj+3OFqNPu41lFW8MzOR0doAKKDCmh26G+aUiq51SVtmlhJedDnT8PvOVOfO0h8Td+xyQJenSWr
t5vR6yF/GSB59xdI0Hphmb9M0TE7nJrRnWhvdtvVrkdOf48XP8xyaN9pfbL5joeH9ZtJCPxd3TkQ
FG+eKxLsBXKfjlY620CUmP+wottBqjUQarrWroMVaCjVbOHiFdP8sa5Lmo7HJFIOu5joZ1oMTNbe
fDaHSiFOf0wnQ5FO05dKhK1OuQPZsQ/xeTe9/ttmQnncGKURqiLhEEO3kQvuzeblzLDugXRV7LeX
vBu5l7B5IEwAxBSiOvbDDzzxcD8H7V2w+qQ2lJNMzMTNb1fH++M3LTMcQranT0nSwJwE/ShVoHl2
WTbiNIIN5NH0GtH8uqGaDHgBhQWQ8RGiFH2fogn9yZGMt7wuF55OSPnwBNi6UraB99uVpd2aX+9C
nVeVE9zNYeSIWFi2lR/60nzRm6XEQyqnFgJrOZD3d7GJxMc8A2BB4q6ME0xJGIJWN00B/O2oOCbH
kPI5XdyBB4F9apI1ldXvuDKcf0BextVweJLjCvw6ZLVldj9Y/+Dzw5sePCCPYSNeUqNHc0M7ksBv
fJCrLDFYAyHgqIXxKLjhs7E4VE+ldXIAFUuSMqytpGUJcb19a/Cl4U2dgmRjUZfz0LhzfYkrHI1R
bypd0EhNOBg1wZAcEYKq6aGJxnBrLUiyPNskt5DSsyqD9RNHUOEHGqIyEQftq6H+kcgJOB4SJWeK
/dH3OtAicYDecvtGjh0eRNmUM23PNrj06OIVQwKl6akpEki7e1+SpBcWUzCF4+PUtaRbUv5d5Lwh
r1v1WWqWBg0hWuzjvB6wBcdR0S6ngc6s0/OhNY2GkVk4zuvsuQAoWk+6ca+v/6F+8nV9TMB/FDxK
zgeEaS+EZgI7OrvXzgPlSCh+/HH8sZhqVfQ5eX6lhsGAiR0OIkqKDkA6A+Jzhk5hGxyXsJ5M0kye
voO4pJv5xcLOehmKSfqRRaxCsvYyPR/Fm03RqsrCKTyMc3stbqgyNih1zYl4q9m9Y/MlGM5PJ3lc
2fQRUl51BFQdXRZK+9im0Fw+Li23E6QNzCgT/NQNkT8SBQ+AsjFF3sViv+TCYokm7NYkP6y3+6mH
pEeop2ol5f+ASTnsc+4jbov9J4B25Y5WFxJoz6BL6SjuhHX/VgHM8kNmoLoc35FNQNg5XGV/zNJv
EiwOm0075XGPQ38l3Am+BNdteq1R2ktSSWfJbKgP0Z9VawVaBY4UbsEiWfDXjiHfpzKPgoOXKRnW
yD09GawHX7zuvL52dQq1KNNZBgALiqKmiNb6n1l+QQl4m5tUJ4kAodxK0OvRQvRMsfNBA7fzbzbd
VTuPXyOnwAUf3Tw7PgCSSt3Do47twDhr6pVqeVeISAdHXHXT6mar8E4R6tvvI0TyoedZRdECKigB
FGapAJrFiMd68suZpQDUmA/XhUBrn9hYnUup53E6Zk7vFg9muPxGGL+M2wib+GEnfjd4qGCgIbVJ
4dntfQnQOOGJmi7b9sXevqdkrci8P/DvyZ1Qn9ndCgZpTgYPMUu9UViUecmn1gp1rcP5KQ737O9s
yox6fm+ox6TTexfnoaHalRTdNBPFZbBpFJ7cB/KJCetfn9sNHHs6iXABoyAmeEDZCfu+H4njJGAV
yeNfC8MYZazNSTuYQ3LfLO14SFDTq/Q8yqm1/NYcRpRyL566BAeFkQ5/X1KF/mAkVuEBZ6E3RH+j
BTVItZSmd2LJ+zwlx7Oh8X6ctKfq2a2InxLgnYzciS4nvbFQj2qfxZfOAyj3xha/z1m4hZNV9tmJ
Qg+hBSbiwwqL92+9YPHMWzqKVQzZWSH4wUvIc44QDzAl+3vJfYZ5RS2KVkB7pm48WENCRdtJ6MRL
YeITiU0X+D2ZHene1nlJv5hvBYKnxZLO2qKWGiyGDtRadhqJ+Tn38XxxphKpfkFvWT2jypsnD7/T
uNbBffiEOQBM74Wj7JNhu13sElC5cn1Wi94qmQdVu1Cl9ZjwckUIsU+suasFkxUxPCFI0tObonxc
Merk9CrEGhQtzVxwYc4BweqI7fsPINVyK8dsv5wKeHuVmRdyjH2ZgZ7fxaCcv6Dm5W7cjV9u5jPX
J2FoBzzVlvyFdYF4L6PSUT1vRuD/QeWYXm+v2KGbq6UVfAzCn0/jvA5sB15YOrSmjbowTybiSi/7
i9Z7LuTtksrBrZplNVJWFqQL/d2CoRLjJO0uCTJ8W1JArVzTDmyI5KwXxQ0ooMWoxI7Nx+PEPpdG
0Fb13jew0xZMMAzTY7WsmNubKG2lgYejHI7sfpgV7S6JDZyc1GdYBVqQhKSZYq+T0GaETaFGmeO3
xr1Hm2Np7Ak2r0W80yKHeG3IO+a+k4gdzrpIZmSgyJsiehpG5YLTdFEKFqQg6gnAwPvJ5Zsc2hgW
Lbcv8ZsOLc/6oqSNMzykvvTz1xOyiHCPQ4GnjZSrAxNFXrh9U5/u5w+3tTTMbEL/sLwX5tew9FVN
87adiYbeP9znzlNpx0CcoJRYQybdEUoXz/KaPq889opNIuNgzkLv52ZvxqQUvCP8zIH2sOK8vemx
5zZTuXgqW5D6n+BJ168xg+6XBDV/mMA/xTxqwtZ5M+F8V+2STX1MFidJLCMI7fbEhu9cxci3ILL1
KoVBz8BObG9fT8maoB5WZDeZJfk6Ia3rV7BffxR3qjih113NFMkR8L6IU2znBXvUIJFQABhTrUM5
kAp2qrA825BX8APhwZxKw1TkTcJnIkfO3SxYhIINm2YRYMdMA9ye9T/d5Q9d2zzDwzPOloE7pfq0
63GcXQ5nsKr561VxAaGetG+QrS49nTzmOHiI9+cUB3LDYuB3OGRQAGz6D98k8uJSSvSGDM7bXorG
zxQMkg+sU8kCK9MkEugFcJaBLZWVhfOhKLPulXtYzvu2n3mI2+/c0qB39RXM6dtexcfHGe4EtVT/
R1x5RFWNQAYL3G7Md7YubCo5aYj8nbSoeoEyfr7rkOs+EeBZUUES5py3bgCXAMmQAlg1C65mrP9z
x05axfygxu5Fff4PtU9k3D6xCo0/aLroNNVdmupDO/0BlbR/LT4oGGum4DdWw6ngVZmLuK1KN4tK
1u0C/Gk7tKbba0eJ/8aX+xhptg0TT+H2j6dO+Zp5yU/R8EzPxmqpkMNUhvQ/ACkJwp2MmNijhASj
lDSr3MQHmYGSBMn89mbawrqEIA6xjN6bUEHrSPE1dJaEL0XWDq2xQny6GP2TbDDljA26OjtwVTyT
O9/dmCxmMnnEn4yUU+Cummc2YXJkZLVTLxZl3Lk6l56K64KzE1JEGWAoqsLOhku1ottUy6zXyklh
CP+BuyCp2Dy8RPMtw2trxU6gge9Cpjg58HCrc/wPrKYQ+pKpMOnuw3ZZ2+iCH3Hly9GOiu4FgwuB
V0/ZOwd4g2bmcylKzxmxSjmwC9sPkT850EO4FTbM1fViryC0jwev4KwrDLL0c5SlmbDLjfnGCZiU
vKj009MIG91LRw6fja/g9Q3Dg0K/JcpST2pBNDSsvZJN31/fMVMKA2gP4GExLto0ZLSWNolSgxD+
MNJ9m0vtTgcHYIR/Hp6NbWxRSpgXw5NznADZz0XJBWA/HrJdvxsXijDVjm85u/PY6fSWIY13bPRW
VOqs9rt3n9K+SpnaE37V8mB+v9otaGlMmn4S5xGE/RRgr4cL7/wWw9ZHoHMrmB2aFbGVtwSehSBH
EM6Vwa5xgLJcRv8myL7JNL/9byrRjHcVT+80MH7pFCcfHvb3gaPw0xbn8//crIvzDVhRwx83ZsQX
b5FyX4oHpm3oxPvd1meE3qALHKjaruiAgZKT3/3WIOcFljoxbYAzWxmgXHcprlYRvwAdEjKFde9y
hrIowUwzoJb/SgKN9o7Zh/x3bVVqmsVrMmxh/UjXIglT0sklmvkM7sJDLYfudQGn6Stmxfd/moJX
iOK2rvMWeyFdLXvxfFzOGc8hEAQsp2v34Ka3gjkDPGGwwPXbZL2uRvacUeV8uyvz3sr0qKk7cwWr
rpcYyAKYAeqr+GpnQi9th4oK7zV2+gEJqfhj54vs4BlB6DiC37DFUH2pxbB/EEgYJfPxHE4MywBf
ANXLNbW+tBHjG2pCksQRmMipEK2zXfvqxoCde3I/Xwk7MvqFjClmGa9ZGjjQoAWYkxZiJMVHILfQ
pK534QXD69Z66nJIFc+VwU/vOz8n1xxOAnjt5OtHQVGquJ9t4bnfxfJJ0dKf4L/a2ZLbTvqSJycT
p/LyFPe1XLYwA5LIU/ro6LE9e8ifWFAtwvfrr2EdLt4nSSQgZUPLv2inBRpwUrTDFp0aSpAhNDZ3
sfOBXLnfvE8xrwEkSybP3ZhIeX22ePI542VqFasKbaknagl1i3hTt3ANQlBs9zz4d1PcI6sUujT0
5GYE/XuGoE41nDlKotvG4AkLHrgL6Uot0NoycolucgyEq1CS0Th4lHEtmA5Qe7XL3coFYoojJBZc
9kj9w7MLXksjFVTekv1u8MPa09ebp9VL2XPPlApQ5SFYW6ZdukYYYVZmWIXkBUAbKrNycifF3xTv
9zf4boPAdRxffUxP1jwUtH3mEBJJvUgrvX6mEdn6BzUXgS1CvUZ1NMQZX6qwBli6PQhu2FXMuGnp
ZDwKH/uhpCHQjGGI3peq3TkeUL5b55pvmqJwy+zQ6xvkfDBnpcLouqLtj1W2Wy5TjjmDLBu5lCh5
DiKQhiEBT8WAp6eRE0OLyLzzMc6yGXyw03QcklqjqUo0okdOW38NIjBSs7mzmGVTZ6L3akGsdVws
1WYnrNaqz8WqRPEeq/OZ1Tqy8/X6+QXz+9FyNr3MYZ4ZkjAu98n8vacWiaWz2DnRPaATnhrkLNWg
pYJD+0Tqdl7jUFVh5lZ16DIhPZRWclNTFv8rlX4UqUfCNjCbcsmINbnONW1I7hdGVxTXiXs/A9tb
5zxogTgdEidhsgLksxfzPGgpJiLL7+s6zMJdrKk/WeqRrQU1q9U02XdB+pZaA7a+fhESkSH3h4uy
ePY8cTACXM9gtGo70AYqk3zceEuEx6lSUeGqWOUp0UHPO61LeK1owwG0fI0J3PmuZNz4SLx8VXOO
hhQAGOgj/HtNVXkTzAuZW2NV/Yjndm6ue8/PMU2jMjwuXfNLEDHAPA0Zdt+BCvMSnW6JomZgUeUw
Mv3EIDTg5pK/8kI2A0wQ/8/aoTkgskUg/tNCElwl9hdrTurbjsK7Q697hlS8b5vPwDF1r0Dg6MwH
FgbwQK8TX7W3s3C1FMY0NWNSXblh8iX9ccPjIshXSlhc6dM2oI85RVsyFrk+cDsmBWc0qcsaex9d
OJHUEj9uZPv8GY86u9zPkqJWsR3IemL3Wc8MOYBt6XqyaDa16jB9qMTMy1u3Ks8zslvCqtXkMv3g
dxg9v6uC9M8nyn1Q2V5Z06DURajvOnCdRyoGGYluAtvvR6wEUkm3yqBFtMvSNsJ75zuX8t4FIxH+
wsWS0FekjOZRurR/IWRIq2/VIJoCmWGlYRZYydLEGHo1BTXWdLHIshCqYBoJRK6ZfiwOmr3cDTj4
I3CTRex7tpPRg5MTYSnpcaQg/6zTXwu5RugC2ldbsXazMVnLMtzhb0mXRI5Me1pEe3GPTznIxs24
ycpVYjak3rZJQC2ejGwFLkguHQDdyyOTB0+/VF4pPIxCfcjN81L3t7cjh5oDGIOMlu+l8GILehxv
h/L06CuxyZQzhTr8W9BwmPhyLbKtveipakIfnE9LRzcgQXzVpW/m5918TFYMZKW637ZjI1oecStJ
12LgS40Lvn3Kf4JgMmKMGzCQqCc2HrioGcgXGmiQAfJ9z2pw5bEEnenSZGb1jtOcgs4WCvbIeGc7
EVPkvNzj2gY/Age79FIkiklGVuL8Y5F9IrmYLLqgQaukl5YS3z3n1BKzv9BhEtLyNv2kO4XLSk3f
fLxIcIhl3g9l3Rqv5a0zyC0Rs7YPQQx9tsvctCKJhS5k7xv3XJNs9kaD63YsNhx/0hZGbXnAn3BX
nfv1BHwo1yaXeIafW8o9+m9DWpLrM5darNPkv2dqx4BORgrSDS2mlL+95/nNdUzlU6UNz6l5xKWN
vZVc764hHGKxl2dVShCsI2XMdhd515xdShnoeqoJatT8tCHRF1oMLX4BCBs1ao0A5VXZ3scgVfCO
8/0sRVuLAAASuuSIrzmtt/KdNvwCfuKsNwYcqTWg5OqloIvNFl3WP3pfnoJwJlkuaMRoVdgGY9ja
GVG7jfxZPQzwPFbgh+eG1bDTCxElmpUHLenhmB8jXKlicdrluM3ixUMCochtRa7JsN7p4LyHj7Hd
H6EDSJi4j4zKgnK+MvXCRkFKSTh1humvvGIDd6/oTJKvtogUg45+MZ1spPAHd1rjG8Y+QiFC81hW
Xnn6Ll0LaIJkTfqb3O5ZZSaAWp4k+WeucApOG+jx74rS3ZnGJj4oVSG65sdkFRHAbsBCh+pec3jI
aU36djMMn+bmV6SF+og31KaAk7t5D8YEAHPVSmerbmbuLMb0ISi7TObS9xKw5LINNcKvWxImwPBm
I8KJIN6fDILv464yhnJch5MPSEM9KH5ERAVnx6tz6JtqFOpzH9zIfCU3mJKifcjaWjTPYtM0jYqu
FAr5T2o3THoqS/3lvudaIQUX3Pt50eDY/AW19qXJSOPLGhbdUflCM6Wfh21dP9TNQqscC/YAI5dr
73gHZnDrbuBWuRTfnWecvsewPUxrFcC3oodq1myZkSIiWYCGo7Zx5QVIatJhCYDmWJe3uk6xTt85
4oqpKKKy4uomQnbVHVm2h//ocdl//P9S6INGf4fXOgzwURLCex0dqCat381hGVTruriMxgmFsT74
083Gp8hZ/8ahSCWgp6FDL0LrRAJ/dWOAmY/wCMPevU0NqUc+wnxYkaKXalR7nk9CImg9RvqOQcxU
K+qAsF1/TQoqhdtN9VUe5/TCRwV6g49uwQbpvlBeT+A+j9yl8/Mr5/wi3NtcFI6ydAi9sm7QvmKW
axyFCE6I0uwhQav3ThtW4hkTKh0+S2VQgUcZlY1oIdDU0lKBp0UU6q9YuJ+3M+mJbYInPZWoSqLO
mvNx/9BF9m5kACUFJmKPB87QXPIYd/KlsmGabLscnfqJBMlVJTvFxLVHnc5UwSSgLZXMtjS1b0Rp
5TKSPnIK9a8M9fUqxjxf1y+3DbD11IzeBFL0501H1j1zDqCXxbrFsE/CRVW4Dz28mm12d6di2ZbP
9kqsVQ+BwQd/gcIeaJyc160IsBbPH7mTET8cGcsZ3Tq8k9ajLyVSH5n7rHoPga5rjTeeW7l5LFgn
4agJmJGhuJ4t/aTH8gNzGSfUE0/ulJJW7RhcwRmZUtDyPVP41D2/gAc1+UT6dc3+O4HFRWddNLdR
EWp0b6dVIA0yFMCzFszIRxAN9+wyaluWYzGdCwuILAFGusOhczYdzSOCWTSgzi9XM8HIxcH8Vy2e
77zsNYJj3zbpKyIK9WoZxYYS6qJ9WkG6agYiVS4n5nsx3xSnVl0m+LlCqnP0VwXk9br+yviaZBGP
vjYAWCjiHRpwjzikfgwWLeqy5CJpL+q5Fq4wF9VugE+sz7ZNBxMhNx541HBrj/IeQGYoTeuqFMyX
J+HZqlvfaJSBThUt44LeLl7gXeWwKotXgyyln0z8t3n0K9350EriJYiCKFhd9kOsLpXlwmeZJKxV
N1c4Bkwt/338vlcmk+xf6x9Gv4cjiY9Y4ulZc7N+raQW2DEPEwBLHiieN63n8UE9u4TXvl666r21
QyI6dQNIv0mf2vrS6mOxup4gHXWM4kJ/VG8tikM7AYaoXitAxjY29dGDi+MZEiGijLNFFpbadd3V
M6xs4b9/ssVZp9t9rKyuluSKK9UzIJuXZoaE1C3UeyPZBxSqG2YTZWipyLNDBgoDZ2k45N3xEMZx
VUd+7oeEgrJIgHymkshPX3pW21BNkXI4B1S0PaHIh+T0WW2ny6X97NfL4IpYPaLbnULIIDokachi
O3c8n/Kb/d//Dg7BwBRBvY39mMu7eSD8HRXoGjzvEm7B1qij5rXskRAI0ptIKsnG1uvytcD3tJHZ
IiWxLGmF8xdqf0RDkzvpfbDyvNelXfFuSwZTMCdWrzHHChFxi+7J8OMzlJKttB0qo+c6W7tXKuzF
GnZjg70ehqB1Ipu3crqgwHTVRURZrZRerluYKAnHWKgm5YxiGNyjXgFUGEMG0NUd6IKg1YSwJd26
SZsGJaoTUL6lAvPD2TVd+qR/OLga/2tm4nYPrKlzU7cMwa97vwry78SUk6XlanN7EDTQRfUSNUrs
dGssccomDDM+bef1krKItl94JqmESxAJg1pUIgpdMhC+jj0pyct6BH9GWqa5R4oSTdF7UcZChaLg
lf4aOx/86Q5PWRv1YeP+/xuq6lVdHN0Uk5z0LDSREmcbQbPtvOpiY0DeoddJ2FgWCl8A6WH5S97a
xgZbGgg0z9/RsY3g7HZvTXvbvMldFy5pCP9oUM1sv00dWZYgslwrhMezV+mzhSQpBziNwe1Sg2EV
h5EGublKUOorrLBQzxt6XP/RCYrhHH6i8wED7MSgJCTQS4ydf7qpGXenoe/wfYV8ekAt8oI7hlFH
K07vkXQ6ppzNUAdKSJP+9OczhHi952pajizpD6SmFRYYF1c6tAacN+I/eDTZq0JVQTPiAAcQ3s5w
bZfSVpzOtaD3DOEidN1TCY7pqQ6ZfzTh5aQQD5qEIbIwwFDAOL/IJWxfMDtAPf9NHzDD3xqF+JIu
7ZO0IhhjMtcUliCxkNBLf+nbCrJ6P68Li5NtM/QJyIBexsOvnNXuhMknk0Z/kT8uwh3s6FYsR3vV
KR8nIkGyZTa0gkz8PS0T4IVbf3pJh+MOjrAZE5YJ+y7RUWSPKnVN9zQ4A+iDCN0kJmipQrYkXBh6
eI2Lv4+xvbzBJTT4EXm4enpJxQ2faIz4KVeNAHGnHp/Em/RQfURVN9K9BVgb2tCSAd2nIIwao2uk
fiu80TyZXpi0AWjirtZRHxmt8y+uui7VnUKcWaL+qTLkqIDTtajYTIpgMoHYg2heviRQqZ7+aKge
hsqZ0llO0sbxiWxiQNk6zB+Fyj3EC3GsaapzREJQvVfDRLv9PIW10hfxJgm4dR/koggfoG8OpiiQ
yP5esiObkw7H5VAxi/3BkS962CvW7QndL/96r3oYcL9txKOBFpib6wcRZEgOZYd7MVVDxiZ5EEfC
vn6kci9aX94UeLQiqIC5FzxfBUdhdgtdSyRtbZWqRkj3ZHIiqehDjRXWhlgBD9BUM48KcTVfDxOs
A6RIhCrQBkkMWjzQtrIjCRi2uratbgXugk7L0Lb+ULYKTXY4ZVE0BalG0NoydwV8psEwo8kf74yv
LmQL3SuDadtng9blkgOG3gi8EnhjLKd1fnyZ3NlYUd4cXiJI9l8D1e0KgDp0mCPLAWfevJLv69Nm
4rmYlVlDOEEnGbk1qv33iBzrvhxP4XyLrazMG/h7q8eTjnsbFypyJKNZnDRDJnTNcrviU0wOqcft
VlvTkT5howP5+dYRrctRs0RlmIKN5bo+5T+YgE5oZ7sFSBLCLNLABIxGCvFTV3xiSEIHNaVrgudM
WL5LZ5OHJ56mf03Wz2aBx99Z99msw0Eyl+giut6kI8lP/xFYdcSjTJDVmQww4BLVerYUX3/Co2hy
J6jhhjOGUBHIbx0D5assxpNaiyjjCkdVHTuDzOsANVJDvNhvDhEsdyNvLUSQ9g/Q73kz9kYfOzqP
u65XLWZukMNKV3dKkboNgLE4IkNrVBIRdvDSQC0Sqy23FaeTCgzrcSoiXwd+kLVtBNLsEfhEsySC
gE4lLmTUA/ld+lcS+HXBqfnazzVXEShKs3OYysuEmVDqsL3BE9Pm2D1dmw516j91MJV3LkZ6meAM
v3fGBHK2uvYIAxQworj3geIpfYXQ7byi/urmQbeUd3o3f67Vmlr12vF6JOE8SKAf0bniHw4fAvWV
n5wC69XB9N/qss9BXItMSsV1jU+rAUq75rFoE2N7d45aWvUrxF4DyFrlr0JCR/dQ381kJMjj04et
NJY3yE/bXCJnUH3GVkGZWPE3mjJHwZkKxpultZeDk0SQ9T+FXg0R9XxRUQluwPry5FZ8Nl3US49N
77T5EnjpG+gEl503Gh2axM/OD5tsdeaDDu700ocbM0Ofe6NUwKm1OhGfzwxF7z2kTBCPuK+xOOx2
zRNqxdhhVfl3LjATqosRiB5tSCzGfm99FxC6iWwtzWO3f2c7zolyoip8omSAWmt1OkjbU1m1fnku
3Ke3XVEAanicF7k5HfbydlmrakHTVR6bTkv5aHFrsmJ96lTCqM1eOBwVqzVi0v/VKbX419Sgswa/
4rS75CnvmpgNmHYEzxFq+rHqdqzTNIMXqlKm+IwAUoYj7rm//VyVfteJixQXkuQzR9sWoQ8EB/l7
DwRla+WviWht9zQwzH94Er7DCqoO3Wshl/NiZG3Itdice2pz8eoRTa4EyEZ74oCsuOIYOUXTnfHE
p8llxJbaM4ZykE8ju660yHBClLbmEiGKl5Hp+s5B4/+3PuS7baZ97OZKN4zNg3sTNvwONnbtLgBw
JqaOIERbQgv4fwWvSm6TtIlDCMYaMrTZmnlGO8yQTulAZVzvYdpf6ra6MunlynilyV7kI4pFgBTT
2GMLahoIp+GZijkSO6tL5KavscVDE8Klw8rB9MwbqsPTpFq5oiDy9oCqsw4Vs/APo1Ry5h1lRgqu
h70pnUB1CsqPPO9H16ykdt+V6baKLYVtbqwK3xeRmMql4nBMcYfjODaAwwbnJHDLziAdk2YHrZi4
6a4/IbSmpicwixf1XEeoS9WVuRDXcnUUAKu2GShWV1HpEg31dRzyDbMnXuK2+GBlYnrnFrlvR2Xe
jiKXwN/MrulBJStO8M30qqGgazNldclLpcpxhZW47gpDx+B7TwflksafLoqX4P40YacI5qtkiLb2
/TsyYlCmKF+eQJmbFcMGKKcaluNARAKTCT0/tDlTPxJSoJhjK7FN3rIJfyVeMW+f/Ufz/8UUKkyG
QCu4M7muylQjb4sO3RMuLJfKggEOQ9M74yefy6rtD7AWUKPTQHaMXMLMxPJwD8+8VpxYoV0nmWsN
x8ZoTB3rAjTRDzUlMwdrDZHi5WCRc92xqw+9AlKfhJz3YRK4/Ks10c2Du0UHMnkHexRbbzO5UMQk
c83d9kYM3ZE/yih5msMJL8IRhBaovmUZVnvy7A2ZthxEg4/KmvQRQeE6yfLFsSr9005tiD+QbvT6
Vvc01ybqeIrW/sBzEUWgbu0+AETualh4pClNzeDrzLI+e8L4PTItbZvyuQe9BJGs8jX7Q3yl+zJ0
LOl0kGeZYJVObeN8sp/31M3m42Ibxcvks/OdQtrrKi3H3WCg6Rsms+PK9Zihg603SW0OWsq6+Je0
nYFqdL+NBQA4C2PoyR8x66fYSjK/OvhDTMH9mo1Nka2LekIZaQqRFC1k3QUNi/fLtMpMmzew/yvX
P16jx39o/JETgy7nEQp7Ly+GkvZkzMsyjIV+C/LEwIqIyuDer5xppIX6CFr1VIueRoxw3+qB/pSB
qRWTgvQcsVfXFU0OW2zeo7ghCQ09m4XANomGUbz6mYDnS/ZcKLGrwsqYz7CUoMMCpJ3YD16vcgPI
ZKUdThFnVQYrR7NvdAk/Jt5eWyuQJnakjDl2HpWRChndS8IInWYxq6s+sR7a1gaA3K3v5tByQnDj
ve8J4X1EsXqjjNitQlgdlDoU9o44YyTz2RPCuiEIoEyFiXiUEcMz/HQ4O0cgSyq/AtoZQlSAnM7K
D71k5s6jasiFKRzosEMkeE8Y8UOOpo8Sy7dsSarIBNLK/jZW7sbtDzK7GOSqDk4/QiVzdLEHzaoT
B6e22kBOjT+cKhOEsJq9e73wWQsgCz47uXt2i2OJx3Y2PQUandtzcf134cwKuqAaXQ85BdN33sSV
HTvK+kwGEYMKTN/VSrhKeEwPbyFGeonaSxNg/jKv/rxZAhWVIjQjHF2FbshbVf4Gcwx1m8MuO2e4
U8Urr8cz3yMCwsDQT96B/lb2w/U0X2ELylhNnDbWjRWpstllFttX813p5/9LHO1852ia4I8Xw/bF
Plwxe5Y1KHV6CxVA/75goaIxSyqc0429/R71bhk3T64x/1fPAQMkCmqouNW3Yb+0c31KPm6Jibrt
4lrcfZFs1nqdkl5RKD3pTEGh39PanC9Dyu2oiFewp7t4LzOmWln2zkXLg7+62JWT0UrreltEiTVG
PF+JXc6O3AiQUOekYhaZ5GsSHCS9DazSCYXekcLn5szp5Vfmoq7b0IVI5R5IevWRbNZvcsVIb/Sw
gwDq+0THKgJ+a5dBYW8hwLEfr51cA3fmFv9vTnzZLQjzT34+tNc4dlGrpCvGO5TEOI2/Wmm25Q9b
L+SkwS+/DYAAxbDPeRMMynLoeham0pvnaErgyLlF7WREIzLz3uSY+8McLO7j/Llqe+5vVFZBYig3
zJLGQ+PifbB8W9NgjwuV5+2epellYgfRkvZ2RkYnq/ieytRH2W2a1jCpXvITbeIzXM0dhQtcyU8C
t4JVCLkxDbDaDJeyy7H+/Rt4cJ4lQZHLi+T6l48dsoLtz+J5rVeQoG3iGxSYamqpy1B1ysw1G+Cl
yo1j6ejjCN0cGp1XSKgGQtvVJqCcUNG2V/IVzaHrblFSEgwbg9zIIiuKZNZhyH143ZxRp9s2nw7U
Nx7NFr905fShMN7KX1Iz0QevDQcnWHaJL2Gt9Vg6xpB123sFPhznXiomBpEdpSklwmDNlR38dmlE
V18wpeABfH4qyyHIdWvOCHr5O4fqVYgNognnt+diF3UT1uspsIIj1EPe2xwC01ug7qP5nKA+w1Kr
xMIPgtsWcWDWfcO2YZ+uBWJcUanYJxNJ8yUup7qg1qFi8DkpjV5tU1CW1kLSgfuFXRBociL8fTWs
/MOhoF+cglNG4VObi1/hUuV6W7fnCNPXT81QBxmHrKLjuWSjxHjfSZO80MUzuW6txRAduXefEFsK
6ah+N+8+Sl8RYaFSWtDUf76t7XHmQXQBzampg0wPc3fCTbdbFmKmfWwV1d1GDkWKiF2iT9B0YIIX
rHieK7fpGRA/s0DsBxXD/Npnis7ss45TAWoYdqqvv+WGB5N+0cw0FW0QoDxwzPYohKBELWlmcGxm
PormH94P3Mz9F9F/VHy2fmSH9ZMj1xY/cGAAlE9hamxjs8gwdY2rFpxjH2fmM5IdvZ9IPjEkpn8U
hRK9eh4oXpdCEXkUvEdKF4OzyFSNnkKpq76pC60/Jdkck1OpxbHANt+Nfwknji4o7REwtTBvDW+G
uco9rUqZxoptp/5k8o2XL6cRGR93D4b8DFom4P7hw4HQMArnAzwaMNy98wMUrdxhIjSBvoW67Q+a
SxugifcrLrGKU7q1fVCDX2/EOQcY6svL0OxK90fq5pIfsSgC8Vs4w3OCSFre6ctvi9pWlvMfWxJ0
C7WDWK9qiqgZG/l/zBZ6U8VjpawEiaUYevLzK8ZxPMBBx3VfjjDZGivWaBs+ymw4141U3+tUdsLK
ZsJJt9GgbOctrffUYHIX0TA9fXYpN9VLGhoZTPjAfbkdhIbJ8ez50wolDbslCwKb1qwbKToTdggg
ObvqmZqERDZVo8WMuK6DgHT1EP2VYJ4RCyIgnvyiQPZCdziBi9OrX5bqxEAB8Vk9X/HqzbyC7wp4
ivXvfQVh1cyy64PkqrFTo0o131LOR1SgcE4h8pDl25VlXD8gjSTYW38FZin6FSyzbr2ZvFjfgKHH
A/8FMLQOhrNqmSeO6W/2yVU/8ghyyG7wm4i6ypAO9+5TkMJLUCrSCksC70OlFT5tEnFmBQ9GakgW
jxJt7o8hTYEiE/+iA83LZm9bpQlq2ZWC/dyW75Rv0eRddwIcWV7lkiIr2JNCCufBe9ieHZIQEE4S
spLPH6P7S9VXW9K02EZCH/OFB+UAmK4h7Ae0qjTZOpRVFGiQ7zsmX9tXt9+Y5+DK2YgxMNL2kt/7
Zs5zHE343bQHKSZXC4zfLdbHASB+yl5dZmaSZLTP/taTqzjjUdPYtLlGekKkWarbEbRQ9VRtdYD4
244Z0ZOe6KZYsarAFCbD3PCaHu6kwAYSMPhi4/GFjU07Oh1J2wosfPt8f1NNvEusgv+XnevMUOZ2
yHy406/iAckMVerDp0kUc2DSyryrmRAbIg3QJSqzEchBEcTX400S6HiR8DpF7GynZfUjceoDMrba
nxc7ZKCx9o/VYBPcx0jrh671/DCwB8sobZLRXP3hH9tu3DseonZVJlGMWtKOn+pEyYW7vzWE/sLz
ixxpz3/qc7t05gNmoHaSbegEfkEJNw6gmEn+yDRpFTs52K2cwVGlyLJhabkxkEyZrEJhJRPgrAVr
rhtaE/s0cCx1qkeM6tbPeWvO1gpweo0YGQjfzmEMMth1wQGVJp8txzt3kBwF7Mxri+YWBJzuf/K5
GpIUxtonyCUU6AWs6EHyrNqDcLztyiucvnHbzaoBWtbLCX3ZodG6ExbuejRgj0NB9cCO8tS4UVs9
N56dH0JiGS8DWrMJ9E0VLZ6G/pvFkiMFH3CJMe2Ys0Qe0qLF6RvrIMIt4Lq7j4XYj5m6NZt2j32/
x4e3IYq9X3EvBcgHorGVWkGLukpdbje8dFak+Ex3P4Qb7vcCuvS/cJQlkwtrE320iL26SxxcntId
kZoZZu+UJuMg5Y1x5bVhApjpnqCDYFM5/25qWhINMV7Uso0YAtmIm6skqsGzSGvdJHiPpqL2duNF
qmgCttsZ4IsDuRt5vVnQ0fgppfNy9ItLlwkQarzqNG4YUmpJun40Bk1qNEh4Jk07jpjI3pfhR94U
rC+vZOsSA7Nzmnbwc8olzSJD7pCxz6lCriGoBgoT1Hyg1hNGjyO096rm9Y3QOYU/WKU+Ly6IwvTb
YDOxvHwT7EaJJo5CnjVlk03bdo55p99rsRkNZKSokALAA/P99JGgASMx4gFN3BhYwOB/TRXny3Rh
8U5k6oHRt+tNVrO3cZ+9lICf8e4WARZieX/KlJI6YmQT8/EguuxpWvQl7Zn9aRXAXJgM8FN5tBaP
HvWfA1jWqgz/mUpz7Sb/Y+v0zsA6rWUxDYa7hc10Jj+Va1xnVIY0sXhrU+6hsE8M2ITX16AVWpYJ
lt6bg+RtE47ObGRcEMgNH2eJurJS9h7lTeiF64VE3aHTagmT1pH3Y8K/rRAOMPh7+7Hzp/XzoIQh
LO8NKu4QPZl563EIFaCdc8N5n45Z86tBbDCV8dRD+5HFUdCvVwtPcfrGUvXXWS8tbEpW9LTxkGxL
8hjxCPtWirrdQJvy1g0OAxevNooL2mHnIHA3BmsxIf7YTjQFWewBNn05Gbcjuhk/vEsYYo3StWpy
Kq2bQiW/4S8Cirvk9nL1k4+uLZ9CL1WSRrTQoy6iT0BSP76U/LqAL9kYfpZU5GW4GO1IGl+CTJhU
7v4TS8wG6mTG3FEkiDFbHVJ3gnvEu+7236pjIaKUnLUEwEtWbCs17EUtv+sdL3waDkpxlTzghqCu
HchrNRytZrXV/EkS3CrGaQSE7cBQqWfBzzeZSw0OdGAnT/ltAo0nG9bxag3SnbYFYBjEJ8CxDLHe
9K1K5i3A202/61o3rDegdro0hsgC4QH5AmixVAtAvu0DFlBqWtmE43P00ptpbBXuZBJKzL9N4VYm
VIP195/kfjKk1N7429P20PGDnVmpg2vAQeloiT2ilveCf45mKUNgUg9DfjV0OIjlDYrQFKztyffC
3UCzjEJz3C0dYcV4iRBN06ViCF+WQlJRn7BN7BE2/s6gvsY1EJLNb7dbTGO6pU5pKYLju/wnqtVI
feWJjYg5WN0mpAxPNyGUNmCzj/r9ugexCMzoGBFZFzRDq4WrRyV2WoOpZf0AwJHjpO1EnSdluHCL
6pyoXMBhIWB2D5wocbykyM9XL0tT22o66lPZTDQheTet8jKNqagR9ptAjCDfkFRgV07dgigXYHnC
s+Ql4RrR3XzYeM+MUEbtXCGg0GiUUQOhRHH0WCnSzC4mgBtf+qe4GAkcs/WUmo2IDMoCmaZ+H9nM
axTU85rFWEM1eXQXF+3qGDi5WnFayg3DTXoKMolk2I/8BKkxbG4zxhmh3TJsiyBKO9lef18U2Bve
TlmQ79jPcUl8xlOpl4ee+qnsPQjU+zWupg5q0sLaeiQ0lv4VeWIwShFQi1nSYLTjIjndNK0KZzhl
KkZd33490594JX89s34UAdobCPp9R2OPgCLQ3jS4nT31D2Qm73BJSPPeqxZv2Wvhx8MtfT+Hl+5u
S2BvezP3pkpUn7DUbZ4eMgj5c1U34xunxQpEgF+PgxU7gLeVSWr4XnblimkUlgkMJKGIYVRCJF0c
jEoL+Foade73ZEZ4k9Nwse6eecFCSmU8c9HOFS92onjV+Vdpc38iKjOhl0soE8SteWN8EXQNhGWk
P+AyfyJ8VV31jE1RPhMWXDzFZD4sC8BUmOPm6qLseq5C/yfOtJWBu2obzKOS4BkEfmmUl2+hvqTs
kEwMA+OQzYYCFe3yv5t1XtarJQj42a8kviDfezsEBQQAWLxihN0HTj4vAN1WynEEzi98JRBUAtjZ
R6USPXxPjcKPsJgvzUxtoWqm6dwWVAj7kGwOigd1dxIpVq4yrdVKAR4nZJNgBdFzjQrV4IHVDFZe
cW0gaFmMuLXBVJ89rQwZWOeyXweiCm7M7Q+CFR2zuFZhaB5VL0HJoLVapsfWsOtYmVM6AvLPbADo
l8DJu9LRS9d8TiZ9ZC8iiIJQ2V3/EcqT0etppLwp6Dgp5/pSLGJfTQpDbdUU884SFCbrACGHtM5V
tp12iz16mCatmeC2mo2HswhHo0wBB9MD8S06IOuz9lAHevg5rshYut2uh4gUeyfIsb/a/JdszSB+
uklHkktUQk1LHgywFwhUmW7N117aialFSOBJkPryKJlPsT4VUIKwo/DAW2tEMHN9wr/1BSxWZang
lbYZxYdC1HeTu+RmnGntroSBS7XZDdrRGF5ERbVUr8v0rNdUtB9PUaVvYjdf3yYCgJh8YMxTMpW7
bqeXar02qTGZYVE8cs50N+GeZb4JMyxKQBDhs5X7WYqSNPoSoCFAaW5zgDJZqCNptd7q06u4BADb
jBKd4PUiuf2RmSvPY5v65raf9e+cS2s7T0ZCWZF9sHGcrmwoa0Y/Ja51el9728g8f/S60A5iOI6J
0TMmboD2cZ56BDFVsIpd4vMTSWUeoj8/hhKYqUB0/u6vyDZkcyo29zYrNiKkrZu2NsQoBLXogxPd
m71byFMhgPkSx64Ikkr7j/ZmDOOG7dkt2/Uw+9ivEMJE8I44sNoChZ2LKDoc/mhFJRfK8APTJhfS
e+980joHGv7NkSFtYwRU13CPH6DYDFI+Suo7rY8jhjSwCaTMCr+WqTLJNG8GT6L5StcQcLRot9wd
PQQSmF6prppENWghjYUJd6LLbWglqfkOXv3QozSeF+UK0xCV8NuqxPEktvKs5BP2gJ6jYcyNU756
cKgyrktbw3xYjVeCrJzcuQt57q1skqZOwbkXk476moFRHarxedtidk02fj1Oh40uAaGN8hLFxpIV
yza/sSFAuaLVpNDhQw523WLsCaWS5YtQru88uTuBR74lB4OHVhkIDkoxxbmZlBuBn0unP5xlSWli
iZTtnuQbvtOTOadl16PuxhNIA5Fyd77Sexz1l4uvDmkhA/H9BGpLDMhaU7YVNgxt9IEEDbIHrpnc
5eYdkWxpPHzd+dbmewSYuKO2tAbFJ55UU8qduWHthgDv9Lrh0MpIRDL9ZkIU/obLgIOIHiQ/k4W3
Ipg8+qAPFnf3uLpHONPmgi8J3MximIMBpR0puCrg9gJ5QYfWqyCbvCDjq9MFQBbuA4kPUlLvljyp
MfBCZNhvoifrtLdQDyGoGl+YnXzDe8NCfix5DXCIKOPrpDHELCQzXyu0UFhsMAzLKYqpWog/2USh
P3tjAJJp2CnI8P0PwtCxX51UeERXfXet7Gp+SYNJO2+gJUrE+l0gDzlmmDs4DtjIYoWUj5asXQic
/bcQvkHdldqWuRWOhNGrFeZwykaB50yikmuxT/LlsrwuibOKr2Zt4cFiMouVVNGfHZ5WvvpF0IFl
r83apZKNBuAmZy7Xn3MgE7rUVDo4HHjLn8XqQdmgDvXXpMsKmj9eVDDSWlbKTp0F5YBnuadpDry8
P81AUAKVgG23AB0v7EnxF+ga0sd3F1xL/aNKsWMl92SdzaUwZlZTlARvO6HchKyd3rJWmFVp7EaH
nJ/MxHOHC39xcd8PAJ8cSNGituoYgHS6AwD8rXpEEBjlYG4UVL3dntngwucbx5RRX7JFtslKRgyK
5l9bt4usWO6CIQ+H4alTFGm35LCethSktoG9L/bRZG63rUed8VMAibZpd2xHYvksqb5nIJ9/GqZV
xudICigcEnhqhyRkHssEMkQ6TT6KUWdVmnTTv1y+sfSD+ILtwitTxgxY4p20xgEYoMX5Xumbep4s
W678aTvApIR/YaEJEFV0gr4rjw/ObbjtXNP635e7Q5WZ3DzUONLF9mG2JXPXml7BvjxQGoDQ2DdU
uKveffxI4JqZqE9d0IT0JefZ3beQZzEM89D10QVXvCwlc0JhlYFXRq65r6DAdisEJ/xepBCWvIUm
ilrVwetXY8bcBijKjQlaQwetYtD8va+PWi/O6T9cDgLpXf0w1xENCZF5CxdTfQ/cp7E93hRdkfZa
zL1wVoJQSlGoHSoR0z6MKmD4W9bfZRdFChBmeBUuns8xQIDemOx/BJu2YwmMyyINFnJPzoCWMo+d
06PITE1OIqnJ6LwI3qf3eyjjEVPnBsFtXaN6i2YknnD6Z/UXH6Kd6PlC5H3m/uxDacDRWSN/JREm
9VXjCafkR0boa3DKGDTNaR7sBXMMGd+QjUMpjqrfNgaBQ/TD7HY3nJofgqzK2J/rj6YET0DCRO5E
TeyjZ/PlyEUbLbIkcSfOdNw423TnElHxGi2njpYJlF1Sk92V6iTz3gRMUGAOcH8NAhjo/l5O1nDE
2+M977DlvZ80GStYquR6Vxh2UzBMBfU18bgPILmTuuESGzx5LEYWQIvPoPSqVhhdezNb26/gL16e
VSQHLKv+b5cYNFgpEkgLB99xXyzt1B8wobqfLT3u+3HlMfmd11p5DkfsgxhWbY+T4NpG/LYVlJGq
fO8/bL8BysrqQCJuM5oBx1TE4yUqVa6NudBMi6o/mp/0/tFQTHbgldsXq/3EMhSN0AG7eolTOsex
5hKq5hqU8cvcjeAXsAOU21J8Nfk7o2LYRpvPCAfBKfj6sMfAoO4uqkWDVl3BG7F8zMEn59ezmqhT
nL+lQvJajxEFpjVfVb37k+uPJIxeUjeXWhy3duF6wCAZW4yKUQxBIFjoBLaHMER0T9aIsBZ9dvRO
1C7VleRkEeyGnoug6WoNiZmGR1z5jiOgWT2A9yhUF1gQk9OEp9SSfuxW54v6dAyBhP01Z9/uSobR
x7WB9mKmEKKjBzOBszKsbhIJrwhioLQ30vomN9z+jKGANMK/tZPcnrzzmzFFlSbLL68fA8iyZK+o
G7UeTcs4uBzj4FGe+7O7FfGJz0vOdRgn/BPvy3gavdu+9Xop4anW3pudO6US3z2LsuoRacwE07wI
IoILvdAxJB37/okzFZCp5gUSD2oZvQbZUWZsvftvhw7gBURYWlx+ME19QdWAd2fhWutMhvyJmOom
j5yv1R52/PnYhXDmf6reMc/ZY4nC6Dkkto873Zm64sOXz+q9MvrAjsV0v52xlhhxDmQJCkviu2td
wVA4JBDG69Ul4xS2ey+H+qAJPKkQeWVjHw+DzXdLzd6e6bSDMABaHPWKq9glqQx1NPwcpRIqdSjF
lZXG9jdirZ84MHV2e7dKn1IwvnFPfzSQ8ZYgD12x/qGVElnxuvzOYcjc5h0ME4MxGFECtxoF6fHO
uXw9wBFIlN+znM1pPE6tF+hwG/UEq+0FN7vq6cq2fwSJ3enPIPRct0/VFXkr4mI9bl8gHLWvrKv6
VkwCbgn+nA/OVWJdLqPr249iqskukS62a2+a7GgvNlVsQZOFJDn369egwXvD23boOlvUbWA1V0ZD
QgB78fFjMau1mGFNIfAtarARBuyCNwfHmImEYBa9uFsxi3sgecRQnDCCPl4T3wVAwMlYHxhhIKLG
Zf28YUg4rbHG4NlZiC65ESVJ4vjVXDFjAt5YSo9SRd0fHlJPmDfRy465RvSJqlsYZ6fzjG6oF0Z2
TiTx/Wnrm8TZx+2k5ah25gbDanSxVk+JWst968/wvoEHzSruAnYv1QT2rUmmPpku5AC49RhtjWQi
judnFtqfCjgD5mLiln466fy29nkh9j8LnGjs5b5QITSLA8rbp4VZ278idxIPjnqXiDMV6i46f7H6
bgiQmXFMQm7r7EjL1TjAhFWO5vpIxmMhDb96HvX0qeSD4SId8m7naqA8iDgfsOclLANbKeSfdMih
/BJmE5fzX8xcVOwZ7Yls/h442r5iHznVbvGKyUhXf5AnPSsPVteCPAR9j7Xily8kgxrTKVUUzQiG
SvJ/L4fGm70Pxkt3OyLIVvNXqgPRKr9D8TSUUdfSk0N1pWVWzG/R+7Q3M//CExxzHxRdmWDvalOh
Hj4ewRpjRYb91wJj1iyllgezIoYmND2D+fCt042Nam9G8hy+EfkTvD1bZldCRzNaRxlKynxSl6Vi
tBGFQUsFW1VocEFiZgsKUwyznDCVdDeFxRaju6FA7sdzWEdFMoyR8oGZruzV2ZmZyMiBLeyUU6WN
5zNjEoBtzXSe992+e0E+YFP9yMprngsCKO/OSKhK7gUWOSuhYqaaS0gLNqC0OmuJLoiTGqsUm0+/
7kuu4fwORT4v1/eh/MGU9p0tPbkr1rgj9LchQRfotyHlCKaWw4DUyp3PitCIoUxCirGDb6BZunvE
NASfOFHX8wuPNmPrCnLFPdd2hvSAanjHD06IKoWZ0tWpDQWyHHB+BV1e5KtFMy5DcSdrxpKbriPW
YcnJt1Q+Gf8Cn/aGrqO/C8IRVj1thI+yr69NUcYSipwS8kE/Vs6oxlApc9TPnw2M1bzYJH6f686/
haG5I9HrusEHkeHtuffe6aj9uVhRe24EnD0fh+T4GNfolkV2Be+rhAUO9nwC0DZB9aIWxLh9u4M8
+qPq4VUZeizKlWQfcukB/XzdDHYuX3ecjHA07rtG5glc1O64tOWhGIiGxvbeHw6VPEEG87Zx8ffH
OhET8GLVh0rAH4dFuD0Qs6ehjRd7GxuIm+FfHAVGCzua6V6uOceJdiSdNK9+UneWkRBkbhLNswS5
lSfENv6K421bbrEzzjTjShkJX38WdJ8mz4Rgv24ni1iltbG1IEyHluk56lLuybpr7BjBev2LvfGC
GrdWL3oQ0vrpDkqHC93uA2i8UJHnm42QM71hRj6+uBkFID5CM21KMhUhRcLMa5N6o/qhkRotKFQW
bxKbRNxPE3OF2RyzjNzCUYlEqD5ToGCOjvn4fJSklwe7vHgczbN/Hv6NlOM+FcqWIgM8Xabv6dsX
UGkzPG0mmE+Kh7VctHsSuoCowHNgPGW1WxYoQvO+K4RXgw+G1k5aRO2t6g/tz7PGZwrWAjcqQLsE
fxiLcafQiViBlvIs34Ra/cr7kZv3KHfLRFxT0KOGFgCL4kDPLZsa9IpS116LzyDR9PljRdjrLs95
s6cRfCxPt/uGmNxL2ybFwcWZHYLSoj2N1odQUH71EUAiWYL1Ja+mHWNYtXhHqoXCT331kkK6mDb/
lOz/3zl2goEXkZsszOH9F7A14+SLqR4xy4D42fX+LieYcdj7UP7ASI+18poAgEA7dfBZdV5tIOPo
8fTPrQZ+TKjLc1cNeXO81thg2YXv894/Ej7W/r5CqTgXzbnBJvW7MiFTFMhq6K38Zf5xpFURLQcP
yDNp3HNdEkmPapc2GOhmGa5fr9RtvxUzzm3hLhxNO29Xg4JW6pSSAvNWwna3nRJ2LMeZ+MifyRsQ
c1IfZ8h4Zl/6LyJhhPdYzfdWaAeQGY1ioXEfjoIs2DwDFgfqBjoYS7AdHm0XQkHqKP63DDFtEDU8
ZkBbs7tAULipDVLW2aa11olu5tLefZWGtojvbLErKVS3Z1/peNnnvcofqN79t1aEwOHnCnUCILOP
GHKQ3ZtClndgotOCfpa7fqVNYGS2dEJJOmth1QnEwKFb3tShBuchIpIYdISWSwBV4U1MK21aYV+c
GZtLLrkqAXS/QZcyt0i2BT5pV4d9eioRcj+ogSuGIUVdfzIh10LrbqsrN9B5k5fBsk1xXdDkVJmr
Lm2z7rY2/36wGrs7kpBPkYIR4D6xpFgWel9oFMat/dtlBFgfrhUHmZdYxJ6OJNgiD7UfUHZg6q6I
oPusrOhZEIYSWOplm1SQ6ga+sRU1UsF/dht0wedcdimxdadP/A+mMhz/rFyY1u5AnlsqSuOgBFcx
BT0f514eNRnadt6E6mwasZpVaGnBFNG0dabBs3XNK4yuIPNescOUgxhkMacR6C1UwnYMLf/mAGd8
D22iqkeZkKo9I12QldT1lP1XXVICKVrmwKAsGpgwL6vVPWNpSj508TMs+H5rKP+0G7rThDgVlJqK
LFKZFeegpsrrVQ082qXVT4vKaj4ou+xVQda/Nu8kEYQn98CrE82ZZaxj23bdioLQIcv6C7Pf0HDZ
Q85zGCTMCT7EgYtKi0sNehOHXE8GMXMvLS9MF/vlXSGU7imqplL2hRDp6CZdijOFjPltelxGRC30
RhOmkhtK6ItMsKVCPftGX815ugfx7uaqvGwTr2R/0kisfN61Z2Ef+2Zl3IVwimxzZpRwPXBXVa4k
/jgSPhBV4ZfVY3Ho0/uRY0iEcy0K3ErX1g/5YKXINbOgdsZsDxPjKbkiXtNSkuw5dWMC8Hoxnwmm
qiwRSmMtIWQ1FITfob7OhKDtgYlsAg4JfoHaGwkKO1lJ2WcKKgHh9Yyb+XCRjLxgNUioQbnQ0okj
vAYB7Raki50aOZxXU2zqO/qKB4CFOi9j3vkJyHzRvjRm54QTPI11TkKHF7Ml4TtzZa6JXNyrskWL
ZCJ5LDXadycLMD7245L7oYOF/hzmu2o6swY7t4h2c2xJnuG+TdE25vOXlgOZ26XCyeMQJmMex/6l
iP86g+nQD+EjIYtjYpgbGal94iHQa5sH2p5l8+AknuOVyPI/DRr7I3JObIZsYLtE5oRiFOP4oKzO
25vS02hkfUTw8/6bCMPZJAKkJKwrCUDEI2mR/LMmdILtAh3ikkGh4PgEtH7HCBYvJV/zRkOzbWIF
M5A4gfYwG3zdiXCH53WXpvep9pF53A8jHR+OEAsptWACmww8pMvqJUV5x5QJ8e51UI+gSkUD1n13
MxCHngvy3bKYtJM1IaI6Ixs6U+MzeN9AUF7emnXZwB0jFjOeeUQS2Bm2YDOl5+t0ULOssgFrIXBB
egqboeFH/ATX6a5Mg0IbtYlrV0aq4K3kGVV2rDvDRKAwNkL/uu2nPq/LXxZ940ALvQXiv1RHttKx
Xu/P4VW6MYY4aEEoTtEhmNXGKma1bu+q2ZXdwieuUu89VS9Ipj6G0iHOQZFJb8hGz5msbBilYO75
/umTnSWmhkxGStesdabOsIW/q0cDbEP91TRxovJ0hNNSwYwImF4ANiaK72Bnorvjtrf4/W4xm2HS
jqcBc9XtTgxkEnMmr5oy30YAr9iqMD7wxbrdpoE2fUepGZ4h+lqhKLEsPxHtNDcEZmvhi8K6i6tb
sgV6VQw4qYy7D7q0I6FtjW/lXhupFcGtIOQveF/7PgD3O5AduBkZG7T+olskskmTV/T0OymK+frL
u1DPSNQ3hted1O8SHTSLazkte+01sINd8eqlCCNNw4DK5l8l8nHNXQHx0aBP3Wbo1DmvbvhlcrPZ
LvC26I404NnO5OyRfneCRz/wQu3JgudrMOSyICmFvjnfdXP3/0QOIjNr7NheleAwi28EXhGP0EpX
lCM7omoh4VF9hm538eAQ3405JrHXNkY0WbTS0GyVHR3Tc36wicCnLUBxsGFjN6fVm6l1wAJIRAgY
p66Y8CmIPNITDPF3BxNxtBkC8dDDZ7uYcBDtCnlNxm8uEJgVeFNYQ88+lXh3gUgJBYOaKx95cfc1
iczeEdl4Hm2pt8QaNTX5DrCNGZC95oZgbQXBHkMsxNgTsbjorUsp6Nm/mNeNe8yS76v5f536gRNq
MAv9rky/N4NXVklMs7HRPhto3hiI/pm41NLNTrsUjQ6jkS6CHKpZuZOz5wmVfIvwpy0eIXCOajeT
oHOzgM1wnexrhQmWHutyvdEm1VRoos5cpzSdR4aFKFKcLT05bMhQC0yFXNstXohr+DJ6w/aQ9X4A
Sy2sAxTT3+4HFn/5Fem+b5Wb5Fapr2p/aK0YQbBrwYWdUCSaZT0njbiqO589d914JgaqVVWEKDfa
375sUwBktcr6YCE5XZGJaDg5dQnlE3cDC1O6a6zXqG9FrLrwAy+Bt8MyzB0xUHmaz6veVYigWVE1
hTlhyRewVWGNxm/35wevLZlwBiyUG4uJC//4qXyG60o5H2LbcnHj3wf9kgl+rEjd53GpLuHK3bVE
qzARgX/T72mPZcxgJi3sm8i9ADj8FL6tvxiXpXytcWfV5lVU+BzJJxNBh8qC8R/gpi9Y3P7f5iSz
fTdR1SdraQ45bnwNM/eDGQ34WOJ9jjuzJh7xGj00yT56BV18So61zkk9dFDsgc0/qmXZVBAlRhR/
8QohEgxqUfJZgDVjCJJQ7X8M2K22CiMNqrPCS2673C5PVIZVjtPFAUoxgRZg+4aBnOE5e1/9GKbL
fciEuHQOR+S2V2ZX+bbDYgN0DM7k2OXsEYlKfmanxX/mVnJxfp25MBa52NHIvBc16YPuA1y8TVvs
triptfo4MXegrOZbpijJklcOK1ajXwGAoYxC/fU2/O7bJk+nSEUNTqpuPyUNXkq8Ibxh6gcmSryy
K2Cj5QoI19tXUNEWEXBLFp1rjZdP9uOJ8XEKMX4PS3J9RHzAdJjjLSwXoNPS2hmDdkZjLSL+RVZY
+SYu0xpCK6D8OXwBkcFE5O1a/AgSGv7y9sbugijiwsXSkXRuIYt29qQQ/RMmrPBnQv9cO/CPlwG9
PLYCb2L2A7v13skULE9s4rWYPXNdXawMYXCHVZUeRHI9V7pO2C2EPyxdlDFf+dwklO2KS2JIAdku
NYrwhjY8dlK6hdxsF5Dbn7+cnxTyPJWDp3/PyELi7w/anNiBDGk7k0EtmJaeeyMvSy0rWtRfnBDX
R2npoIZ62dQEh9M5Mevuq1SFjKXlNCebaAcC+FntdDvbrurUbslImd0osb1J3WmZZPMG/ELygCDP
o8d/3/384t5glgrh7FE0smUNpIWItdxJsYeY6DNz7c8fs/fZHvVSOOhajhyhGxJFoOsXJvjqhG9W
4CF/+MLuK1Za3wzxdKgVRqifc1r7m0o0dy8ICpWYx/4zy3cZdU3mfxnpjfKT9DzHVovyAS7wiZJT
OEWVMhid1X/M1CMb0OGrgBTshs+NT5cn6nQv49eoP8wfsS2UPo37DnhCpG6mpoeI6y1mReCupIxE
3TjQOwO+W6a7DUYfqqlkDWPPlljOgqMdehrPtQ4ojY0nmFtr7tZMealTczSgz4n1orJS2J5s/h3O
i6ZFwvw4BXJMZdkPwOj5bPraZl01PQUVHwOZcxd4AiWzR4iJS1z5U9mZB4PQWks9KHgoory92bBV
+38Ca7VkryNVCSFmmumzpUp0BPUwFUNq6FWlTg57BPEbjkBcaOBAZuzXjZ+rYvxOP/sWGANWF8Aa
ct0cvJ3veManj+q3vQsUIJzGbb/PJA/MAaevNHAUUwPhFs3Bh1atx50D6P9+cInF3WagNA6RPiQC
PI2jCVHHJ8RC4kmTi00UaQYmKrLI0h8hZSX2vshTqW69cNNoC+QWZRJNLxFVXB5HetQXcjB70xx1
+xuUKWJopD9sWfcO7Ghh1JTULkdRpSjEv/2W9dC8RgfmrbscH2nxLM9yMuj04w/8zkCXe1Pgv0sR
pm5d61b1QgZMpH/qBpUQw368oxTdi142goOAw4ucdirkSBN8WYjZ8BuJqmj6Hz+CNI+8zRsmDhwf
9Ii+hZs9QEvzZgS2hDrYEPVinF2rG+IuVW/OmFPzUF/YdsG0whYbvCEBUbX27NdiT1sJR75+yx+U
Pz3f4KSlpfUh1Y2Pc6RpoLkTmxUj9PDD5xNMnNZcpJefMKKr5P/rmgjjjb6bksSK00nPDpcYp7aq
IxaQFneCh6y3pBoxQixNs3xWgxwqbCuGfKYpWsR813HgHrSgnJ54rnDVeLlWpsohUoS2qigIhamp
Nu/DV0x19+x7Brk/aoB1cIRxQUlUHrSybTGdjzl8ynp5xzkpMsdUZp1i6DaRnzo2/srCjzrb6fYg
+eeYyGKeag0hwDdcpVgQ7S60lE7hMzMq8BGKn0leW7wFai5+GtC4ALgRzPe2hSoXOi7Nh2/BO0QB
pkEdVtF4lWXiLn9KaYzTIEFUSaPuFOLogRgm9SOOba33pNdUjOJfyi1yGgVMvS+MLcBHrP65Sf9t
69KLlWtQQsq48Q//QnHEp5FCZkJcKgI5xhpSkwYb/LoI+gbor4nPQcaxg5xop08Ubrb0tQC/wf29
YVGEjS57BrbKqkrzoQTUOsao5FuMsHgk4A5loN5Qfg9iJVjKZhmqaRjYjmZb89qwtWjRsmc2Lp3j
h1pDdbJ+U/erxouPpvSCOeHKFxiZuGBStD91CnuIXMFKj9kEgiW6a6GbX0MHXFuOuCOLChXWtjnt
Mjz1qOXuK/T9aLvWNvQC4tRXueGhMuMUxdJz5PfQ6/Vl5HDjQrU/F2kT8bzOJ1Qh6/vGntUYj7v2
r6ucH2o0lb9vgiFj4VWadKaDQKT9Ub5ADXMpZHEMT5NHcM8cbaSsrFTapKtfpMhgn8xGe+EWUigt
/tuncpeaZXB1N7k8D2kxZsW0mH4jAlXl4wlWieDv1CFHnUf3/eakocsF8uoHppWt3BPVJPF7pr7Q
3SWyNVaGtlW4xEEWQVp7MAv3I9aYuHNnXA65X+Fu9fVotx0IJyizUrWn09CM1i1a1/0SDYh+z3pJ
yhYjy1hmxtMGtjcSxtpuRhusq9mxzxljrjuoYy1UYVfIViCbY8ToXQ+8g3zJmUiAOhVsVgR5sq7I
eql8d3Op/Ng9vroFxbr8yak6ftWC6bGu400KF3WHHdXvkJrIVD0qjVPNLRWF4OQz2V8dNC5cNq8R
9w2yojUBY2cEOM3ekOkIwDJjubeVB9gnEloidfqTBNWcAolrD5tP+50ShTtjOwfnV0NzrU9h3OaR
klafhX5iIGuNeE0rTHm3b5N2bBPx5J6wBYnyKPz4mXG33TfLfBghD/q4Il15GfgjEEkLGAXY6UXx
R2G2sXCtj73hTZ4dO9Qq+qyxN7QmBgPMP1Cx5nKsTHgXiDjcmugWf2XFiQrphMbtIzw06IPRft+8
VweNwUrIVq+HQQvPTYTiZNtcUlolz4LBUmaY7JUCpQOb2py2n8xtQn7+MEoFhHe5KAh90Rv9tMee
W6iQTWkdUtdL+2FJYqSSmyA0F53QsN3XGjrSy0jIBWiPTLYlTJbqZlqc116thizbkbpYNM/XWpVF
frORSCsP8DSnak3WPw6rxdkh6b0wXRkQGa8nx33N/Ckj8kWqItOe+g+y+k46uuZ/BhGnRWoOvS0e
MFAGI7Y/xX4qD5r+Gl30pUmQJGrlRwTO0jrlbhiUCPxgXPfx2Grl0pTG9+XBSIZ3zxO87xRpwxTB
OpmW3CzIie8m7GM46El1eUJa8cqI2dgDgHTNOMyk2pWxmAx0ORiHbWwwsHdoB3Y3FUO7HvJ0mxOF
WkwHCPz7Y7hE/8QD9ReGtoVqijHlrvcUW3XSsnZ4jsQiKUPHpipVSA7jRlTLmvoiy6gea0Y7/WV5
1NH/1Ys6PoPByTWK6QB6tK3CdutES2CxJIqk9sYCg1lZeYMeP8/7F9hzVfXJjqxfttL6Z4LIlB7B
1xV83XgRnf/B0/7TIV0ZEQdBYfnXyBucIK35swoTreq/t8iEUEYQAFS0xJriZyqhvm/k8RnhUrCb
RC7iYOYxiTYGn+0lrxHMcx1CZd6qlQUACFewRqP+/KP3dnVKdMbk6/Ysn3AVfeWbSzz+JXFTD04I
Vgg/rjLyA1Iz7mqwqCRI2ctnAhLsE0illDe2VnlOHnAxDQfLbcPMwY3OWX7jM5jB0z4TuU02jSs4
RSuakRv7+rlFMDBe+tW086WzwjT4FdtGMC0Y4Tu6gvxlKLOB4RfGRN/uaxnSLwERaNuWRk5Hs3fb
WOgLGon5Wv1zHp1SlhfWaZaaGY74kF4d+MCOqS6xth2MCH3iBR+aMNGes9AF5xxp0GP0EXxmB2pq
r8qNF1SjXjkSkcvDrDqpl01FPfwMy+cxxACDw1cArWURktCFOVW+ClrcK3W1pRA+QWoWct9aLT3T
NWk0ESMJ1AQDWmZdPz3Ij2hLInbr0cEDXV5k5vB6vf5L+iC5QzjLFODyfTZz2iSvx/jny0VY0MMP
7Q0zlYlxntoi684SCt6KOsyEPEhTCn/FX+Nf/cyXUK6OyjcqWuCHL+w3JuM+n7a7aoAEb4uxlxXQ
2BpJtRq/7PwxQ4pTy4vyH2NEbXJWn1wR91QYOQV4P5Pyclax8FSfauDfngvNyW2N+x3BCPMIHs0V
8dLNdETcyrfFFMlXH51TpFGsw0yoVEkNvAY+qz2bFJs/luXa1w9MYl//LiW5fbQX/YeMoV1WXdbA
IDtHVUs1IaDo3Me3b9ft5KRoTLpJRJRnVeEcbWP/TtmmgiODx8CEzIXNhPTx0gT451NhEdheWrjG
RTMjoPcsIVz73CjbrQrc1BCggaDVWf7aCFfbhEwVoM22hgyOVKOqCtZE4ZdC26Se7P9tYnnOvO2H
CmKp2eLjcfzpQ6742D2jpXxIPTMj00SXLYMeYt+HIIS8OHIf71Zn6q3g22oUXB2up0eK+quOuPtv
GDRxLCdR7a6LnRqLA4gYTPw+hLSfXQF82CbCgIWqH3sY3Vh1PfoNMbDdZUne9q14RVjfAhiy412h
lwPIth0J0DgHj8IPimJYM4ebBXltwjd9Q6K8G4nOMH4zPd9V8yJ4PZz6bTaTB5+aWBYywPqN97Lw
zD7kdDt88S9NVkD0S7D9ldA20J29FUiRGCtBmk2B94wFMO9ivKyyudlDVg0ZYJKPluTxpcZt9Sxz
D2F6gY0YUk+O4YMkhsmM1jWErTB2J5idm4WvFw588dMFZApU6tIGDKp3qCr/aD4saYy0s1jk4DK7
oHYA0o+Z49Sqi+7yCjC6AvpFAoznhi41govAdkDmhqNKkjzh1toU89wCHpgGSSYtT75G6pVxXQDb
4bpxkPpv1dedPoX1iYx3RtWc7ehYH27ejmtm86aaOgqPKFyZTP9YlYGiolgwJZCLzPKxzrHKZ5wp
awSZwzqMd5Xd74mrsDSdCz9+PGcA8071YXiH7vDWWmr5DJd/Wjl5H/t7hlRpDsmIMVZNeazJG+De
jSm5DbTaOTSS4rg2L2wZrHLBMkH/HPNFmXbXftFiz4kiTUNLxKrQ1VdvKNshXHRnpIzTwlR7GftM
fKdPMEO6VyKRkZuETnGlx1skXxNwrKpTIS5AS8EoPpLdkm4ZRCgWXlDdZnkYLeFwCzLVKK5jrIqm
ewlUW4/MdQcQOJT4IGrPTe4lKBoE4nxQ5pHkDLmgPdWeMxzdKh4mQkEX0mGwtyc4X0UyeMejRBqu
x2tHlvJA7wk/6h+hIY0fYOWWucu58j7tDaxJX0vEs9sINSFDOpCqpTGpMCujcH+Sn89xpoHZIXE8
5iFD0XLmziPiZSD6tgdkGsHKYyCcLi7e6xwDaqZLHnKcHR+nvyoENPNQOTgt8DB9apUQ1ius+6wA
QfdfzkA4CJj9M0vzPSE9UXhUkuATGlEaTIl3hXs5p+vbsbDL9DLq8shTQrFBTiMTvqqV4eIGe7vk
7AWYiE1wrJzVbW9s/vWuwxsvITwPXuhLhWCSgTdkQM0PQgeixrBvyeYh6BIxTPiVI8QrOSqSezxp
D+ECEKhBFqwiulop7l56s9dK1fa+k4v0FVd0XaqMHQptCHIEEdAz9K5aGvAsOAiDILed6k0YGMq3
ibQhaDTNiilKfOS2AJNWrHGWTgTQVlg1nxSohw3V+M2nce4sLKnI3tK54Sv55DtSiCufDqxbynXe
psw7aV2spWDKW3nMWvVsOJ/LfI9Ye1R/MH7dVBy50RzS/TEswV/MFeEZp3Hlk+KJpopyNoADeliu
bAnnw3reg474vT3xhPF/vJqMmuL4HVKFAf+I2AFSLXgi5QVwUYIjrjCMAeI9VjAj3mYOsmgNjY9z
VipDEoufqLqKiQHWgftQo1jzMfxMx3oPBbfT2SZptZIYFIeGl8Fn2PSGsdCxlAdGRofFkNoKHH6g
ok8xlacvami7EdFoQYF31PjQ8moXgCFe3t+ZZat0qH2VPaJbBmOCVwNUM4bF1xmw64IihtkK3C4J
fDS9xwDMSTEUyeVVaCF0QEurb5KM7YfreZqRuH0mdnU2MAnYh54KVUXcqhvjdwcPJPPT9NNsRpBT
J8eMhvY61riWCtLYb3JdwLAPyEN1FBamh1gJnxWll0SPHGP0xeDhx0v/jOv7EGT/ICgc4tanAgTz
JNy5SbB2rClEHhkfxufEDVUsOdHmYTwfYg074H2XrxNVSvXUvI2Pg4fiX2o5ujZZkzqgrJYlTP41
bbr9623ASQCpRta+ecZlu6bTPbr8Rf4iQtLwk01NOLCX8wVHri7F8+t8CunnAkyzJVEjDTtO39os
d5FihDgQFwLMbxzuv2Kel3bMDrhL2bOTD+KvBSuJa4XGcBW9a6yHfX1eW4+33xIiA0qJtX781NzA
a87f3OsYe07tU+LSSPWvKYAhTTm3hUqjHrutCNioDndY4RD6QsHhI/8CBsnb+uViCCEE4MD+ZVtm
sWgpH2g64vEo7jKvnIv27TnE7g42o9fB6Dh+fu5dL+FEzc/2wNR+YhXuN00WuLD63jawX0GqOLJA
4QzY1PovTG/lcHcankUqwy9XhTVfiGDfHvEo4VnMxTyQnsB8yzKasYZbgkowBbEwq6MkbYdrhHPG
4k2+2MiNKDW7ZaYOwDBLonCkseVT4CRw8/ynmgem3YNgJsuSJxGOhVl0x4vD8r2y4+StJT9B9T95
V8LdHH7oiluSG/GkKudlHRQgM26+IU7eSh6Mdtpa5h8Q29bGivX2CpejklHqO1C5e/RXZwXozMWK
CI6HAp68otUdy0aVLceerNz0QAMIAfOCeAfWCWuetyYJznX5TttzEjUmAmQicA5nMqQdcusgC7UI
iUNXNu4yc5nA5z0LXGfZIE2jZ7IXcWalnZrD89K+yDYCddVx+jZa6CTQ0aHJhWR01q25ULtMMg1w
aOQk1KSRbgCP1I2CXueJjZL0j1KkQiy4TGZi2CWx95jp3JUk1VP+Yx/eYWHQQRRJBD+NXiksPq+3
90+Pstdfgzg6AXjxMeZAHp9XHmYvts26scFIL/hu5wrIra5Meiol/9oWVTJaY8QakS9IX9UGg4hU
giI7RLLAKYXUHlzuG4vNmzJxBmpf4ZSRBPKa1EYgegkbf7JbleR7jIXCEsVaGUxMog6SBmqpsRHh
LXF1P1lfowkQdsiVH67FCfKsWHrSxREZ5/MCSf0sKqpxMqLfNsFk+lu7agtkar6dwXGL4Lozj9Pi
6HfKzjWiX0scZ7Vbu2s8Uv0HM04xL6wRFXqK6cxw1T1+Y4nh53jFT6PpxcRCp0kEJYF3TdlCxCwd
HeEhD9nxI6TzmCXg12hQx7YaFH2BnIUtAPTYFrTh7G7iOT0RUd80LRohAZzHODDo7b+DLB8/hYCx
Wn2ZvMI2Yjrqd1bGIqs0VhsCLJ4G184GLLzUpQkimHVzViYT9LRsG9Hb/ovz0Ha04iLRAocJTwcd
CvY1QDnGoi6hV8XaI8D560qEUqq+2wqfNym4YTQagme/uy0ZQJktzLUboS23FDTEFionq+n6RFiT
2VvxdQZMTIZFi5JraJk74pTK1dzrxdfuPlm1iv2t1v9zRUM1OfUTrSVcHOpICaTLiXsb4DpixdYJ
Fmr2gq4SCZYC7NMUCsidMuWhtEbmOKi0mu0Jz/Hz5Ej+ulxD1W5Y09kkcFvBDHppm6aLQTAc8Php
x07xlm1e7KGhOJh874bZbLPKjv++C41k5/JmKDmHGqPLez6F7v+kelGI+aeftXUMvv4vKegmYCdB
CjrtLvmamNsGLIl5eO5n7gx2NbaFzy5jymRQv5IbqtMzec974VaEK51e3YUboASertqhXjo+4WQi
ZNiDGln8+kEyMHAqRui6P88YCzFTZiNwrMMQsswE5mpJiQmYEymEdyNBdRTCmzspZw71j24AyOQx
aIIqg390eqYNQOCzkegdHsfxZSJ1gKr+AK6854wcmXLV69Zm/SaAE8PrlVww69f5Ye+SCR0R6dr5
oT2B8HI7Nvbz+qoBaSu05SF73IHBdv+/xVrevo2Qu9HfmP0qTL7yLbDjAA/NItGxszw0JmCdEZf9
+9tGpZcwkjJj5NgBHotYYHRH0xLCSNPTPQJbDsLtYWIvKZno7eYHdLZPGRw5RQCMd7FDfa+JtZoJ
ik7wLE+U/9EhiAcypAwTG5Dj9hodnbm+lSxko6ddV5uhBt4mzR1JZXBUbaZtwvU7axoZBndpYW9Z
51+oHERACwYtQ1J09d35SBcImj/34gG7V3qcFzIrmugpftkVmbgIxNaW05vQYOF+VEJreGpquTnZ
9WBzz3DvnDhL7DrDG/TyEx9msb93NVBc6RNV+vVO4FpeLRY7bnwhFGXvNBSq9hpDbwzr0iUOLlWq
WKvJOGCTFMz4TpuodrNUO2ohP5w6QXTDhjnniNtJa1hBzVLF4NYMvaCQZ2UmRPIh6sPsxlTR0CVQ
R+iAyGNO0V3wUGG4pxPZwOBQkUcTpmh/tRmsZ+4IZ3Ggn5onsbg+VuHoKEcXyy/e1oe24yp/z1fF
WP1LPsSYjx/DSS4VSz4t07GgCct8kb97ztOQTE8Qwei1YwnqYZpeOSsDDHZWXtRLXgWRs7e/BQTF
Az1lMMOkXrrzPOyNqbhqDHomaeICFti8UfQJBxzMzJdY0oksfLUfpfHzATr8dG3+QaaZOB1rLspo
xgUgconDR/gdpv0uvI4Ppjw1ltWLxK25yyCr5xlFGCdU16cCSYA8dJz2nOBXv49wQ54ETJYwTjCp
LLJ0HIp5SO073LLB0Ta1/oKtDBJyHiC5OlqATJHEtzLuxkPKgIIHnV5wzRBWCUVApYJUt9VlxOIb
T5iC2EY2XdlQIIKtUnmDPKyXq1KIJqmMmdCo8kLKYwLMvjaqzmY/O8XBWpDCdeeMlA3/f8gRUu2x
aEpVOIMyOB3BSPKfQOH2BMTxgJYojq+nHM8lhweUTqBfI7v86L3snMCEOOURfSny4Xr6lVICJHZW
+OAC3zZ4+x5SSekGYxlmvUjr5gVIFLcCZ8K/gN1Bdt5X+SCbOTSnCGgVRTgNsK03JMb0wycHwRSB
UpZ//CHQKX3/Z3ytC6M4fNQU4zNdMom0JmiOnegCVCJip8gf6+4CkU78riYLD18VOuQsTPqlMfGX
GpbTLFizjTgRttz0NgKFkfKtd2qreYHplyrKglFCdQMmCagwK68J58Wcp0TS4SDStEMlFrAKhC+u
916ipl7In2iHa48eqqVYeiyHTmq27Qv2eEgmYyntt2Zyy+BkjHOR5mI7Xgn2VIJ0qqD3iGs0pzLr
Q53X1EcLkICA7OejDtq2j/6YSf23HpUBVxi0wTtg0Q4VSEbhHwiXcAagIUZ1WrqEQY9+ZkXZVeG4
g6S6DG/zYPVXh577w/lmBPmF5ohxSlZd3+biCaMbNF1+/yb52i11RXvDlQjfBw5f3HkkQi0CE/0h
k9/aD3VHf2axPgs7j2+aqLU8HsPWzydrYijU+ZVsccB3q65Hq+JE00ldt9qna1upDQYN8m26pRKE
gvAQJrbRwXkYXntNpuWMs1etmmIWAbnrD7NoufA794IXNIF+pT14RmLs/Fe/6RkR19uMf20FFlRw
d+upk6DOa/9NA2w2dm16RpQ3rO+BO2LjI3StZSwRKxqPD19wlG+/y93Lov4DGpgRsgwkWeXhA8Kz
i7xq/9bGuA25+ccio0w5+JOv3MNMB6tsIsD4wwfYLjjD2SaPdEFKCMidHbAOTd3/nWZ0/N8+E+HQ
iSyAJlcF4o+B8i5g6Deqr9aHIsQ4PpaE37SqrXqQ7boAXFY9satX8FUnC1BCpv7PssZi6U+h1TSw
sU8+mddDyFuQ2HXKBtBNYAaEi8DkTnMgxsKodIs2QFQ/DEwAAjYqvBr0NpsunzCDqEtjdUiw4K0u
SjyXwa3re4W5j1u+gsUmqCUpuE/ZpN8KLk3gEPYV9zQbs2OpEDcl2tcS7oB4sIjtzpbxnz97bwAZ
mdHUj/EhnFLCnOBsvHFYrBs07kghDOtsZhTZ1czKuvP9IeRaRTweckcDoZ5U3uki8+B6Mzc/TRIu
rsz/04sFVD2IR0gMML6hUO1qsbjlHnrHqJgQl0K26PIgMrcWGTc7zAV9R4KHc+Ix9spwdvHLa119
ETe7j+VuCsWQfyqTKhLwDvSHlpujQTiT/KqXw346Sdlipmw87SLLxuTOLOWMbpmLwyP+BSZGURcD
DkvoF6xRHKr41WYi2RsZFMfb6VKeGaWOtHuSIWGxmjhw7WxA6N3pfQb2xK5JE0bT+5I9eIJ0YW3T
mVhUrIGlfOz0Nf4iDAi0J2rKahYpyONXrPBN1wfajN3PQP/ijy/drwxCB6IXpWriSz1IJfTClTFb
LgZR8knS0HcvLPlCbrUdOUPlJvCtUnlUQul9NmFnfq2JG11sJDuVEEVQzOOA9gLuvHlGXSHGpIxt
ysY/ekbs7KYSFZ2rk02RvI3fVxCxX2t1JEQy3U7KeYIia1MeXeTBGk+wV3C+q+N+O36rJcole9YO
a3w0qwpIw9UreRO6HIYcP/c0j57SOz6Yoj9N6Thg7SU3DwfrLRwgLnZl1zzWO28vaVAoMShm5FHm
IjUYqDQTXys3nx3MfZmWxLmZo5AJNImVzVvAKtiMrc+v6nuCumWlZ+fW61KTpiCSk2D1Fcmj/gOQ
dFuzfdcxbPKe4M7q/+yqhYhJORISWDEcPAMmmEcV2jVsjdh9I77W6PNFfHOS1GevXqjW50bA8FMM
5/vTYIK77juW4zhxxHs7g6WY3GPE83jbiisFvAwtKgNyfvdotGSoNRWCbg0f4wgf/npxNkDTA3Wc
9q9iVVrasP9MN5XEs5ptKEXcpNfTR4/6ERtQRMuTtdXWcpg+JlYF3Pp2myPneM2xUbFUNBAip9Wk
2G11iuzJ/gUf1nQt6QW1cxURL4/0RUcZgKQ1poz8/nqfJ6ruH2nqgKutaIro7u3RqqjkYRDkITw6
qoywijNkAhRQj6X6J5vxPkYm5vH0k17Scc4jDS3N0P6qk74bE9/DY4r/2tZfQBzWMe41i1Dy5+LZ
z7euMG7a3dIMjO3Z2EsdJoUx+4jLtm0DoG625kbkK+96Tkqmzaeda+tS+8pmEULWLbAgB7RldQO6
U9Uv436YaiNldDxcggFxMuj4fFvMp4BI+qWd+uUGy8NNHa8pjem1w2r2M/ZFp1WtGp4/Fq/iQedq
2USMCjeJ6W2Fo6xgI4nwr9pK+Vx1sK0y2aAUT95LU5J56PaqoehkKJhYUeUOscO6KNwPQ9Pjn5N3
jV2ieT55yd6PeSeXuwlBkW01iM+7eoxNF7rI52xOy2lcdQlxl91wI5YSdJXpl778H5Bsn/wIK5ox
VTcZcWNqxZ+WW/O8bld4yycNJ0ND9ByTXKondDglmCZESfKgrhf6Nwb6E3Eish0O27ft3eJwEDh3
ggxkrzuXW+azxthKH8WGVG5olwoJZDSOJBT1MOlst23E3DBnCb34pzCzRmzQf3G1JA4lqF29u0Qq
Sv2BrL4ht7D4yxwWCSxv/bkRPcGYeVqtWQFKKNN9JGVQVoq8SkWCaAoQFKJbWixMEj+8Z3OTqdnQ
uat1IVZvwYTGwTOif3bB02cciAAIp513NqKU8geohyJLTZJEvBX2AMExFc4x/k7Afltb5D7OJVnS
L2hpXuid7LyizbEpKGuYBj1DfoTx1ayz/D+EhknrO4rfiO+DWzCwWFbQfAQb1ZIDMAZzJBEM5iOU
rczKMb0X+PAzmPjxVCi3CQPrWKN3QC1yAYVcSEjIAW2NvH1lJTR3NdCPZcQfNbFPHE55mE/OrHR+
kdb9aq6UuQnJccvQXA9oHcMsNCXXsq4Po4s2a2z0adSuRLOIaAwb2Aezz/0Q47Cfh3ZDFrbBfeUN
198n14Ci/FDyN32WVh1J+DDENjtB/yCibcw+IeNr7ufkWg5qlvio9ln+ON4ehI3nDc1jVTyo/qi+
1CFTChPF4RBR7GUruUjXFmdJI2z0uTfTz6prtmeiphwiBdrWXsj+5+7Zu14cDYZrW5yRZnryJPKk
ec7NIraN8bZymCGwW4g6u8a4vbnIpKpURLYrw6fL6P7EsVBtLoy413tIl/OORp3a7ogXdNIH53Bv
bjpXS7yCT8AthvbixSei2+thHN/HaeGqiq4MOSLz897lRcukumg+sjz3mOYgW9SyKAAFtpZ0Uy/1
VdasIReOSW3Uap/SjIF9Iuu7TJNRn3klBUMYbN2cXgjuVUm9tfrebBEayvigQDKo7QCBKFmk1mSh
Z/3/ZMEWamWpC8TV+QPIY1TtocfCU9FgRHzrfUwxnqDXnl8pui9HqyJGUGTDEq3hj/GsUM1dspDb
6QqpIkYdKPCVpIekKb+pl39rYaItqe7HkNGY0lcZUSLJhIGzc3q+nLP+oO8hVQiKI4SVFRtwDptX
VObmqI/x8S4d7wNj5Xbv220ISmxw+eJ4BKIk+R89Gzg4tG6uN+XzGBSiGnemYodyYy24kAnmbjIE
isJPPzs7waKM39yG3F3gMJ/E9Z8DtvVOYKzh9GKqyPXxtqchV8M616czf142493a6AXr0ldkIa1o
KCeILIfYn7ykWtpcSe8GUGujn6rJHVxFo8nxJT/2MEkorK+yoUEhJfpe0SsvnFDXhXw09QfoF06a
xo/5HpEg74IU+2Ia0bqi3BHBnG55zztkinrOQMjGa8NcwTUY2HkRIX6XHtq/xjp1NViQco3W8EVp
okauUo+7/+CtWaJNEbXqXUwMfyzC/Y5hqKsH/UjVG9BLfcIrVxm79jVwclpd8lXdWqFXUCJmC1f5
teVbLAQlhvNmfiaRm8wxDCtfOjVPOWMwCqsaMC4lCaeVUqncP82qC0hJ2rN5O06Lv8STDKxtEM0R
eovEhiZJr+EP6ZMqQh0NVMFFqhaF08vNdSLWYbwtozTEp2pY+RY21Rq87f/wXOOD25Hul/SEbNOe
oEN30CM+jCPSaMFFc2YTvmjW29F78+Z8KaacpXsLRo3hOqb1y76Xprk/KR9r2ut0VDvNZa0X7IPP
U8srKuw9/bUwqNaivOed93BWUJp99YTelHgjc9GQWeAQRMOZkRgwTRQ7CYNjrnjzRY3fCE5Ck9jL
L6wnvn2u2XEo2K2Fxs1NiAQ59JXglBbKoqqkTQdqvmp3XsNNsGgpyvOm5dpjR76hBq0pH40tSwqS
/cVXQS2vcJyoba+2TgomDJmHipWP9nnq8fMldLu3nqZJQ0hledM3nwGWap05pGy+08jVVCfiE2/r
s+t/Hb2h8eUCsRY35W5+ZeXJN1DIvgs86iG4s3R9XTRjLmswRPQZEr3djVXtaxxV8fX8Y8uEEB9T
ptu9AFlEsw79Rrdz4nLPyFYMie9AxyyYT9i1CZOb+b2FUNjyVhSqhJy7zs2ukHQaZ+V32nJgkzGq
tLQBaDhYm5AEhOHSms6/eXk732sOHyrrYSgFGqJtZUecYXz1mK4hgJcGrvVs/jvKhLJbiUxvLYnk
paUDJG2pyaMqJOQ8CQHKqhZ7bg1TZiiABJO6gc1ehMHk5MdL+4uh/5TXE11B56a9L4d3XDM2eBUK
FsbawyyycZHu9BcVWEp7b0O5s4QosaNCZypMHm7T59Z9KK3gGhTQE8hHjFcAf/IuNI0/pwFFe+QP
SGQd4u0CCDLFANyR0Soh1MmyjQXLIvl2Dnrly8G24GjCT4fc0kwNxEgdwpF4Y92/rFEJVOV3V3b+
7ITQo3cSvwfJm49p+3EOMZAyhwM9ko8wjFX8ppvW8tBgKbG9wcShRCUFVIlIh6fZSnYWsVJ6rhNH
x9+pAS9x9k4x+FMcFosyZ6L7ZH9LNN+3Nwq0/o3ySxhSk94PmKUpD1I0jHsqxUMcb3lp96npz7vk
vlPVIyrYFb0kirV0ZWjINvrr6p4d2mui4FGotKIVctVbfP57veetQ/4kJfkEAHFUTW7cAf3CqMEA
HR0vGXh3DP9kWtVkg//6aCw+EZiidDJPJ3lQ00W4Lp5AYOKyf+NoD6EWltnsOFVHSUpPU5AIAU4H
Lz1gLyLsX+6qVcp+hCtqsrhw1RM3em5ZAEBr/dwJMDRmOIDCem9nDPvusiFmCMsEWYC7QAeZjKL+
PSmDew0UGL1PRlcHZwkGYIOM0CJLxW8NZ5u8S0oex/SHMyF6eDMaOeGhOMVI6GZrfIVIaN50Fclr
olitqABJMbTKEbfqa1rFvOLCcHA5YTO/xk453bGij1w6xBpT3FtDRLxkdu9p3kRfHQ8FZOGNkx9h
+9clFgjQe51ZQ7linBL4xt9thpqxLTn8J8hLHj6V13yaImJdyGTEi2fXW4V7Qd2LBmByXuMU34Na
x8j7XyIMN4Bx+cpCMC6Jg1upvcxkCB06BGL75uDku75Lf5UFpgfCQppcWoEfyr9LaHMTnbaOVDTw
moBYGjRoT76WFQrF7bDx44a7ipFTa2lTBqsMrS3gN1Mf79u4kAB99wjea6QzmbTnw9YIcUpRwqTo
OsWaaGdlQHy9j5JabjPfgyn1z+JhGjH2paZgxslilkn19QHqpq2EwjVKrO9t84AvaeL0FS3wVJwb
1PWN/Kc9j/7AhVAt94/yke5H+MkHrbiTXFp+dWt1iHRP7KV9KGJ2xm5DWksTV6CfmR6zH25dKDjs
7uFoQV6iG5UL12r2yAyIPxt9+L0Z9RmIW1cbRzwvESpkWhATlagHkY8SrPrEH5kVm5YWi1cxkEJh
nSFAwN1EJfKgBlfhC7dSV28tJ7Wzekh6cJQg/kQwQWGR2++soJBzyZgZW29yHALnC5HDnjciyo6P
HWjEoV3cVv3OJiQalvKudrR77MmrOR8/2wAt3PYRyFYZMoNO1LYroWSDaTsQZKcTE0J4mf0K6zWu
KO1LBNdNhkmTR/2g2Fl+goZycas53LAxx2HWAzSvQqplUvoen229vGfu/i5U5UkSe8F0KjkzM85y
F7esdUNx29WiDDlbtpkQFt8q45Ibwyi7yUQdxhCEuT5hHqj0UXuZXjUfhZCWxUTTHqZ1ImMWkn8L
FAb36GJlz+PpwkuVQX09BonjDV/zOrc/L06sPyOJUCEuLXL2exggeFJ3Z6EViioEPL97NXU/Cl3T
VywGNhN1sTDbexI9LTzqHwY1nt2arCT2cCUSrLOvTaTSBUVf3IP7AU9x1mAJIWTSM869w4r5Eg5p
Yajfgpn/d36nB+uRb8kU88UpWIryTmX6REsYqXTVN2tszQKhHBISbWNaOpQ8YgfjOwa4vnKbT3CL
1OlF59GPw/KYoxeJ6G0R6FJdYEzLMaQJBUkz4fvuLmrVwUsbfyo5ES7A3NlDTeGBwSupgcvlKF2U
megvWIJU/7trKyGwsa66WYfh6Can8/FIx9MSfoxtkTj+rwgZMH0eaDVnQQLowv3eHd61Ep0nblG7
H6oUO1gIzxqI3vjxKlAAYrLqPtmS8XLBu0ksWJXV+WXskL2A2bh6E+xKV9XJWFtS1Ipd8Esf9aPa
267JbzZC308S2x1ANXQRY5Fc8TyhaD+C/zLgdZDmf9H0HYrIlpoFSpNpmhes7wp+FO2WNoBalu9i
CBeMRT9tPF5Ong8Wx0bNuz8En8Gv86G2LA+PQkgWZXllDUySQjJf2IxyE/zbtrCKEsvRXXEH6Iyp
kp6wb86e4BQ4YcSANBzzKI0n1Jw94SL2CdCVQ4ICuUVp1CN51Nwb1Fsd26Z9MwtO2S5yt7b/O5g2
OKgx6NSJkEUPjyQWaJPISah1fXdou2bhPc91hhtOTumRPYNaKp8bHbX5uO/4winereyQEVtccQzv
Rz+XBUOSR5GW5J5D1KoHQG3rusCHiGBtlu4tZ1DIrnfpJQ6PllBIhnV7aZFc7eU9QJ3zowofXeqF
VXjJ0noj5Z3/Y2icFIOhQ+amGvBWVEnpPJlDW/jsbEyNw9ihlBIpy/HroadDLjj/B/cr1lYEPsQJ
HubuJrJam3AF3BMk+amxW8Ud/QDNWNVyHbU+042iED4h9lDEk7wMQQYVWNT2C2rqYAn23tROFNi4
5Fl0fsRuGpV8Tt1o+ivYkJ3XYN0JxZg0Vd2eedyYjIBqAjnVcPHY8cs+t2vsul3vIrWn8E98asYK
MxFWCV0Bqav5jWZ6gvvQ8qg0l5KsxAp+PMJUPqKgnF/N8yUsQI9QbmKUF74Skd4MUmPoR7kyVImi
iWJhtXut7Kvg1j5CbCUl7xsvKo3OamLc4hpmOKtZlQRAus92IHGz3ASXO/aiHD4kRf1UJtXYMjp8
Dk+ZjuY588kEd72ZhnJTopZ+PIYPTMWiWtVf28p/yvmW6vGQxYo/oRo4hxdtrCI7ROIDWrH9pCDR
KLrCkD9w5rW4DdC15GYHVU2keTwtvC/AER7zH7Wll86mLcM0Gmc0QS/fGf4NrLVq2X3Duq3eQ4pr
JBf60Gq12rfCxYtEMkK+nx1+7YNuwCrBJGQHertU01pbUU0Bldfp7Kn1ug4PfjrZnVpnuezFSLHZ
h3iCbOEjf+7JYtrf5hOLz1FwlfyqUkxVcIbM+Y8hrB2Kfpn6T+b9yN4UqNb2mHvH8pWaVUKzXdA9
Yn3zRzYda0fLjrxPNleXRcGt9wlRiegXnTTrOQg1gzn/30nlcz2PLiCHeH1wWgox/ltH+PuafP7m
fzXz5STspCsxM+b7r3lWmQ2eiSQ+Ed6yaI/pwJNjCwfzb6ZxWtWoyBg8xsQSnRgYIy0bTT6XFJ9D
bMS08pk9Xc5NGdkGW7CfHg0BlQX7UxD1lFSAE4KBbaE6MvkLUZCkHNejo2mbg7yUzv//BWkCnC7D
kfNqxg7qY7GN7OXGBNPaL6V+mmGZX15Ems/MfPVDwq6vC5wmS1au4c9EZKiky+pphcgaPdjmhf2W
6rd+5est2c2WMB710X0DcuimpirUEzKQF8r/r866m0HPhWQqlhdQnhkk6Mwys5s6fw9ze1PP2O0l
OwTXSZXKSZznkETYekd38ecSt9a05lKjR8j/nRqdYajlNW80pByZh+FiEe7JFb+kPB5KzVBvLvGd
updMapQtJB0rwK7N51hiGu0hWUsYRG1i5M2N5vK62yRJ9nvURUITe/4iZWi7JTzAKILZ0XgptXje
D6ETv3SvnCLGvPRK7Icv0g/LS1ekz80bLtopIRTBP8FXBXXldX/rwbUuH3A61oXSdyUgYEH9viDA
ibLJ4anZcAPQHWmIGVkCEeUG9Tfss4p8MOIvUwOCxz4ATGzwlCO16ToclTSqQKi5SY9VEMXO1MNE
Zvb70kWgJBhYLuybXEeElpx1+sNuX224RxFBrJUd5wTcS0MG7k0NT147QKuWU2pzkyGoFC6w2t8G
YxQoYSzgt3xSGlc7IDx2XKB6FAIb7Ip3TqBTiKno4uA6lueDAkDstuFe3cWTzWAXEiqchnmtXZvL
ANojZOjFUEVBnAvITKtJFOgGasOcdR4TPWpXONErAXWptiElkzKzFPZDiIHNfbrjEQtFXF3dHJp3
Ku21HolspYyblenJusu/9J3mDzPzpCylYPEDIJfTbijbOhlc7C5tYpGTUsHunXh8fZjWlPTdXSRk
CO7K+bFRHAIMAPFra6EDw2JoCAnfD8V9C1Qgd4B9RVjavhc1iLnkTtDrXnVrY90XeFc5sA3G7i9S
IMyfZCVT6yEwhWrnUtq5XpMPxIbe7c6T2t7rk9asQhR2g6wtjN3ATp7UFGm8dMcgON1XHtj4o3AF
dn48s7TROB3b7tKoHA9In/9lT5V4Bczif3SnYLorO4urn74iJPRZTS6IXZevEG5maCaEZobdEASa
9XvPE8s0j3KH18FFwdu9ylGb7Saq39rKcZHQ742xu0qwi5nr4YRasFW2ajVW3j2KZADN7/HIEoxK
QYO0djNwiZPHIkxiAAzbka/YQypzxtaz8P3z7YZIujx9p4VBsi1rYspjyONrkVrWSaHDGS2XFBk+
ar3pamLECR7XMalq5gfxSkTUiczzsbtPGYEUMhKk2D7uPXz7svCizocK3UWIRdFzo6LeIAPHm9af
7RLTOaQ6uX/+Kl/25zvL1+oxqnPLbQGgYf2X6KEuRO8Mlsl5hYcSqwSeH8efqwXdn36w2zWMkSWY
rf1T+K2gVOnaqJ+nKD9Ee6Z9uvJwUH9cTr6OOO8XH/dIRtxEUmmblcdrKl0rgnRj+beBoRdCsEuL
dFomTVux4fqV3tIXBniXkHMZXPbTHFAS26Ag95zIHBOI1PazTiPhyCzXxJmoQDSwXLYoDSfGI1+v
FAugGgxdfi5AgQYnrwQcCBG8fMWcYD8ku4KXLKMBQZM1n7wObkU3Y7R9uT+yJctnfzDCme7ncYOc
U+flZ1LESVL/hzBWBOtuilaFJ6zkK9QaupP8gyFky6RbW5i7g0wU9+w9YGHfcBce1DRju/zT3LHR
ksTdjC3Ir3WSFY3RoHPX16Lau/X9bHWerPhnAB7Xzu9AlG+Y1LWTzF035TyHiG6Oie0GLTNmZ+yI
1KQ8LgN9kyvG+e+eJvqZC0+7QpRFXaPCCtV3dQ9NBOyyGjO82/4u4PZricmKxUp4ZE/aTFXwXGap
R4jpEqYs4i40mOB1G/qpbg6WAjaEmoP2CveFTI3oDGaKpB4pIjLysoHlTlSlUGDzHmWwom88ULJs
zncJ5h1PcXOoSP7jnAFXmsKqYoO4CvjVML58IKyJJXJJqJ3JJ/L1fqJDseIJz74pXEJ8j5MSEY4u
IClG0JUIT6SwbTV3dBunbNDpPMNUbCKn6UBmvj3YBzw6yk1hzFc/0k4Vas0HA6UD4OTRwkK6BiLX
BBwNZU4yLuQdbZwwytWjMn/R/MLuBS8hn6kVAmJmwvIiFQiRaQME4zJUNlwU/u1V3srybiicbh/j
TY/AtWYQCcbIgLHx6+KS+u8NCldN9JLWsdiqxFhv4ny6Yf5sw/PHooED0327VrUsODwu/YfqkrHA
2fDtaQXl2HnJJFHiaKeWmw0UamK7sPUfwc3YCDgL368wA/z3roTnmPV4+0wfaG12sIR6BcjoNBHT
x+itn9sXVKHTvkiZqKs0Lm0WlGuC0Xs67vMHPbOrD7XHGAwl2LYiW9ezRudUP0MDj1i7BnOqkKVl
+hhJtIyuPrtrQrF2eLZHwUm8/+NLEDx5ZWLmFVQqmJpbycRDb6YownhaHsx4oJzWT/gPKRAfvXJX
Y/N5avC4PNJqq47EZEDURuaqv1OLimWxB/yo4HvIA6Zna+3BlQdQh2WTaT/56T/kmg4nXdAX7Cxi
SgCxfUv7z2e9vA+5UocTYsx+7FlBw1R0qJqtAarhsYOVy4J2JZZ/M6R4Z0eSUxhZi4ImKIQ16lKy
E2eSZHhUz8/C2HcVn+GBBHFw1p4IrZ91TgNFKDQrtwRO7NJWY1oHtiHFDSIEvngchrIezL76UIUc
M/7plrVAXMrS7oyGnwdYeR31O+Sv5f6UwsMaogoz1wuJQZVGOGd6fmbtFQuHPiZtNTyMGXseHGjh
TtULfjemg0lIl4EVJmhHZRS/5v4EKhgJY/2X9l3bxq9uxadPi2OujEZlpLs8vVqOY1Jp6pMdGDUo
Qh/eL4CCDn3C6b0twfQ+5jZDl10GByC9EyMUfRlSnVl9oeLkW9bqz343GJ0+qd0OO/zxpughWIMl
2Me9CtYJ5pH6vEx75Cl3DJZ9n0s+9mEzzHOqAtOTXp623Wx8dUIVSFrj9Q+mygp0MgzXGpgwb3MA
lkBKJq0vJU5hyosUgx7fNMt0jo7Q+8EBeM7In6E/eupGKNSjCCOEV90iAZko9xdYC8v4JtWN2oYR
IGytxali+HvvHJQBNBJeLSnkviiG9FZxJiwNH56FPVk9A1ZOqJ7qTA7oOqhKveF6Vx61MqUBBk7I
9ggGm4+ZpIoUi7C9DHBc0o/rI0O5wdM746SXEC/RAiXKUPNH2uSJSxBphY7evaZBPRcpPFpzrxOp
upA4aPtMPB6WPZCaUbRpmJ83SNOkOARmByGbVySikZcSy/7QnYXQtZkkG4TzqGylPZzOwMr97gPX
hBSLXhYRPjcLRU0tTQs0qKSVWu6e+U6jbJALx6xm6IMxIqYc8FI+A0/xeHpPKYD3Z/bf12NOAYal
qWBaFJKqRRBLQGJexFJeIarmmVicxnsCcBgmqH/Rki3EYlZ6dcfNYObntQScOoDKiZ0QUi6wqAeZ
llBzvcQtCC5hoejoa7ObOlHDT4mO8ZTEMTa1wFHtDIDtmuL7FHgog9zTHlXE3yixELLOvUI1Gtqc
FNVPST4e3ukbf3Ri+1q6s0Ttaq6VVCyy/mV7V18NfqBtNsEQB4YZcWpkMJrRDXFvwLjKtJeHVmMj
JYYA+/d2DV9rQH2JZqSUWgaiWvaqpFG61yBwWygmsRnlGQGcL4mL4ZeWO+bgGs8pdGEO4r29UEKK
FMY7QJyTsk2NP7eIChxNi2lGTNIxEDjUgb8cnoFwb8oz+HTYT4LmSaRp7uWaoGj4dSNwzdMuJ/iE
fwn0zblWhLRs2tQeg1FMWtgGY2nShtPv2ldJPDfMYtmPtS5kcnYsJ02xexbtMa/QfT6LAiO6P+Ih
a0vSwCAc6WlMcKM4JJg77XyfMcSC0MJ8ajcK2hzv+Ggp7nki6VE0fHIpAcTtQ7VwqlBMC/rz1dzP
8cQJfLD7aiKzTmcFWQAtt0N1aTb2QQsk4HhsoB1ufF41wIOHwmMuh5DUnnz5B7MZWZFLfJO8ggxJ
jhWhKc1fzmXqT1AqmvXdrnHyvUC4+e8PNi/lDF2Ix/BQu+6MZtwjYaSUC333NJX/fhcBfIIjUTlB
pVnrH79iEa3y8geEQT2QjrXQCR3EeuynCqxcZ/7nKmIpxo0fhBwO4s6TWALKgxoVKh0b82iDfaXY
XejEAa1Tdi0PrIYYxbZliBqhRsWhNZHwxHuOsZFYZSfOy8hz7JblHpqupOYhuvMLlJsQH2/hkka0
dLXY5bYkLn+PdepglpcaOSke2mMz4kvUOSL+i0nRvNCEqYvVoRPFB6/OcLVe9Hr5UBLBxklkQcOx
uqWPYboj+CfN95veiM7XjjZYEtJfOGhxieLz6T6cd4XKPmXsygm6IntmCRSNjFG7R5seBn7xLNuZ
QSIcVL2ghlK8qJ4Qn0TWL5YNM0v8s42vLoId7ZM2p7r4dUICCpYyofDII7j1WcaD3xQf5OHzlBa+
FtbqToMg/U9d91wdwlbkd+Z3fLKG3YSOmYE/xCashojQ8UYmMlQMQRARs5YQmyH6yac2wHH6rDp1
i3OeJFQ+luFGJLqlaY7b4wgx4v+qc2mDHqSt0olJHE5MstNCBfP6iYwJ6kIpTiUKZSa/cDPenQ8a
flOjH4cqrJJxzba4/M6zQuboDzfuzC1of65YFejhjxSSIcZnK5fcSPU0Q1ZIrpAJqQ9IkI9gTOvW
nVD7f7aHuoCh6aVFZyCZIzxUcgY+aD7rs/5Rv/bfZ4EuQQI20+Uq4ZlPRlrR6wXK4aO1IJqmnQWp
uwad0kfsVXXNn0evXeF1O2JutNAq57FoOqgjqYntUp0jxlIjHwBC1JwG2zGoldT6oMGdOp3b0Gld
StDqomHkMRFHtCbWpWFwjZ5Jg2A0ipP6Cx7uiSZIZ+d3+YVEinq/oD/o78z9H8c+XQt+rFBgTait
NDIdzAqOuo46ZTj/B7H4sdvAqU1tdhNDp8i6Q0E2F26m7w/dEGk7smRqdRifHYp7Mtwu2u6gIsjd
OU4EnvPmYTonj35Mu9r5FH85BVuDXKoAAhhBI13sCHZfXJpHyMK0mrsf9dC632RlD8Y/ERPkkZ64
/tu4AWkjTHRgB9yxhdeOopUvNM21yiwPsYOpar9BjBGT1TYnw2VxMHqTE6GSoqzPS0tRlMWB112w
+6XdwC3/tqbrIs4ksKhVX7Czgf0KQT1URnPBnGEqcScVwdOvXxitk4wA+SzUumUi9bbOeOwilzL7
wDfHUV8ll4verbGBCRb8jN47bQbZc7EdJOt1DNJcbw8R9cYugP2+tUGJfmZMfFLCtGKBdL7akBtH
ACt4l3R0zM/PjKZRVXhWxobccaVtuLOaVIAGkPYkjBTmq2xB4YBD0qRwyA8cxxwSzymUF5y1BmfM
Ji7OtbpxlnRVh22wtlqqP9LXyPxcNYPMzCO4a9ON9fSLFAZqqUukOipUOAIx5HSmybqRzySLK+0L
QLlrmoxAiZI0JrWceTyMr4Rl7sCJFXExPZAfz1/1NkRYl1Niz4BPc2kOdJnJPzhQJwVJJSN8Y1RM
V0CK1+Lz/vka0Ij2n1UYd0QBy8zpBctDp+N21i/SUPbTL/yzxrjRW9gHleiom5wbEva/dCOUHCqY
RD9t4JuWr9fmxumQED4dEgIaw78Qo0uzrmS8NPAOS3boOKGYkXUw6hpcEFGyAAeKH0fZrzgFy7rN
4QzizvpqTh0xHanyxVLBRQJWDoiSH3+UjDDATQf6Rb70Q1gnF2c1dqARg0yddO3yVjaUv7/A58rH
wtuPHzOI2oRSSrdub4RJOdwWo90WBA84D+yazwbxjuEdz8yl+gOhZGQ+lzxZPeSfj7d4XtxnqThO
+drnutV08dNF1znxutllVfvVPHXixUbWjcIDYplW3OEw1JxjKmQHjfbBIRGbDAJKxDvG3Lsd7dw6
uw5Gbz5CjhagRKkGbIBFDriJVtnvLFowYysfORZqtsElXI9e8fHKCw5qM8KGVyTBS/Epx5YGEd7B
lqXhqAHy5vCAY+EQbnc56AUiIpkU7h0TGlviEz9p/wBS+sto/zh77bfqYrJJ9cs98qkVYBlPV5L7
3sCGR1nLe72snWIJ5iydezCPEtBIbPSzobydT8TzP2ktTJ2n0mt6jC1/Z12Vim+11kZL37oPyq/r
mKfFNkvDiX4EbX54zheOPr8UECnArUfjmH+gpjzqIn1vuhofWbbb5sroPJJzlNLG6wcd9rPtfs+M
XRBmtDBokdfkP9lnX54KnXDmyhTcG2pIsPRUgVyqq16uCW9iV1uqyhwW7whPODXllDpaVj0e9cYN
51Q+RHniFAVMyJM/yFQHYKH0hGoRsHT2BteHHEm908A2TYrVZpgss4yxkFPp/OoxyAaQqMb9tNhr
fYMY59bwMoEO1E8L2cXkvZtBMkadbTzeTivxUXOp6XNzttELPzQ2rSa/XGYxbRURYsDKxzrTuX7u
pGVSur8CTa69HsugELG4CS3Qe3CN1YK7I5j8/sw2Z6U+yHZqJW38VX/qwIXTqLSMspXp3R6YkyC7
V+TgVu84Ld6HnowKnR62fgem7yjIEgCJ9w3kZu7BOhvzSXnNXYPg3OPf7/rOjvU4UuWsbS8CM6bV
kxBhR6NHuSG7TAeH4W5iVIYcqKCQu/FEmdsV4a2zdCU/9WMgbFJiJKHJ1z4QVNdEeKr7WUt5gwOc
uj/7zpm/YmPest0PfHQGL6ubf/R3kSsTh7HYsd/qfL9tmcO2v9kvmn4OH15Huq1e4kZbqEhVlBkp
sEpaVbGnLDGwlL1A6f6I9hQkGeqWxoLVV03nkjdyy5M6lhC9rMWh73U6M/n5VD1gotZblCU3PrJs
boB/Wehj/tuig80o1jC72JuVx/esTDs8SjqUpsyuLitucAQV+VWGWE7fpzKKAE2q+Uh6faPrGiXV
jqjdxjHLzrqVwjyzCNn9q/Ole9hvF2O3FRvYUBmEZ5sL8Rt4pKlFUGRKE6a1BmXVPx6F/I5J9LjH
lKVL2Kpds1ug7zaOCADCgbpC1xbVBbs6IiPdsEIv2oLyOOKVczcsWTMKmcZewdNBB/LmmdtLnCfL
6V/c/Qq3zDZgzuxZZXXFYnv6JWFPAnz7c8nDc8QWK31JtPH8rxVFqtrQnrHO7iZ6bKB+lk8aMSpU
tinrtEg/h30MM5bzOwpOoGNiJoFJBjNGwXCtR2WB8t4aK5xMOsH135DN5FuQcu/Wv7931yUzoazk
mbWHYdFwO4UPfdiXSmB0+IeBFX6rp/wAFo6SLLO6bMQVvXbB5U1fhcltUOBF9/JMLvkNkjrMSy/s
ogFFVPXkUvvhsSyYMwVueP70i0Qn2Z4HuGCTTQBI5BfxS6+zX0KoQ7vbfPy+0FY9sS/mSwT1phbZ
EOu5pZNZojpM8ZE6Tu/o5tdyj0fcSxnV0rmQADbaEjAXuR8Xnec7VwbioP/eTltSLSY69kwrUMGw
TQooo3BMD/iaxgarLHV9NZmcoq1gsesuLjILxf93QJ3c23XCbPRtW7WM8mQxGKRsPm3rYJnf6Ltk
dKgyCxp5G2fXuiFeTsthQWf4CYn188JIYNXQyIqgftQ46edGeOsTuTMTY2Bw39lyJGrskdWkVGmz
CLdxTIwSrB/JQr4WY2fbAx7nEceyLehMSb+bbBtwaHSed9vIWu6Q+NC1qp/2tS1BZ90scmyMi84o
Hsu6ZmTbEgZpPMh5NRGe4l9wVAIbCxDWT5t62qoCZr0slC9l2ZN2Goq1QHGBSmwDW1wgqzMuFTtA
pAIIAD4XwLzlh5LzIQzoJvlbn5r2uQHUusp1A5QGpjL0Jf1A6GsQqe8lyge0zghh8qoaXnkxQMSj
QpnP8rEBdxgPUTx8fDTyoz/Zapsj+e3Pp6qUWpwV2opm2InT17Z2/GxVJgzBbCk4Wzdm9UOQwN/u
q5rIaanmOMvFrTUmpKHFLFnT3t+/jiFkdnVRZJsHhLXnYKWDarZIz01a6nsXyFILBKf2z54m0fNa
PqzYAHPPR1iXjRQHQat83mSD7HYEUQ1UuJlM6SOtbMHmRJGbGNrogU9TgR2K0altSMErnXpJMuRu
ujAnAtJRm45RGxLARgWgvv6Plwd01jVwj4ze9pzmU7KZogBqpNBf8IdZaJskGPWJfd3U1SEKN6jP
5ltSHRSDBfgl4tQ0lAO7Sn61Lh+Vp1trmIMJZsl4hSNy+3KQX3gLl1j4kv+h2GkYluJFIlrukQui
9zDA2QX+tD0e4e/xO2KpRnI1NEfP58js+lfRLYYVmxIAUk/zqN9vhJtUNnFQxGi/gW7qTFprptRp
2ebGUcoKCAo8OOjRv+Q/1A2+d4TbpTRKPQCq/hRzxI88mQwClRziQEhrt9VvkcuEh3NXNo6cVBj+
53dsG0Fn+6Q8Jz4x4ZhejuhJCnmRnCkI8GBjhGXaoPwBKc2QogBDkI1gqFPfq4GfwsLFzU9F3f0S
sHSXG85EUZYPkFzvYyL/8qgBo4YF3SS0L8FUBnJ5WQVI/U6fycyTNRr/LbKzwWasnyNLADARvb9B
ISpLVfJG6nWySQZrmDzWzvDcrfkx908ptV9+mCM99Adn4j9cfG7IFxF6LqLQ1T9BvES6OtPnzLi7
oErTugAN5CGT/w/20E409/dX347YmoEkOVsGRuJYsZxdjG4rezD15t+t9/u6nWf+JMkKd7VYTJCD
B1WtV9PobL3wXzv6xP0a1xrhtzz74WgI6yISRfiZcRccNo8gs4yvqYOc2YZfM4+jcIGchX4yoLMG
6o6cwaRkMmvCOC7OJ7DIGlDaTG8d5E7B+mLhzX9yXuTwV5fbwkAYFrxAd+JYBbGP7aDhqxwWS/oQ
q+LR6+gC6pClRP55EMNUMtXyGmOiQrmMwFnLjGx+MAJl/0iiauS5rjT+EY05N27iPqciRSHMJsfo
IMo7xQW4lJxDWZ003HkWp/CC00r7pMB2oYdxIahsQDyFXBbcXD6m3eZWNYOPG/raQ9wP2yXA3HCT
UBXqozaPq/y6hyMheuT+xKL9wQBVTeBP4XAC7ellXSf5kcD68Mo6bWiLskV4mpFlopK7QTJuspYj
RqrsNiexbi3CeMHhZQgwrzEWTsh1O4ZAaDIZpAozWF8W4e7uE8OV5Yell9ryFA/9SPqSL473bPiq
/03Bj+C1AFYYOcGXXdTmxo/nSJMaqjHOsRnFNHM+I4y82TAVi9mDKHi9FAhvq2gONYXKMsh3QZsc
ut5748t069OgVb5md62jDsyHHErL7nv2BuL1oFOUH8mnfXLItSZ7xSYxCHnTxtKH05OI0jNgscZ6
p6KmCoaRG56ANexVOSrunaxUDq3JsG1xVbpLYEDsc9yojgPMqZdiilSl9iG2SvIGLM5ayW4WjBlO
Au0lfBY4Ci+vP/e9yQ+0YIxXUfCApmdHRc7eadWxK13eT1QqDCjZMclG2FL8mKLhVwes77Im9EO7
BsCw/mRW97af79dfGg/cnwCTWIQIIslZM/LDnRhjDWmvaPqtmmhWnjAhxNjXfT4zP5a/F2svLF+S
sL5Pux37/8wB+dwuE2aNoqYj8CxygBfXhHI0Ly6zlDG7uG8okatpu8qrRXfbgBzP7FvUc08BCeni
m1ydYqVFlCMy3OqTtOXoyFJ3lMkvB9NRkHeA/RqK9NHPPXjQ7qQFr135Wwo7znBKwR4oydKxbdku
j+b09iac7sD3wIJlq5wz6QlH3wX+r8am7UHNtqjTQQoLKUpjzoofim7DsgWISZZHUAKImXessWrN
jAkWypZMxnAgK5kG5K8oaDqNfv6pzkr7n01cVaLzbhyH5wBtHQnIkmRm3ZdFt+WwQxz+V/+TN0hK
TNzZIQQRWFRioFSBi1Ec6Lle//tioLwIGJcNauREmQhgnzPqNMPP5F+K8trHcwl+fNbKSMAlvPpd
xFNZRLHkTITBZs0Js0lkeeiiDvZS3+n/sE/hDUVQ0jtLSFu33Du1rk9udOm+xLQ2NEgBPxPaGWya
389CskUGc7PK/xOOyClINGL0x0dZdMwZ4mp2s+6/2uEolgPdXIcR5LKVqBjm+Kz6fqlSjQEeggsH
U99qohTQStFrRiSmcLFvj+kvlTDDZjOd45t0UKB63YdbXEUvOqRgkNfqlojh5kdA3a/Q8Y8FVCR1
ayZ5CfTYgS0u9DnywfPCbU7oDDVG3zgnUFZUDWPxnjb/iRztDXiOdTpCWI1iR+fbQ4xLc5oDRKBM
zF3n9ZaeWMdGD6+Zy4rX0vANiUhEM/SlnjN/zBWoQAIPBySY8WQ8MHcmwxxbUQ/1JllzNtMLjUs5
zmmLU5CkHt8qbTvOMMYn+zfjxpxly4OP1mtb5ysFceWofMFZFjuo6HefmCataQdsswDhrCtQeBnN
hHu3gwLXG/lCJ99mELXmr/psYNhEmQVvDE54xL92eXiv9Tk2IgYv5RfpzkyKl6Pc7J+HrlI81xY8
vGezggDH/Zm4xxvaoxQfiXmUBUo383aE72R/2C5ZnvqPbLu1N+3uxf+/DpBx+XSW3GT7GrtblOP0
fNOpB3jOMbQTjMyyyzU+5u7XzvrAqQciYiZXNSs+MyCgmdgjJ5xkblmqRhJ6SuuNK+uaeqInI6mT
PjoDl80cT0U1bw/sfClCw85nl4DGo0tbRS0InDQyfnwcFezdN7XbdaAfMW4qC+V8cWdjGF4aMj03
kCtUwDRsmuNhX3bc2neOlpKmxkyE27qASlDkNUarsaGUAxPGdSjyvTseu/LnM5tUhrqMS76sNnjr
MLa9Sn0N6as8rLDFNj00H0YJ+rYOohD2VKElmsCwQrH81l4XBocAPLrl6jRXx4enO/0BrSGyNF5N
V1YP8dB31nXVvf+Lp/O/oDfkzZMUp9sB0Gfst5JdWp8G+dFMQ8OBmPO+AJftSz109Eh0p4NRRMil
1sF89pRV++P1UYCYi1cLBwPlthjHF199etWsdHsBQXjvFbd9a48MgqWRhV8+5gCHVcsDe4+eTte4
uozSUIKJio6KMO4mPr644faqfSHkm8UCDh//oVi/1ywAWE7MLF7kl4eVw5bHF69K1OXIzfOSBxtv
J7GsfPb74NXHtGy062hORD6+OhLgnndmSdRlronHH7BVftAtARW9P9ahHHPW94MkRhgp/iNouE94
xB4octoEel/trETwlf+eRRirLoTeKx/CwZaxtJfXI/Id0GiPjubkfknCnZWpPABCFkfnVYqp7vRp
KOU3zNWXJXj3DuKsPHP6VfxHFsUmeC53CT3BY614vPDQh88jtUp++kWwme9NK71cyIOairHTudaL
+DwGR8CzhCT9mPBKLJOAe9gnsgVZ3OH+jn7LxxAi7topMNYUAJYGCxlHRVf3WFRPpUNWS+dDwWdb
1nR7mqcv7QJwuKRnNvaumdpumMcCoRsZ02icVQNWsXrUz/fTHHA0bUWja/oPUuZPu5bQT2lGRzPj
rG7YWaVIquEvnI4BMAmRT0f5ZHC6nVO4C7o4CUeaEUG2ODYLaAccQKuhLigqWc6Qj8FyoImP2Ply
1YwJhU7BqnoPIq/aYYf9UlaVhqmZSfn3/FduWGeX6vptMQCh/sfcDm4L+UeVAPS8tx+Wmn2mOLPB
UrockuVr93VZKn84HA9Y/EaTJWnYUXjJ4oj83fOfzgHhgo8VNz2PquX+X1HVtx8rbXi9CExfkoCb
RQxkoLxxKLYlIcWxVxB1QV3RevH9aV42QnjnvT+BHysde+/lYpTs07yrcXJx3FNzRNAnVW+1nEcV
qxmVW3G1JdizoEYaQOfA9hU7R0mYlxSunAGFWF81EekrQDuOTivc3DL/yMGVQzBntqHqxbdhFCMk
cs0CjJYAQxi8qiWTcXrQkQHpNF+ayKz9qNdy0WeZPGkD108OZbNAhe2U2geiaL6zkbgF9bO2k1x5
zYmhhE8gRw2Qd6NnFoLGb949e/RH8zsut7XbaO0ivohzAo3KD+WaFF31V/5/QQJU9AzoRjjgJLtV
7RyvTkITaYlkchiU+Yf81I754/Jb+TPabKg+ci2s6n7uI915jQf0cvgsxq8sPWmYE6E74mOKwQ1R
KNj7drUuO/oER+yTKJsLtVkJZmLTorSI6N5MUhBJ15AdH7Q5mHranvKVbScaSFPb0MoaBidEcm45
Rn0REJ8HDoC8VOD2/yjXDZKLV23yVa+oD0VZtpjYCDLDcxol/eVvM3YmbHCHBlXdvLt2LStp7NAT
zpYsJrsRcuiRCJcrzwoTMX+5QFKPegVvcftbSvIYOpRt3qJcEZj2LCUWrOuhepR9061TEnvH+qck
P9VllCHYRwtK0Ub22YLqgoBI/I93+LRkjAq/GbHcQgmN0ilVNus+iRksEnPkpyxhc4NzgY/qnAwo
/8yB21ytkq06nCJYVo1pzA8nxW8DOPcF/sJvbSo+YCFVvNDWGBd6nHVZBmMONkkcJuPa/TRKyJld
1jtOKebEoL51+MMAPQSZ7LrEQ1jq4XAW9EDsBms64/jSFZadiChs3rgqi+uC5wKr4wbf5ItFul4M
k2z6J2jc3zHEuUt6F/66/lYalpYnQO7RCmXfLDBQ2b8bCzdO37SLhye6ZUxGBKqo7uQe1iKqiOoO
EK7vaC2oOMBpMVu6iX4MRhRY35+iEdacyzdGdf8PxjdlYB8hDrF9IZF1UdIyLnelbIeZpGc8wMFm
4U7vFe2IVHlQZyvnYzQFkfenSB5Qzw2S0dysfHp/xUR1X09QQHoYqGyyV7LF9Ne3FAh0r9Pi29e4
HC0izuEuNXw5IEgeLNQgzZOcKaeoWM+8AVenAr1vq+L5dhmFJqd+9orJpBRSHe7BaMI8sRu7sa1v
eiHJGqXZq7UehfvatK7jOsRASDhlS0Px6VZ8ejgPM/TnblTuF1CDBFLMGiQrBGyd3/e0tNDkAkSu
LIFCiqOq4RcqzATHx6OVggvFpEZcKiKFKhqt9wwwiIC/XgbwXANP/oeuyEWwv+j/UZ6YP5VuJ1w5
vCGa6BrcCXXhlaoTZXXzwwY//oyz21ZCbZjkx7Q6j8c8PjRAOjuDVJriGqwdcl7B358xZASL0vhD
wzlsyczL1lrBQf9I9jod1YhtGCtGjDz9abGJBp+PNqWjEbk0m/mn0c260nMAkVAzdC7en/ExDh1V
i4a/ptIMtZheQk3YS0z1hf7Cj01w41FcNwRVZhysdleSIPRbCJdn7t5bQ98X52NGd4vlM2LNBAdk
EZlm6Sd6tCaaOzQ+cdYFBucOSzwFd5BslrmGcLVCo7R3enuTc76LuaIJYzA9LwcVzDOzAevSgVUN
d4vhgn5IgpLusT7CwI8oi9wam7sFqB+Qcn3+YlH8b3BK1sWujUcV+Qr3MgKWiToHCCtuKddwf4h0
QTLaQ06JudFAnvKePn3ujHfK1ePspomX1YXAjI6kXuTwMiNgNS/TWI29PYbqW78A9NXehvcUz7Nu
2IviA2edsOgWDUqE8mmbmn64r739QVW3vqR7tQHAaho/3F1c7swrZ9vaXh28vqG4sp6lPrqkcWeN
AdQxz7js6tNCyNJaCHN9HPP2fL0mLFzlGR1Ky0v+Bp1xMKCroz07Kw7I1UvBmGZHzn7lgjHMohXY
eTQIsY+NzKMX5d6I6b5gGqyC7Om3VD2C4W+i4RDKpYXIv83myjundnHHNKsM7hNaXSPAAr3HM4pO
NjanQrVN/ytNALZMfFv7VBIkR3Z0p0SCvotC8Dk8FYvR3DtCPn1ZDbwjMAIf0dGsiTuABWq3H5qy
AiIxOs8Suf/UGiyhw/NP4fC6UQ5RBOVSP5g+FSde1CvXKzrxmAF6rNvPi8VPwFvhoR3onFBpsrgO
cdeQcA1HqRMfuzfQDCUFkuVkaoKmVLSiY0Ri/WMyzpCZzSLNZd/rVjo0eWicI0qdAz1d2WCSubVv
ntuLU99Mx/Dzk3hS4SptYg/tj5YDsQRJ9hqDw+pJK5gTbJAB2zTT2sG7hrMfOwaFhpUMpwyDGoXb
+2cegaz/pPaavNMsNDzArd6Xi750KZ+xZCHKOtrd2jUT4OQBfC+RC0DJViNuYdmIYNAF+ZvvCaOJ
6lLhKV2xUWtQVbvmoFAsskIILU3ahz4UMi+2wkI1W5UX20fz1lmdUamPKVhAq4vSPzBsXUMaSKES
Z82eAKfBDaPVKiP/OC+hcCoeHcSxOzPaedZC7pxEGzkuxWTmmyYJoF8Nz4n+N2i9bAXaJZJGSShi
Pv6MmIIOmG6x5CO0RiUyUNR1zIZmVMAfNR79ie2WlhfkC/aghwERF4KuVTdWRsG0JfGKdDhrDxKf
11T2mdwsyQgfnmkT4RUtV34rnmOXy9Z0EoT7E3n0gqvkuwIvm7knC0SHujsxd2ROo/LnEgUk9CKu
zeMvlnEzDBkoh/3uokW2XpVCKymi2qC7YJQTmLSoa81dKuZQpyLu6XDWPluEEjHY9oLgxV2ntsWf
z/zy1JKhCVi+AtfowFuD7c6a9i4aR2vMa90MQDyXjsxSEczzKjcLIM4dl26PZU8uJUbkeSYox9JB
pQUVSrsiwzqvEvjERK6tvI5YVCQs1j+KxgvHN0jUO0/b5XxgePHH9nacgMD7F2lzWyk3bXJYJNHw
dgl1osB0HRY6gEuVXHi09Xc5hzQQzEA8OTcnN2lb+H7VbdjCLF9WPwDjShu/StPCx84/MhC7rebc
m5TEHBQ9y8dASC77OsFECu1rquHIUKbgptJTFAjq3ceQ2EYkY8X/BDfm6aVFU7iOQ62FRsXiiHc8
Zu29JKauLDWEypiGHnsvFW7qJiqTX2kegBQpHfN7e9/ImHFiXienCyDf7bUtleZ6Wf0d7mKXabCs
6wgLcixO3/9jOJ1RRlREFjE2/+MBVYrFJGo8+xFoiezGPy9Q9pOyNynOxkO2dJcPvbsWZfjY7WOR
3JtQOYAnUc1q/oBg5W4cHC+u9LxhXzpGr3I1YaSmpjyN9qvmRNyOzmxN3yLkPLJ3tD9UucmXrvoD
f80kD7Dyw7J/diqmQWralY6fdX8G/AXwSSAMzRf8SvYKXx53Lvd7TfXymRhNuCBSqEnPcPmaRl+9
JnZnBd4axqROq1pPqnIMSlWvM3LEdhvy5rdxuMw02PrpZdRh5OpEXw0woQsUAU0Tj5kP2NjOpp99
Oiu3yM+AkJznKan4oqmgePkn5Ga5pxhDGEIOb6Y9JdtHiZTzHJYUms37tJ9liGTLXnosSNFl+Poh
9k6u5BLSqVt9RVDldX0zB/gN8OvsJuAN6XaianUwPnwzgJqkkuPW45yoY0w3lojEm1Yyx4bWGBE4
FkcuytjXqpUtB8WXKovP9rV6qq+wLJoQ04bgWuAFRz4cIZUx/5x9Otps6qyTZXs5ZAZ5am+ORuBg
YgYQ4ETIHqXNWeYJsNdvWCNpsiW0K0WDIdojDDVxC+kzJndnr9uyVZEqKICyzIndP0Z8dHy2lOUj
FYtLbImQALyTC+KPsju+vMFDnaPP388CQiVfgy3QxVBhublVEIqEIsPOHThzm6DOXLTjeB7/HO5x
Q1laAU9wJ7NR8/HlmlcRlWShDFxjfWqZEKhPNNclbniGen+akV/yd/2f6ySOwNEkdEe74lOoXCyi
D17jUAs7gh4eJRWKGt6KB0KB2L63t7FM7y2DKkgb4xECYAHF5cTLMlFz3LBh5IRpTqMtlNAkUXb7
pkGHwP9BvYzoZ+rGVt7tFsp0Uq0Pbp+znc47/Foixo2wTRr+cAXWI7mVGpu/i8N5ue+sXu/RO86Y
OlTH0d1YwsYmSvo7mc6oz0vs7E/0pn+ZDG2tvJkZmYa0wZ/fMdmB8AWgb9sAXzmCDzIfUpA2qO7p
MCjojaRqAC/iAboKfrSxJswTJ0EjY2l3a3NCJppQ/I7jxdKwE+mTTo0gKBhzo5CnLYosP7TH2y2H
BXuuGcIFG6xIlCVihl+o6DSxqK7OZ65Q63ab22SbpkHi1uZa2LjFjfVRVwHxHJk4fKgIhtqVvuZ5
aI2p6dKIO2LixhMUrK5Y0AsV8L7O97ImC3BMYWa1L2w7dfsPkupbVanppG8bd0x8shY0acVX6gpH
1hf1Cx91/EkkBvIggtBOcd4vpa+zOODGcj9fYaMym+RYY8FCJIqwj4PWolxgVbNjLGPuVkELnDTS
Ac6KsnYipZP7qEDf5bNhOq/xPTFuGQ43LQMqPs9VxsWBraEVuxxb0jyoRDgax4PXGkIBrmGbNnfU
0mx2oQ8YewGWgtC9PY0yoxOXuCFZ4AJB1TgJuy8h+CYt78bz+Czr5rc2oLyeQa/0Syu0ieuLWEMG
XjKV6F2EQyo2t+Mt75w8Ti7GWc4o01fGz/i24JF933TQIkw9ZMf2NZtIyITsDg18BUV7XcEnGr90
MqKJ1Amm6afbSx2/p5NJN6tKR22x7BHUDyTtZtI1IoppekBgnU03vwqnrNGlSKYt+oD05ZUqRQkB
FC2X3MNVYgvZmYjN4P7fVODF6SZvqFIaSEi4ukPCmI2mDuRe47mqfER8JtRMRHEjldiXpoaUccuZ
BhNIFZUdeN51L6gLV55WnUIf0RW9NQ1Q3wyDiQqkPZBD3j0ebsfZgRcEDG1TUEUF2cB+46QUH6pj
OgbZwPMcfhcRFBLwt3o5CgLL7OVIzDWit+jprSKHEgQvOLc91VzNphGb/yuWi/pC8NpPprHzIsgd
yEGCY+3DI4HyXBgxVzSZnZQC7TF5eW1xQ2X7fYnTzLw1YmG2oJDbhdYbSysGgIzrC2wynEo1nIus
MHnnR2tV1/TtdB46e6sJF2PEY99S+N+QgcV2vu6oZ5ryj0wQh7YbVv8/cmii6wveUpmJor7fdJPZ
82KbwfGXVxHufXyTzP1MrfogKL3JG0Q767vz9kGWfSENGBt5o+Crf59oZrCKqYNBvVLh27wIu6my
dneQClNng1brMEzsp3Z1s1mK2zmV24V4gcdTHFBUH32RnRu+X18rc/hjb/byaT7pkoyKTGjeZgxg
x7yr9LYlI9THJkzrLk53tpl2YIWfjhIYZ/kIdIN6pasqIpHkydPPEaz3pYejFyWDZmhH5VZUSXbk
4v2nJ9Ip6R+YBHH2vBmZxWLgMfG+no1m2Am/lh11RyRZKzTofxxuRdHmm65l6wqqH4c18YxyNwIv
hIIBITcDBpujsNoQMEoS5+p4jVG/0Ub8i0CcMLYC6VVSw9o8uoF8yAMMwB+yKgL3HVtKRYeOC+AV
INNuVLE0GAHREGv/Y6b17YVYdF+ZryInEi+fYUGQyEEDE9BjHYXEfvrsevJ25GFsUoUCX8rUHGSZ
TsW3gjTfAW8Q0wGOORumT+69hfUHw9aIXnUxkG+Ux4BwXmpVTd+XZoilxwve7/w75V3pUqUvwpRV
+bHMRBIabE8DhRTzpvuL8K6JmKeZ2ZyJRvv8rx6VNI86Dhdud9kJtLkXyIBHLxnmy1ZMvfVXROvU
ZoCpiqOwpxU4CK7cpLEcsj2RCf1a9pMqeLFHG5KC2AvdyoQvQ/dSnu/WhYBK3NmzdfdqxVBm4MA/
vVjxGWh6/2+/N3eh2L3yHEIoxRcYzAk3VyL+vcVl2GqIpAAN5m3nB+C6s+KZPxIXn0kaYvy2Ka1r
kt9JSb5QRGCVJfacEYNcZVnlD9lKGUKEsXayo3lGWlN9LTE5GxfYKQIUWfFVOKP4/hv6zUWdq3+s
qvZBA5pcy6xdGbjYXKKdTufMB6HfE78ORdA60F/4RLhIdvZbHPcGqNwd5bGlKQVOXbDRofZmBLfW
nMoe8wd8O12opsy79NQ3CuaTa0ApP1+DNEkTe5im1GIxVQ+s0dj4aT10xz5vnQLL2XtK37te0hhf
A+v1L3UMvda0mfeuHDv/ZCkKqjJQsa6IKGzJqR3mlu7h6If4/PPYYgFq4QqOVbsMgnDLI9gBFo18
t00Wvi1M5j1MrpwWBZjQip6mBucwZwRH+57UkBy6f/llFIPhHYEvQPAjkAc7QPzj6Z9Ff25MAH4U
ptv4RwA5TmSYEDiR1MHnUmT3YAGu0yOzTxPUjI/E45fVnkO5ZvIBi8n6SVRj0H0MBeFUNRxg7kVk
7WbxthppmkIbo0xgucvvSk1jUCppycfLSWq43Zay5xiUlY9u8I9eWyeZFnYmFCcphcNpdatqikeq
uzzggrJVajRRtSHzbbDyNfaSfI/rTulVr2f++VuTVIFOGJ4cdCQi7QVJvEmJOFh9alRIbEeNzCyM
9IFUSyBmllYy92kgSx7YCVp06qeNQRUWDqPADM0e8dK1PExAK3b6b2EHREXtQco96+Jmx3/KEts4
f7hInorkjVWkAHbsXRdDvvzyAINGvpHfvENDXMrulZwughni6az4XtWL1KtaJp1Ac87LhLJOy8/W
+rgrbUgysXTuz/gQ6tgxBj4qVM6uOVIaPnKfPDcspTq+K8RJLvKmgciaWTlKTvXuc4NgRCbSZEg8
0OKvPsjju6Q2PchSDWPYa9hcoImSqcTFG57bDD8e17+TEELiqM/+Mr+amMwfV0oYSe9A10esdLEz
Vig/gUxem+2WWWA5GnD1Dl4rjs5e1FbP0NUnjVZUCBVO0DvmetKw8/GStK/f2sKrafpfAmjFpn0E
D/k3gvzD2i2r30KrYfuecbOqJedopuLmPQSeGwIe+F99oM2zRp1AlzvOZAqgAm5Eo2FnSw3oW+UM
MxJUQmCe4qFH0QyqQ3mhz0i6FUOZX8e7OJuSL91PxLrNBk9ajXIeXAUFS/1a/d9R3GXVRLwXSXC5
BxUnpnGjtopevm++BeLgKXMGPBMDohsBrYG5LkRYduY27nBmo5YzQV4loZD40q91J8Wuzeis8A4o
D4lUQoZb4RmY5OGfvUSp7dOmDlu3rkl9XNhY71+vd1zVDfQWc9wp715rm4/vqOs4XiQGHKC3tV1Z
JQCzv2CmbiFW38fjGtCTwt2OqYGQLHDMJw1pHbptycjHVY3VuHJTIcY0NiP6esFqFXLmglXCnBnr
pTIoG3eG1yx5L3g1aDL1xlWOEtd7hpoDXKEwpBbZgyHuO5pKlzpGQ6a1jY6PU9ZRbXAhj6PFoIY+
FZRa++NXpN7Brbtr8C/aqM+oj7j3KhYd2iDf/g8h/IrueflxD+KRbeWJAVygt7RCRMuUzJ3hWOjQ
HPXklYPLHmrvMcKc353DzHsd/OD9r7/KmSkjD8AD9CKL0KMRI6/8tAslwqAx4IJ2PDGzj0vaPAeL
ueE+VcheDrIRV5QlN09R+YOFREdTX6ak+PgRYKMF1lCEmtm1SkJ2nWVmaRHRRuj173bm23OMygJ9
1NcwrsjE5amgn5aj61YJlKxGncz/cwC0sXknLQtlMOZTFZhEuuSvRxlGqY5v8ekv56e1ABb7V8pw
GHW/1jBHDK4uY0o1snJtarF1/Q2+rzSnm4nTuyqRrk32kwDJQjd61GLvbEm1DTtDFLbFwgtflOlZ
iqLyfnk4+6RS+KU2DPilhopYC2amAcuBO1qakcFgxat8Bm01es36bgGyepxSWKpODakFSLzkXBQ4
4mTZOxqbbNh1D+2ukIrumwU1EH7f9kSYIbWaJYZ2AYF4MiT/wKbW9LCAw3fh+or1gLWukR24UwTF
IhqcFe9iXhE5e5a34FrX8Nlcur8GvRcZZPrZ5yTWUDHpObVvoGB9qIajxjIPAiMTfbnFrFdCEgZu
nq7BP6cO6vVc15e3exlEmDfhmkmZv/KQLbL8P1R0fsjZREy0133WxKflE4zKiykjPJAGhvuEmNNY
WEC2FAz+Y0+4Xj41dah55lHw0EXpT8XvpCtxmlb/TAtd4go0SNKRBVfUayjsjLMaXZae3eeOrwn3
dc0nUWaLzlSb86T5nTUwHyWZSHVpEMjOyEYMNDYvkWQHgzjZVl/ynjtrkg3q5Au5sEOoQ29i4ON1
Q5Za+ocNoekjstbX1aaFNZ0FqpLf1DH+nlfZfWtSuMPxHWhMcDmofOGAm1r2l3CtZR34IYpbkdRJ
LlKA6TczVoGQIAfSdGthEXHfeTbW2JXtNtkaB/tnUE8uJ4c0Fdbm2qYEWQM3Lo87pcoN4TrpPEpE
I0EUg1QUchOc2IZOcmhCqYymQ0nyCGlT7XCnKU0lwMyhV1WFUZS4x1FOfu5fT9XC7qmpUrXJcRwg
gJae+N7SQW3x1jg0ZqWf1K9Ib4wHaH4DbceyPCHu41eiU1Jfp3+XOY18oZfktjUXhhDQP0hoOOjh
7jeRUTpA9a2rl6CG/TpngV2vKhx+FKE9NOWNsILaWfXO7ZMUi9b1rNrFGO8z07oguRHp++iiZQsX
HI/TGCWQUUP1ondQepTW4xNzdb9nVWyfcNONVBAsRKSUuXplT7qz0Y20zBpYUlkgMeTC9vYhMq9u
xh8KH9P/sj3PcNfG/Li6xFTlNvgD+sUXInylT9WNTwPzsER8S44k8d2vvX6qdwmTs120YxiZQChi
CGwkHkOeFeMG1AMP31I0DMvkgU3o7Ahr2r+LmV31KSZ1Cofhfe9pPrVyrFQi2cxL3aHeHiQ/gZlq
SVlvyPKOXjnGFaiEkQ/Z1/Hyc7jYwjZxLBR88LEWmyGcIqa5DL4hsz0DcJVBeEBGP827S0P0W1Ud
HEe3+u6XL5u+qBRfrQGxIWz3vUSHuQjbBsIAfCY5hGR0bTVUWA36nA3MeCS53V5V+SHWO03E68rT
zPpf5o/p0NMqf76l7TUK4tQaMTV37OU68Q/lLAd1JNOq446IcQ+iUrclotEj4EnZztMWcRdyfI/c
dTp8qGA+Cs3B+pTZKg/sQ9+E4krp0Z7w3cj4ziTqVIn3aBA45h0Y04Y8ylYbee2oijLciQpaxL8O
Mapwo2FDUPv4EefKl+8gACv263S/cH2M+JKM3GOv6XnxOFwPZ/iZexVv15zLbX2uHclAa5T/d/33
iFdlyMBk2qK4uN3QUGL69ShOKG8qtBS9K9QwDH7JTqnCy8wY1X+jxbf20a1GLnk8rN5X958BrZRG
fKTKKw6crnQ8zDFf6dpMGFypGcVEj22x3I7votu/vr/t47LwIlqYGEwmk46lV6/Am3El+rW/IBED
q3ger0sdufwQAcQugzbLBW7Y6eir5L6nTDZd1PzlE5cYxaVG85Cqk1zpy7ncXUW+yRY7gbQr6ulD
4JEHRKKMu7/4nkR9r6u9yqQENp8BaxMGQTYip+puF7VN9Bo84a9nGA316OqF0ik21icJHcrX6eEM
XsU1pY9pMYZxtJn0eAdkXZM4OBzWBInczyVu59+o/7iOBU8u3SXHxsnf1/esJN3tpynW44Iyed20
kXJw0NwhEnKcJQLQbkRowGdH2uH716g7wCR+plwr/nLIBXSnDqpuD+arc5TdNqeTGHfewPjP1uFZ
5tLdU9N1eOHTDz6owVj49VoIdYLWajeTlLeclcAhUZT3t8GsVmY7mTG5WpEjF9JDS2/H7AWkpiXO
wZfS1vwm8unPXWMOFrQIhBJbHS5Wkn5pTk92flI/9fVtYSuLEfp81FVp6YmvWislOvK/Xg9Uh6r4
N/v9ScgkFTHmqiyRbKmQH6JlcGIbF64QzCUSVOEs4xi87GJkEBbqstmsODQSSktJCfRwc2eFEUAk
xY5J/TVTRIBhmAoWOB283mT3HOMstS+QxYrNQTlt+tkwU/3vHh7c5wtqAAE5et4i94WnQf//gvNf
OR7jqEocCS2emGg2pO4Dwbh3Du9pBHbu4cxMUq9QAFn4pEYhCnhN6XVM9spqdcOy3u81mEjbK9cr
hADKJYktSL+AkikOg9Y9m+CkhFhQxdu4raUdXiN+9N5ygPlPB22SVOH/3BDQCVbV3R2tQJqbUeW0
5x1ti/Hs6lT7OesP1dxsg/5oTHWY4gGE84RkMJqwZq6uEURrjVhUuILhiYKjYJWeEDsCBh7zc+r6
ungiOoubsLPwSUMlg4bPKhtClwfV1SzNvBYs7LT4jFV6/ev60+NOqFJCmbJ5yJRRffEBvtmOTK82
bZwbJVj7fMtoEQbdydN5FBsdvNkBKi1A3tC+PNXxOb6vyrv0Y33i5vzqbS3XK5Ly9iLPpjOGpSYn
u+ln2/ySJlfo0QAdQlJvznBMmeXh90hWpORBh128I2W7QB5GUd2m1PvvEO0hSFQsNUge2BgL/d8G
qaiIOH6nNrKYwRhL2J+8lzM1VlvQWAGgnauVq5V9XEsGDHjn95/Ig6nQEuJoxq2bFxOFLWOQKIaq
kr1afesMCJyGdUpvBiIGrELX/dpvN44xilkr7V3f/tFFO4zwNwxsMWH9k6xWynkyPG9TTAr3TUrj
A7ehozWLBSYfEoEevyCqOW7cKXce+KFea5dD7deDGy261VdDcnOB1bWAHlUqvDzQvL0f9Lap/2g6
7bp2vvev1iK4VXGy6omDf84LZOEY9yafqkDc9o2j3I0bAy+yXsZ7ydmwyOYoeIQAKLma22m26Oy0
D2cGJ9q1LG/2Wpokmkoe4wC3EwLQuACextfqRvtEZXteX19+vO5Kfu7qdJSsrzRmOuEgV2YcqQV0
vnhFiO4hv/Jgh84mv/OKhmzVxajEX5YWMX6MGNhkDkC8vb0LphI9tDDkeDC95Ntrj3Td5eblnV8c
Pw5B4hppDFeYmQARXxyE2rM6sId148TxeMCz6ziFHyPLriaD4HtVS9tWw8d6Al9huO1ssxNogZrT
+ZfLWG4Pdp5dyEaqvFFLT92EvZHGTTb81vsvI+JKEbYrXj5xcaFChtVG/waMeP/gAmcihug+Yniu
pLxG/rhjg5V/HaBeqW/6Z8ZAzj9KXTLS4Pdbg/4OSWz4jB3I8U3WIQ7XBAJ2AXyzsO1p7W6n7vDX
qeJSq2Hz0Vef1nRiyqTPHwlTuDVqd9YWFaaxoza2qwFdlv+XAPojpfcJ8Gy24a42gn1YDSGbSrm7
3/vPf1ZlafswDhHQgFvNVuydd3YksEy9gsi/ZcjmWBlPBOvqi/lmLpoo7SsYvCkAsp1nnqdBzqBi
96UWxhdu6B4bvJmd0YCGD0CfeYi/WGtlZakCfLEsc1zniBOK12rZuI90J+p9hjwpejaubDJV9/pQ
5HtLGR58/e7Snvs/xE+JgV9lpc8B+Q2QNkqoKQesbeFwja8YzthkcpuiLFlqQ5MJViE4dv5IhFdY
qt39jJFTCMVGnLbFIOBbH8KO7c+WG/LZoWb0EvSqABfHi8Am/5yrulC85U5UNy20IiGR77t5+oCu
zqGZshBj77mS8OPDVhyQ2TKp56a9fB0JmvKxKTXD0i4tALVN6eFiHz/+RiDNLMB8BbE6Zs3kCr90
upYDNy1Sezy08+p6DJbFPyNgKuos7DUlcOGtRLAtkEREXnvHWv+/DcLVE9d6Wcfvx2rwEqsgQN3N
gsQE+a4yJrG6B5lHj6Hh1tv4mq6fKylo96y8fnWGATaUGizybHHApminhk1KSWGcymakRF0x0XGo
bGuAAsryKU8LuY3ldlpmyNDyUIFLOb6LyqDUSbzGD1gNMSZReO2J5NBFYMiKu3LT1cbDpy9UCexF
Jiz1OhQ4Qws2ZLcZLppeCXkZSHPE+EbB9o7z91gpr5Xf8znWawXL4jAv8a2fS5rpvR/P9tVVsn3q
xLaJmEBJnrrTPXBl4iaAc5gpRV80FatnuRxsi7nNJmh5/FADHGzlsTZDEa/elcO2XS1+9/1fQDUS
+Y3nBnkNZPycpR9tXJ4cowoSdoQE6FnsO5R+qaADPoJw5uXjk2oFo1hYZ6SCVFwCIrdMpXjE3W84
mmaMYtgznOoANcmRvS5imf+jVU8gMjPsJ3c4NX8qPZcqcTo66shTR5WI4OLPyaSO+hsrpqOt44XB
8ZcZQggnyw1fLDst5qwfpy3dZmx/EzMLi/vJeTbrQkBMabEJy203Uj7JZiW+hK3hyyqccRuyhWjL
20SjmiLf3BUS8klrtwhBJhxUySIFV4lFUXVg18EJC18hQV0WAHvV611eqx4z6tCbzDWorWzc5P7N
+uHbwnM/etg3643o1gjZSKapBZmzX1JUl3Xt3lTMD4cFC6FDZiTIno8EXBwQp2DPlKZUylbL9/cw
vfHJUxPNiLfpGCo+ctGqxyxyR5NsYr+y2kgtTAdTlbfrvxHRbh5IyUkIcGP0SYmt2TrBZ5vkvF+K
nXGv60izKWtRXsfJwNz22JpugfDageNvWVYZ/0KZF9BjjaV285Uz4Lkj2hQWlGmGLklKJc6qnyeJ
xJfah6Q9azL27Oxl0/TAgAn3P+hST6ArbNP95EtsP4kD23RdtBa5+TWyYsNj9IgMp4QO4WalQ723
kotDLYV5xYrOabZs+H1ezS8sZVBKt6qhSRGIgB7KDJZtNcxj4muNwn9YdaJkwaEZm4mztOr7Zv+d
sY2Pozf73aY4bnhN62rSdpnIQDamAqkjUV5ipXGPhfT111UUOuimYnHkmmIlVuwCsbragHHhez3J
JtFb93WS0gD2U3z4XNhcvWj9nKRE+icDVqxKrnn4At9qmH1R0G5Q6wiY9WBDy+23fQu7e09eV+IB
40PXKGqxKHwDI/y6lhgYednzuVQ3NoLfk5QISS3P+ExWQDGGvpdCPZ97Q11/9U7TivEt8N7918Ih
7NdbR9bQybsX9RIp0LWyanPbfJAqWRKIahu7Z045XC49oXpDKb6i+kGlAa+jmuI5MAMTjsqvgAOX
E7ZNl0Oil+VM81B8221HOii2xU1yQHsMfrWfhB/ckTvxwjlyyfX//TRdbcPqFK6CwoSmjInF+Mxe
0RpiIpuacn+tc1twYFaSXlGywxRqweevRtFDPhS4J+2dHgTN/lmppetwLqYDqAIySIudOA9a4LlD
00mqAnVuVPBP/5wb/jVzfrLvXN9HS27MkrgmdYBC5l3tncPVqviZ8wBNKA26UCEZL3B7QPf/Y8vH
yO/imJWzOYv0Apek1xzFNEtywQDW0gXugMx8GHb0isOgnUsAsta01fo7AOLlH9SGSQS83Q3rasAV
yJnInC/3+Leaqi7AVsk7J/J7czXEINWRRSD/F2A1n6yGcnvYYzBPzMPeugBqMq7kQ/qP3sxIlMUu
MpTv2n+3Yby/7igYrCo4HuEO8HB3Njyei+/964wCfbsDq+59X7/g+Ob6mVb/eViijsJsM/C6oKHn
U9+85sdkodWFRI5mLMD1NJDVms6ebXMILRsRg/uC50erUD79VIWii6ytBvf4Rz3pVbLmMuvb7OtU
pllL/RaslQvGqlyRCIMTbIreLXaazPr6UZN3xJnGBG6lI12MpZCTeS8oFzN1bP1Nhstx0w3zbzcr
IcwhoTeelDt5ryiX5b0/Nh41ckXi5UHxz5p3X+yFSk2cO5ATIc2rR97YFeezP502B8WC4X0SLswd
cP2d4xm1cTv4Q/8F7noQ31dWhthA/0bnvXYwjDKWh1Y18+6aKpuYsp+EpuL+ebctOE6Q3xpXKUeW
Mb8tbEkZuqfDs4Tc+qsUDVBbtsGKa86doLBzIy1lnJ54gxVkdTWL2H9R+u71e1OEPUyYioPDpRRR
1dAotSA7G6G9VaR2MAH4/z+CI8CITikks4WIbf+sSQIlV8sR/4dT1ZPFWU6VZEXsUyC4Z0w4+FzN
lrTtreVM1iEBcsjbObLV0oTTRQMzPw3t+BMsoBCzlOS1HchaY0DmZyTaXZCULO5gkV4eQHQ8Ksad
MHbGPWJL3tg1LjGlXWf3OF1+0jriUynUJZz2wDEKRxpw/H4rISDjdFQCUWCMrQ+/kU+EdGuByC+T
KcS3wqEcx+v6cMDRTdoUJaNAq9WOwdXpe45fgotzcwWl1NQNCX3P2pNNOYgkIELO9D+u/17KsCeQ
IMZqKVXzU2V9xC3YXPG6o22AVNdyo6wCi4+gmI84ER5K1OhA7Eg+olDQOaqAAqhFTcr+4rU3YgdT
95p20dwFyztqpjU7JOql4Oi4c52IyTXm0pgIVfMR/aVdXgv5sNJX0mz4zLeAHhucmiLvNJkaLdLB
bXjK+QCtLG2AEoNDidTjnE9E0ZYBQVrRr0X07mu+psMOT9cuhzvW5O5HVQNexDqH5+Ml6ovmHfOr
f0yolxjM9i6x6DJTngMTXXrkgxSq/HTCDxbS1Z1ImLpfPOvrpSmY8/eG323JPUIhlxv5OAd3oXvI
8dtU15oJSNm0aJFLMp/aXAKvwWibREv2CkooFB5XI+RWopBW17XVGifNpzSMMylyWpOQAoeE/vSK
LNw2E7VXxpa7JNjI912IItY742KEx5+DIUNQ/WVXUvtM3OTlDrS8kL1ftBVl4BKG2yEpYFyAhspj
gT0ONjg8117RcBDmjzP4qJRM+tZmacvXq4fxZV5pJnxnRanP/cLxRPvMjGqfj4cCvpoltDg9oC4s
zKxLW065Iz0FkKraOfs5YDQhAhKKDOjTmogW5WL6FUf6D83H5DqfPTsAv9UrQbt0wYF8r7r34IET
j/UXXqHnUr+0aWlap5MuXoct5TB9C8coP01s8pVXmekvP/rc3yA+tNdOhTevyN6uVJ10YrYbKHYl
KiHmwc+sWrFPz2mjMtuKOirGHu0lfEZovqn+TMkO2YEk1rgp415UMQVZsNJ6lD5f9LKZI3KdIQUS
lZIuZlMmsk+hzMWxz7AACI7HkrrbZuDfOXxWPyhGeiDEwCXcOPdYc8bnlv4RJCrJTjfZYD20UNC4
U68nu3z2N29HIyevxrQBnMrSR1gJd3gcFG8iYId0rEn7/Is8dNFcuuxQnc4ntKer0TzH4x84lb53
RdvWBG/ZpQCt7RzpFh14m5rqc647yPPZml9jEvXfS9VvLnt+SYUSy1E7Ih6zCm4Bsb1NQ/ISwlf4
CUJTxQrJnm5p63zBNqN9KJ5Y20A8vizIelHuB4TecNeuYSVUSGo+fm3PpR3REEJx1lwkcCgAvyYr
20N3YtmEfwEUo9/XeOzpZMUvTdk2dN5ZYoWxeG8OZpbk2ctUCIae5prG0GeWKDsWqweWFj4nOAUL
RNV4AKr/lHEw/BazlVoCNMRCjppiCbDrKPxHitlvNLufvycZFsVWMB7jJiBo7+I36wLvH0H7AQmN
CK4VcDBAmIU8AFJkNxMrPhO2Ou/XBupYPc0bV/DFBMH6FdPpnbFTNxBUj5zJr6+eC5fFmc8mVgiY
/Izqxd58A2nsATC/jyf9WWeOjpTCC0b6RAEtLEg888gvh8Lmk8T15dlewCJRDYgyyTqDbcgR41x+
p1oxk1uVhYa7mR1Db1HAAaHZQh1yquwL7iKf02DdNTIfRBEXKLM5AFsjMdMGnwk8jgz2F9/hYHO6
KKhCvXPMDPcm+AQKeJ1JNwrrIsArga4PWqUYAcNkmc4/M/iUK40OMxqX/O/XqfR38FBY00FdE7+j
5XKPFKjCZUeK5aiwql+7bKKLs4AXRbWjuMLNKRhbMa6Xu0W539zAc+AQmprDSm5LMW7v7dTdfFUH
YsQAexWPE+LF3e15Of7PPOW1jKRJp2wUGi7nWHaJgicvoJG4lVB4LqbFDCrQ2ofCd5PGWRdBw2Gr
DgmGUwq0rHn1l3Fwx3RnLe/4a4+7qg8EvCcpw2NFQDqyQA4NrvkN8GjfcqcCX30fWghVKu95+OX7
fBqccMuO1EnTfo/6KUizK63u4fvki4Fh3V4WnGKQduCsLFNHdUTx5/ZS5emZZT2mRCMScg5BitzL
3V3bpZJxaxVziUwSNbQCRCxp6v3OQ9lDTygK8k0ylYlEqXE077N+dO7R4vtbc1Swfgdyrtmxlk5K
0r45JEgzSU4CXSxnSJb45KwEa4J9UuDShLmnmrdSMWfiC8lc1Pk8zBXDvyWuxz1FBfbjhKT7J15N
ihMaoDtYzE8meiQaBtKI+CIJUyNGZl+CtdAVfbrXkLClEugG0PZdNwsh22qcCkgcsmAYNIwer6xg
DgmaUBrpFapWBnbxW5hk6O3lLOO4xW1IvV2APEJWdFt9xAe2wSSvSbW2y4UxXLo7t50H+YYxWUNK
kIas4rpRE6yrAIjJuOzCzwBCn6AVK67nYJt5a8FtReYTUYltsVkBpG/U5n+GLTOcRYQAeb0GRPYE
ZMSCWi5PAx+4ogm2sOMJoG9bbzfe8Cd1JbVlvTAzk3ra9c8MNyzV5DO2oOa9ahYB8ulMydVOe0ex
aJsAkeaYyu0qj+gdMXlaEYJmC+5JrfNf71NL8qBXCL2ZDq9h3CnaMmg+FxG10zR6MVs7lewgm21l
kXK6+WBYcTC0CYQDXSMwGdqUD+sGJDK7lHH+4jvc2RKhxHHjhZ2MsBBQq9hjP8EdvjGnqbFSoZVM
OKjgmAOvOdBhWEYaHVaIdC3j/VSVtxDxIcxT+QDfyHb2m+qmQnsOmRf1dznADVtD/LbXxHbgKWQg
vVVRHFKqq+iCHuQK0DRwE2rVd3ux9ug2PtJlCwc6jDJQO2HGqmT82WUWTFHeoENwh/UX2EyLH5aE
CqjUNufg2WCVTrb/+4gNsH0uFO7udpSFOc37ffuNq9OQ3GdgR2AtHachzupY1DN4yDWHcqG9jUrL
FUOxpxZXhprmN9QqRa60ct6HoRJ3GQXz9Ue8VnUD6pLiPb6WtEdoTeJinC+gU7v3xtKfthafdjTz
dnMyWyCnJlPnv3LfgZzcxIC9NRYHPXzN2OqKu7Y7OsH3PF0pQIs10uQgGzSnjn6gqisVD0qlRC+m
wEWl6svgmTGVtRN2mAeVxyQMIJmMUpqBdJ1DdTiDP5ez63AXxstmHb4NPL7ll7kPTeZDnRwai6XV
xQJueTFOAV3LdNqFZXB+HcWV9u3FmvfSYvb4UrFPc/ZUSOsppcOmDESyUV2Lixq95lOTxfzH8RDx
2Z33Evn1TOa6UhLAwKdMWhj4UbPH8FjaXJJw5MwPlinep0W0/Wi9TKgFil6UfycHZ9hYa5g817sc
Ek4Km1NcnX6v5l0Ow6Gv6xbYw5E5yHhVR7x+ot5Vkk3j9L2QmYgnma24eXvXaDalz55Tu2bUSwc/
8Ziu8zqEXghoDP7bBTef78sUP65+3P0Skw9HVYWMfQTmYf+MBhFXXwv8k+gbYcR6NAw9FICajOhm
JNiLUOXfVCantmjbscfbREgaE/Tld8baTo/ykQlZyD0/P1FEyHOcNemSaTPZqqZMspHFvXDQNPmW
WTzQdcDQvgns+sA1BRb5Q33zd1J/oy8E7yy9JfG8SybbUgI2ADKAJdVioZoHbKLNGO7ZAQZ29bYG
aGwYN3wEK7Pq/z509nwnXEpUW5HSwxwB6j9cJr8PJWCq3WFlE0IMnYUWFXrvyhIg8qD46T0E2uPd
cG5mpMGTjl6wyeoqYjfNh+0F+gPz6hI75ZxHZIXC3LbVdfSp/0M978+xWoIIDs1owGNyJZJzliQm
QNV3nPgazVswZLs6VF7zIOIQFs16N6Bs6wPEQFoLPdiM4ahB/AB3lWCwiuVsTrnhHV7eckhSRFQ/
GUmWuMVd9cXX3rC8NqmcIzb3lgRKr3cy1pWoVTo1DTfumanH8Cl+wNKWN3hE3qO3pd9Fk3ibqYx1
ChVRHM1z3OFDDK+UC57bjYtuKEbrI5LTfp1ewBe/A5Pp+GOHsww4ynR608w10as42OKHvwXuwScK
7O95QP20xkvvDbxwnJxa8yhrEy71gOxU48n0tOOuZdXc7j0ZLyXSEXR+saUVJrVbnRaIemFpZPfj
LLgQrGAlKRNFLMy2uazbtodx7QftzcDwdv+rcHC+dpadwIk5J03R8iPt4cvBWgiVcaldVxbEJhfa
Wi6ivqaVYwwmc8Gw+wARMuR+PnIv/0LtAlbljdm0x3QQvkFFM9Hiuynqjp9ddPiy2OSCK0ojilxG
JdDLjr3rqrFGSn4dtr0Z1+vZ3a4snKfxAtYqzSIJ4sia/O1kkNtJNr2R+AuN5r8/7eeCyADUqfWE
7+gYM/ftbO4xlTLi8P1bKgkbJ1TBGszoupCm7Bc+0E58f7Os5oaQzmN1Y6k/ArCE9hrtH6I7yHk9
uW+vXlNTTb6iPWfvb4yXEasM0LTGtSkgDySgXltarl7OKlqFzMx34/CPK9EzwQlEnySVdEV4Oyap
0vJRcaBGq+zSW3I09fa5FPepCwgnwhxmPuYBOcHySKnfx5xjqKWBnejba+MRqVx/UysW8LGlxl+h
TtxaZhdUIszOiP1foMoJlq6JsKtf+Ulgwgjdec2Dv1xPtwmlRCf/hD55cdyzobMjmfXzhScPrBye
D6619MYW4YZH/Lf4nAR+JVINgKQK14zuigk+yukCkPUHjvoo6mXHLs3O2SWhrxJILNhd47gHfCKd
usxhSxow4+VQ8VTJDLfEANgxZQ7qU6BsxqZXldBFW42Vcws5EqERQo+y0cSUzTCRJ4kFP9mC8xLu
uC4IK50OHIP4JI6q3r4Rq73pcgZKXvai/QNaiz7HfNg/EquMxIB1jJVCbkBmu/FzaK9QRNZY/nRN
BbWoLPe5YTGBScHiy75tSLeEl6WevPMwNka2soEwO2nmRfSAcLuenCELzXyla0fZlxdQ32hcUOOL
vUXbyv/C7TUeVzNQ6iBfJHUf7wzJXHqXAJj8g2wW0lBcxZXiscDBUKky1OQ5K5cESAIUXJGfCFsX
MzNH0Pij+hG1yiyj0mxxOEfBFomFK3F6ZxN9OUoPOfYDxt+G04+jNam5bkMXDlQ/Y3nHj4XM7rLQ
EZ+udH2qhx/TzJIiAPffDCOHyjgot/fJiJKcHfTkGggnmMk6NVBxLjF+XqOCYoumHizCrUldRwUZ
P+uCNayg11y9MbMNn9bVjdpHkcfJkfevdnhS79Goa6UEAbWJya04pjnWvrggGRYgKpLL22oGw4SR
vkBiyo1+vHhWa60LYr0qMyt5NF56fuF6LiWBjY8UkROx3uGPOxrnUnf+qH2tu7HXFyJm6ZEcKlP4
U7qT48fj5JGL9UdxVojgHnsDZSDTGR3eWTZnF16HdOw4dvrLnf/joVbu59vV83urCPDhRzIGlzTh
oALr22fs5N4uHlUr/H8EiaY21N0ot8kRBF/RW2dqSOaHRG8HHh2T848WQRBDmhSYwJ5mNEzTYPEL
Jy8MAMo2L3RWoh+RKGTY4Ir6Ra7MA4EedkYd3Ltg7H5sx7ewiO8si0DulM/x0yKj7/4nlsyKhuIf
v30GEWp2Bdb3lZkY75PPiUgiAr4WrM6Ww0yXS6iClTrTLQmxtCIv+WV10iuD8vDtGA2WC+2YoTEq
N8xgBQlT933xV03SDGbBZMRJTd8YdQMWYipDj+1gTeQGsgUSlQ7zrMxCtzZ9SAdyL1CJ7TCQXwX3
QzMSbahKFm6LiXBakAY6d7gGi68fPJPHFJVFiZrzi58kU7j7Q9MaUKQ/S369aOtvs51w0/EWALmj
0Yh6Jcs14NO1MBDSyQrFO8H0TyWdSx+Ccc02l/sgukZ1HomKEe82gzoUhfbkcR7crsRWOYNwAR6b
91EuJZBlsmF+3J7jvWyFEsEbcvfAaKEkGskEHyvp6Mpz1xgfHtHDYKVemnAZD4mbGtqpASpFVyBS
fAPUooIWawjQb8pEhSliMltWzHmLJQ4Q8CjH+MfZWTGFsYyQQg8VwN+0gZyL3+xnR+CRMD48uXun
OcNmeoq8FUo1QHeFNDifb3mAVKyQLFagcBHFKZQKYPztTfDT9cQKNhqvSkTuA1fWvZGR/f5IQziH
LJzODGWJ2pj9R6YenzAVzmgDqIZT6vD7+/vXumTv5n8RoemJWfRzvku50rREu0RqE+OHplg2Vn7q
6UdpUSbM+bbQHu6onLrM/AooAtT6hmYIwCxwshM7Ztqf2AxBkWNMRNzyp89PTg4xb86kv7ZEzvRZ
6bO8yXcBg0GKuuTI80RdmLqrdTq3l331CevWjGiwUQhfAIwDRTJOPXiOEBKP0Z7mtt8fS9HfhYPa
f9PPYRen9cGYGzGrArP4GpagwGnV4PDkY4pkYJ0O57Poz/ZbgwTBVZP5BCTJJ2gxGKbuG871b/mg
8SWQLxXHKHzb3lTBMaC/vWjBf8V0JlWnA8LtAcq1+U6AIypaJYjb/LbXtWxWK6K3o0GvwpJv0Dm0
ZXh2CtMQKcKAub8oBAz/i1ugDpsMlre/zv2XTH+TYLr7IhFxg98eOi+HbKUlYDuhVjYNKb4/EagL
HR59ZBwi7jZxAQ4iiWNWdP1fMpXUhho+bN8GXnh0lUpMEonVUt6W4fXkgA1LWAx0DKfmv/CU2XVc
R8OtBn0Yh89uz0rTitraV4xk31A9AQpFLnfxGV4fa+u17nq6OPTH9Zc41BUpMX7BLdpLogX2/QmB
hcFd/PXQekkE+8PdoiQtMc37rtEZv0pIA0hQmRRdfGGFNPFaoY5qP4TrcA/JVrKmXDlPXCsUyE7u
0PWTzBOPa0i1nQCFRh3JlOPMtU31jPQdSXOS3sRjONKWJ+npa3PWe+1O/+ExVYWeor21l9tBDuIU
5g1difR2bud1xxQodh3VnkW8hcGT/LVqofsOvqFQObvLxDIO+PVsofnExMSXTjni/JBudoImZ3BD
h++KrVOrbWFQe7cI/GyOSv0nAVLavyOi9jcyNac1+jcXOExlSu8yU4KATT5NbXcFgNHW3yLTajyQ
Nql4YHbx1gIt2bs51RXfeUX+d4MIsSjLXQTPGFToGD6gN3N2wvojSAtJhbGqjPxyWOAHH+tlaICq
G5JU06XTRs1B/eHu12LmylV8VIL646ETRoHuBMfqsj3whNGuR4+27VbGTPNkwBbbgwIzr3ZRj+Sf
diPd/BvdzkGd3hLc+8nHm3HzPMReMw80ppRwBJyGPai6ZRzr2gdnb6auo+pplvw6/3pEKt6Syj75
QP/Rgva3mPeZRe13ct592guR73oDyZi6E9NUS9xZy6ncAi2ESK/vM0EU8vZoHY3Y6csoRUIEt2xG
OSmTGYxw6mQhwqxN0c8oYBKc2ZRTgdnTT5h+LdCjBYg34W6/Y2E9ow8knBpTUAsf9kEwXbAisTKl
7ZoRGWXwKGMf4Lngwzz1UBWF5ziHveS/gd8bNCLHuaNljST7dc2EmDsggk/0KaciOuzV+cqMFkqx
U9DHMWancFFpthDbC5JwqS34u9DP55OPey55/TGURiF1tCfqJFg8wwURuhusnGXocHvLPVppE70d
C/dBKY2hxUZ0ZG3vo3AmL6zdKujbCgbKm3FUUMFfytk+yxGSeRZUtIGctOyngzrKZvxm93HdgFDD
rgw+Pwlz7OPHrgcT51C4vH7x435bmidZOOX5ZdYhrkTD/WUhvXHYK+LDHf21nk0+TUSMHzMckPVl
aNiXWzBIizgWUgOQNFf9G78M1YVJw2Vj7rQkDep+VTk5luz2BEyidZG6Y5W2fuzHQRC6HJ3c9Urz
GsOsfc8TXiZRULuYZP9NeQ9lQAmWj8DMtKoHPYj6ogGkJGAXKnXkKWgNCu2P3nIjiyPNlsvDv0G7
bAGeP+3+USwsT/27sg9DzXC55ZvcuZG6RgrWcxmVFXhoXnKUVpHzroK8PIDKCtrCI+5o4OAaxPeI
f6xty+wS00tYFG0QPydBG4Uh1jvu6raqGeMj9ycjdHZuWshqodz/nDamiYaZpVC6zE340PhKrPx3
p5lA/CjbuioTw9ualofaQTzvRERxbSeN3wv73/nvL8yObYD08LH+LNhbJ1uNTMLUcandXqA+/6Vp
5rEBzjsImLbosHLqKUS7HwF6HMNFtzvzIpTXlW/Qhfl1kCChJyShhB69x9FKETO4RC9m+pOXHmOo
MfJvcC67dG/7xcQs1Txr38Kl/TTPZe8dqIWB19SmN3TUUhrAFyMNYxewIIzT0Z9tzdzNvGjtg/rV
NLu9/HPgXr7FpjTy84jnHjwIEGVKhvuQAnRsyV+D434UjS+rLoNZRN8MGoqR9wgdpB/76FmBfW05
Oml+pRvvQ2ICeXCLXvCfrhI8aN5ZffOMXaOImYt/+UufWKxHi5zdioDT9XD6IdyzKIyvLhOTKjsF
LYKoDehxX/gxCFQcrQLINPn8Rt94VXaN/i85GThkEOhY9y9tFtijpYWmjtNmA+GKc0wgUDvPMJat
A1LhcTs0+m+TV41h9mCtPAN4sRFirBmmig2m8B0JxUMmZK0IqLjjm4lPo/HjJ+1v3KRlv2sZ3ozk
SJbmCIhF4W8qYbWhK9vz0GH5m5PvHkQK1l14DlTbWimPtksQ16thzmfaJw874ZpIm6nTOFGpsnHL
f2LE3UBcV8fj6n9NhzhY7RLm2JSyjkqcrPy7EhFh3KWCBW9oXXFgrSfztCN1MJNwDTOvWOPPQLmy
R1sxsn5rqda/fpsGHd53fsUPVtL/fvKUNjX9XfMxB/HeYi1PE3/H9aAZH8QWgrQUO39GDEAYcBhk
EkAQM7ECqs+DnvS5Bi21Y/RPlaz+cBDqYQZmz078ZFJ3XndCgYhm9q8Tw9r2XIMz/ZtIZpgPJBIN
MsHa3ntQqeGQkFczcx2AqTjNTUBlz+oVZKm0PzlzMcGJ853STIGduqyOrhjBfrNYYXW1VsoQ+6Ys
9rN9kmiwByezSjfHx6qBgVUOvdCewd4A/zs0BUnMJA+EP6yZ5YECV8IGoiEEKTCF9fxK/bLQ5c9s
ZXb5woKDMlKpCccRCHkbG2J+B5FDtURClrnENn/mwyjm0Pxkr4rQOU+BqptwOPTO+jDPdYjQ8KF7
XOrxLDCepdhEoRXjuWvha9QJGCaw2VpG8qQKeyrPHkIN4dWMOPY9qBzTH4qkjIYB+KF/EJL4Cl7V
hOTI/t8WWKJDYybCrM1BlGyUPkmr+R2Twpcd0YRd5dHZwgH9y1KLrVLq9UGiV/yCSLwvQTdaXebR
R/6Cg3wrKc7dD7UHVc9cI1rKQbVb7IJ1HNx4LO80nHxsQwYQuDWoLSqM21f9G8q6/zXN8UhlZ18a
kWwkAWALbxqqNmaxjmVQ0/qKyj8UOwbQo7Hy0aKxaoIlSKDbY5d8tU13YdI+jh1ZoJ+8EePjZdEc
5q7Qc5ds/veDsi3nTnl5a8teaeP8cfKmBaXuzQkcvkuBLFtLR+yZexxypIvl7ttc2eM9K5ndLH8S
2iIAH1yflKGdV2wqtSsxdEwzxFwotvRYt11T7cd+YHZvcg3hXhlRsPRdDKRtyJSCc7SdVFYOwsz7
951L5AuBtffloT7ohz65rC4c3PjAW/80oMTr71qYCo/LDicIPu/Wk9YPNkdBw4WKLZDodB6wv5kE
y63KFzJrilMO0IgOXdNvjlEJsUvO8w9wBr8OVSR7YjDGb8Sz3kPxH3HhmJxH0hxhGB4Ueey0FouR
w2n4BvmMvSFwdRbdcxhtYI1/yygxcbVxUdQhAltj1t4lfQ8qvXJlBuxXczL1QUJj1Ha0dFOL/ILj
J1kfgz7RhCoCfWfo/4aCKiqZxxlb69DaF1S8BX4G3nfeSFBpkY3wXPd4+J9zXRCWsVYUQHI9T/6P
8ow6qnOdWXP6OpHcQtAHmVB6NSHuX4riQ+Mppc/5ZdS8GNhy4HhBSMt/3FwRpNhp8YeHy9gR7zhq
LZGd2n9ONFBZQo0HdXUY18Y8dfmPNoSrMfp9nowo48AAfSK4dPkBZ+JuYBb+grr2Lag0UYlNJeSS
odtW8H6kRDktKbpIgEjOPaYHxxi+W/2DEKospwkzoGYxYinMzHAlwnPBPHYywe8pgWFRz7uOKZmw
3ONkjTYE7uXRl3SC9TZ1h1qJ3IN8eY4/Qm8I2pI8gOBRiRZZqWDPoE+h4LmgoGGJB/M27A+K8xaq
UqZrWmttENmCDKL5Oll2y0zI50rL+5Q2jwAJ0/bNq7Kt1IpRo8p98kMWg2m4v0udZDDPLsY/eqHM
9L/p2RUjT/98yl7Ob0KbCYD1fZbSv87IB0dD2fwZnVcLOJSuuxztqdJoIg5dSq74+7KyKssZSFFT
3b2E8ptnFMoNFKqdGLgz0rl0xArlRl5r3Kidjqf3itVQZHt0ZhL/9Cd0xBb2kokp2pkuwmo841Ao
WpHgq34D5O76u0Elp2yaBzFJT4xkJyJWvq2Seq7g7sEIiCLm3kojDXNPJw6k9k3MJyurx655De44
C9+zke/pklS/qHetb1jo9BzY4SZeo3VPlYZCKPr86+2mVw5ZHd7Ry14GwrzN5Y41PuT4YnqDnmsh
NeHxpeEJYJun8FKi8RHwDGLSJaBRaiinHbwe6VjMn386YR2HbLNpKxsu+Qi+wsPJ7GwWCat9rooF
BGv/w5VbWK7cO1TOaRS1nUffs7PyHtxtKkeAmkIr+pAmzUjA7JQVBqCj9E9F6Gjiue6W+pXMq7Px
iZAVIIug9+pmLcQtNhErmecF/tHHF/mNhVoQPpEJXuyQN++Ds2BF1kheoli6lqKp+yelJ6o4mNMG
h07yyIaryRdXgLvual3HHricClDm+BaTbpdnmiJg0DCMqKAOD1MkxneiXADEbSjArt/dn7DloYL1
19rsbj272A0sAwcPcbeR07KwgWQvaoiBABYpMc9NdTznA3ySO94IbqFdIwkLSb6Q75LrNDF46VAU
DqZufsOkhaWvwnQutXgcn2CxWBVf7RpiKciW2MwpReAi1hF43BtCS4kZ3Aw4u+Z6K59GVF7wU0gU
2AqTS1brhG0viWfAXFSt10AdSlezk1/3ANQzOdEyRTpqVU2fBj6+1PMHa52I8vvoFe4ip9eAJhUG
7dCQ+B4Sg9EAon8fjgdyakRfPeiDoPX8NrfdXY/rWjryCsecIdPhpphyhciBcJpG5pIG5fu22iXP
gC9gRrEPc70eNcaIen2LyOiNyowkgWE9T/GBXiDJbn9dGzTy+NVw9FY+DYnnzxFmKUAVAUx0PJ+j
MIQ/mm7bLv3KmDrhABUll8R78hy1Az8N9A75/ZILT+4w+cSv20l4/y0XjQp+QoA8++qctz5RDi9Z
x0B1ootuEdCKg7dUBvJK85TpPyhOmoqjDk7cAf7n+mq789GNnEh6r88V1D/tCOuHLmBByjtzM9SQ
M+ZsZNGklQZAQFEDe22lEN4EjBEs+jNHH4HqDCCGA+QQa07FlKwKHc9ztKhO0aYlED9X880dHISZ
hVflWeskjgn4a84LL6TFdIPtL2YO7w2IhE/2AIEH9Ab1DFk1brNrOSQQjOzo3Nk4hcBvbghxo9ld
9X0FZBjMip5hWdwnxwh6MvTFllYbM4hoX80CBmA2DAhDEVba/d4w7VyAoib439wxW6Lzb4NGPsmq
qCQgE4IDw+f559wDPsFFJmcyIYJPQ4exS5jjBnqMlJ7dhLZoGo0cgT6YqPfMvvPG7Ux4CQIhxeJt
LXn5Z27FMLG5ZxvAkj1uF3LMpdjyiOuq3EN/+O6O/HT2hKfGO/LJFyF0iMzmJhdKodVYPXTE8BYr
DaGRcS+ViXEvtaWIqBgHEAy/w2JpRCQupza4fWGOU2IhtP//0BIjlJZY58r/yhzpOmaN1883x6XL
+fmmMlTejlWe6bAL//zM5ViAfr4qIg/NX4fDG7LGs2FFsSHHXDj1mMTnuXCczjQ1a/5EqPWWLJSs
mtZfSV3BoMh/wVKBaNC+BuvztlQIG5A+xKdKuwNioPILNPFnfTYqzwpdIgS9PlkdJ4Qx3VNvJ/To
Vp5CourCAn2jWwEDs/hLemDVDI1jmpCBY0Bk/zGkHxa5Sg8vARNR4JnkGRDRKgXLgUmu2gsLQCzj
3YCPxn6FcIX2Zkua4Gqjd5jyh5DLFxNrLZFMPHj97Nf2tUrWqe0BK7Ro1+z3jS9XUJlfD8V/cU1b
HZpLdH9SVGHVYWJsAzqeNVm5aCTLw2t97Yh0+dUBjZ4MMDEOrmoGYSEJXuktEus4BTdVTdZl6qKo
1e2EOv92dcj/edrqTaPxnvR+/TdPKQDKjzpommEPlUYQRkVGA+tvOeBwHbYNMWeARQNn1f5g2iOD
iHV+XWPA888U6rNH/27REHbEBx00Hi6Uu4sdDTKaYez1pyVesGdTUxhaagmWaySd3ZBIkPI2u6wh
xQzV8L/JUUFy7wWI9GXFbTSwASJIOV6BaRrnkaxCF88xhy+VH6KBP852axCyBaF4vurDVpUSxBeV
0LXyMjpq+AL7Mlhlw+lSgdT3amgMVRD1d1C71tNUvAp+7iAChzcZgetpWT9YBn8Pi+Ct3ctscycm
rC0eKxAOF2jip6ofLiK+J61oG7tse/nViiNfRu7oz2HiMTc1lH2ZZhzpquvRk6hPWleLLxHmAbsh
SahqCK6zO1wQOz5FSVvUrE4k73IxLXydfbQf646Aky+Ic1VU6RSpEYfe5qKGTAKcL9b6A67FJpuI
7UpVTdX8uzulgox6WoJBRfgvO8NRReO9N+1qnks6PBt+1No5iVnv/WBZOc+VZEvzLvylRh5iZCgN
v3kHY3NFSmeHfWL9HgSsOxbbIfJRoH87EvBH5az69juKJyQuqe+vA6z8dq0NbBTc2zKPYnYgzSqn
qFaZGFX6ZvzU2K8USGqhblBuVKMekBIVbt9/gOnSuEjDeiMkGiCt4/pHYX6KlizcpoH/0cUBa3B2
v178NM/eSQjs5OyDsIWG/yss+ErNNl7MOge6h11KGPuCDtWojoSCTLYjedWMbVRft4XYmLfIoLXO
VzJleN0uE1wgOxSiLqjoEJfrzgwKIMGDDS1EWZQAZaFoUsPmyx6YSYmS2l/i6pKv8du+hB56Ree1
F/qf3HV9BKSdfMjDi7iOaus0dAWHMFVQXutK8uToTpIn1TDOmElxNrx8CvUK2QhkTNjwSGoo04t5
aYCUpoBL8HiGsK5CpC5uAgXzA87JCu847Pu3vi+FXf9A+KUR9dDVJJW5mLbG6qCJcKF72t9P0yA2
3Vob1iV7Ul472JsaicaLlSFZf5tURgK1kK0PFjdgEXJcVm8k7pNqrfV04e8jR1jKLiKQGRNGryBR
4ijFEZ1zDb+c9Bdj2dfs8mF0edZE2yRw+29yhi3j3HRD3GCZC5klkBR507t/X2I0t0RuYOT+3eby
6bRI8HJZxuHJA8sfyos2//NoSAJ9ZKWd04GEnQa5b1lt9Huq91D0EUnfBU833ygvFH1a4CkU3Shk
czrZDfZ5EHYEPJes7HV4IgwN+T13AooFFfXl/TxG7Go01r4Ovd8lOMSZvb5Ww7XdwyEq+qNbBXYX
ciTtUjhjtYcQYBWDYwcVmVT0qAPpjC2TxOrTavRey+VOv4Er0Os9eek5tCiRAPkcLIu+BfCAwG43
XPeaue/CQ3uVEgIDdkQW7AK/OS5Nj/28Uym1yUvvEVlJCtBaUauYtBSUkV8OiKTkLFOODJVR9kem
3qvBwQjhJV2Y/HEyWY6IYFDkfATYkMeuftYHtE0DaNpN9jWU5iDbN5Jc1NOAfseUonIt59Lsdd+3
VGBTV834KF2xcy1WShAQ26f3lAtJwLwF8MyuJ3XW0NC7qTTdcLooHI0dbaTykU89I8dmEn/GDDOy
irKMPhAK/px8C07r/e3bY9EP1pIZQn9HxTKUnDHpxijlsV+cm/XaS/JHQzkBc9zQXJAyu5q8Nlw/
bzJijpYre2ROeQyR+z53YlN3A9VRgZahKzB1sVjIvVmkKv/Ka4EWOK/xRvsCaEa0u83NUYBto+u3
GoIHPsyQiLUOHUCkdYf4pq8dDrcuzShWYLwOzSCAlvELs0FJTtax0qFDsyHHIHL7lRipmEK1lzG+
lOXRU/sVXKbrJO5sNihMJPzyvZ0fu+A+Wt75Yqz11KdX0isugQuNbs5fCrxCaIJdI/vYSSlSw0il
/9NOPxSj48uB/5duEgADq3MiIXr2V0FEndwdae+jkYbf2pFd7amm3K2oxmrNFBbShn65YfNJdVNB
tkZqM5nW6KF7pVMQDjioC7RmkZmitCyz9UETWEL5tpubVFfxnmD9Ol4xCiSss53CTNG+ZwxcfM1J
iEu6IX3xzZ3Q/iMB5fNxSNl/eTv3wdxVqM3KxLOe1dGjm6iiCoSSDUAVPTL8uccfsZhc+vO4MF/G
VPGC9o6vt2t9RcSnTzqhOjsIFV/OSNDF7az/poCY2oJyu7Y13GyWGXhf8EV0dWiDep9OzaxX9JQH
XjhAuMMrd0VkauWo9kvxApf8SNDCqXcfLZxVw0tzXL54DLGiqNovk2/ZgOyLks2Ln9ZED5d9cb9w
UqQW7h9/ti/3KL+yGNYFd+snK2aLXJWx/DKnzebcNEervgnvsR/VfrbQZAxS3kRAupdBf7p9JPDW
7xsmSktYLrqM2zCBZE+rezRMt48cfk9QU++3SV7Q/2Ro19KByQobsRy8juuzuzL4BBxMEvOL0NWP
5+GEWMIU5uSmSJyFOPFPWCQg8af1zRQ+++3W1DxS9v7Agji4x1swlUZteDfrG2lsz54bmTy19Yka
HB4Tp61/R9PM58Z9X/VFk2Jn8+nJE8/IdrV502cRysTkK0C35r4PfGTzQ21JeLgj9eJeDNki52Xb
SaMnQp1SEUZZz8NqGgY/GltfeGOO4Q8zy7tAynl646hkIPOQ1B075/DBVKxSAP33EvITKZ5stnjF
dPb6gMX6JGv6gHzwIbg95+oGsmR8Ylh8WdPre8L2YHximo4KeCjizD2EVNDdYpeEDbxYM6jbrX5c
QqmW+DGNuz0Ve/UxAWR/0KwjHf8SlEszTG2cRev1REChYedhX0brVpKDDFdYJHtK8Hm2j9WkYsbZ
1N4Qz+3SpCQT7BIgKz/4dNbI6hUJgeaRaALO6BuRf94nEqDU63PH10YsNgbwVm88yCP9liSWTg04
OD+EGk8Apj7yAKCsgEOXzOW7eY5pHzWWGiqhEcwxvLCCI+OqOtEzOmRsUN70JI59vhCzqBxpPPg0
alHJK8wFs332nSwcy5gWYjBgJNNIIqr2bpwgz5PuU3ydib21Ah4KtnZGYxHGC5xe68lh/D8PdsgE
wKj3OHppKUA/ILCw0is77tbNY029eXQLeqIWXkwuG9tFeOUYCsl6M/BS4gN11qHOWlEf+oXT7zFo
tX1scRtRXywmCsPOcWRXfiafdSt8hKOcNNR6/N3y0eZ3gZPxJmS8QshezdgINKUjcUxG7jmGKw56
vX+aihwaZcCTIABgzNICQK4ezEQrfyYe2CbGsubKix/SE32P440iwT1pZo+bSDfDwGF6KCrQpe0p
XAZjxbnJlX2iuOUIQN4nOYi/Sf5Q6F4JmGkUUxdDKJObl+dJHQWv/xL0toOlU89slq4xEjD/Su4S
fr/YbsR/PMp4PzMS9IKEKqyvx6OdEWi3wJAWed8tIxjNN5Uh4odFIoP7MaNk6rjeAHpmxASKe/x/
eDiP5dZ+4Q57yyDz8j1oIvQNRSwgGLQV3ZnmeLfosB+KpqIYXlIPiUIh+aArNsM+QJCcQ+sCYFQC
HNt1UxSl6WCfEVHDP3rYouaY9tMp22Ijp5r90w6Ip+syh7FuDAR3wLDPrRCW97VOPB7zu2kUUdVR
UIhAQcAma28Vyw7nizSLsKqGOoKlkuZXs0XpdpRIaH3g932OfRhGVTh+zaarwB0gjciVHHF7Qqrc
pfyYJjY/eQp6LQttvSmqUOQroYd43K+4jgtpYTHRT46yMfh7No33lwfHkbieYKf+HbssbZtzz+C5
D6OSx8ulhW0boDkzWMOgM2cScD0APOO6WibK7awXEeAw10V3wkOzNWOtoUi3H1V3AkICllmjXC2o
u5RhSm4PsRumWRLjQeyS3ZdmOWs/HithapzJC/rtTFmsxaV5qu35iQegVXpsqzXh5qfZhgxYFPid
uZwnZFuSejtZCGO4UxxGtTh+YsvNNOK/QWHTvie0vzvqDw4BacFO51mltS/Jrqp38ASUugjD/G28
QY8e1GGGnzh5HlBZk0HXrIWsNOohMsem19ztQgD9m9/7+sFbmKvTdsRg41ZKw7V0UpR6NkwGEtV2
ck7muwfzMx7LNOOcaFDMu/WgbwCajx4XK/MBu9iDKYNboJX2gNbJtbw8EOiT0Xybm1PCbHnX+/PN
1phV5iMFwbyq5NPCN/oshWlmJFAmxEoNbk64xJuzWaa53kDLjGZq3CEKCfPBgfAIap5Un5/+F1xL
TQHGJMgdQgNlsl/9d+mRurSiKpsrxFUSrdknnjajkzFryA0Nrr8x795mlKsk+mnqAzQjO+B7lp1y
hR6nMNizEd24vEKbqNriVPcCFarx0GujoPSQ7WRokwaJlzw5NESYwgeIgDwLONL9MRnVgDy6gPdj
oQGStIumGgdREoAyItv/BzXpZ8S7tjIRBPn5MW71tjiz04DdxgQTp2VE7I8NgxK7lf1sQmcS+3ml
RaPwwpfd4BHPQREhVLO0/xVSOCYTfeuk3pukRVA48iYGNgER5U8mD99601E1iQ4U60ahfFeQE7No
VMGwE8LdcldUuRCoKwxo3YT7VfGQ0Dy0OUGMmPd4hJ3c5mBIIbxffI/X+nO8QQ5WFAG0OoYliEXQ
Idu004R/g9U0P+vT6rH6Nbk0ujqIkIQyN6ct6wjvHab43l48ATVKxvyjiApPnHz3/5yL7EhrmArf
fsRsOfVDsGygKJ73kZ3Rl9+3Zd/FIJF36BFSYlwlKTqcXA5G1qHDJL6/ORmWQuoFDUUuxIE3Gycc
Q7JWAuZGq9CrRAWOBG7xanSvZYLNQyGQXBp++UMVQ9o8YSqT4cIs01aTIP1uP+o/JqinEoGdISZd
ivsq1F0fWLvZ2SzirlyrAFF0J2YPRCynxvnkSXCECPBj+AoqAnBVKTpVeuIkA8cADZvKPB2fZpL2
aZ5wTW2rqVdW+DL5xT+q6ej1jcAvhUsxAqUtNbooWj+13TEUdCJeG2XMNMd7Z8MoDkHF5g0GfHVm
B7XLNqKEpjVKLn+1+/IfWWVZNgOlSzQQkIiNB8x9+EsyfrKBDwVjIYR6fTnFvZmsjNcj6e9QvBOX
o6QHKfbiZjuWNWEzXsGR9hGu0GOr6kQDTutfQy1vpRpffrHCtzudOwZO/31ECiccFWBVOISjt/Um
F0zg4J9Uy3U3yi0mxbuwDzfuZthqFa17+2aZk6cdtc0g7qwZ0PY7Xn4MT4uVic0HnT4JXDdiz68m
WgGCRugVnca8Egp/j/YCJX7mjn8QynKzt1abHJitbroxNU90YqepXMVdx6Jd9oiVJt+tCCCygvjG
dmgdXtrIUPFTg6G+FFnuzjMzPJLk99rJl6Vey1kpJpVHE7BCmSzPRMurC8N/C3+enKhsbr0QxXEy
qaKl0eS65noNPQ1/sgmdCsF5Al7Ri6lSDt0m1XSSCgWSpxRJNhlRNRFDRZoYSXlo9/nQweLs9ElI
Fq5eRP108PFArP6YS5CZnjyqOPXTjlCevJDgu2BM67hKe0FdQPdYCfphMRgkuksEM+Ft6n2p7gFQ
eJbAb70CMmy3e/JoS4In7/LVtils9L4yFtsvU71otnDEJgiSG534VZ5+RwQf7Y/BfrYbSKcHYOxX
qmyMm83HStsIFNRZicWUN6c8g5qsw0TE361udMMIxtgguvk7g8oLKUjrg00WfHR81UUiDUvT8DPh
/2eyp7KGxKuEZekqpvIpTN+qR2zPxbJw/flZTKZZTZSjNRJYgRJ+vh7rAgxNWNpU1DJfXCAPN27m
gBcEF/Pj8XddF+lWYnX9Kc/UTZL59ZFgyWL0zoUyLShUh41CrlClgcPvlqcFO/eXnOPn2DJDf97n
VGi13WDf+rG+gGf3iJX03PO51LRvbjA4cl132U56GYa5ydD6jZno5VANzkVcuuUDQIkxUFUABJiE
3TR3++rLsvveuyg6lt1T0nGJQzstK6nUA35tjR4y35+Nh5a02vzXIDfSnUqbQemnFTWRiLufxyPx
BmIR95N6yo4kRALNyrkdhvUIUSzlDrurVXgXwty5Z8J9W/9IFwSoZNbbnmR30cXaNImw4fj0UmxX
N5nN+a46llDaMiS1HcYP6b3YTrDI7Id+Uvf6LxJwO0N2cowuxRvEkfSu4PIvqRUs2g0PKh5gUdMs
UwoDyRqPBZG46agTAhe8JQ+sAFUBbvp3k8NW2/nvuEJwUEZUdC6fw6NL4VMGZH0ceC5gSlsMBA2j
pDNo+IWDNCIBzz4V9E37Gjr9xkefI72XqnG50XGKxqa3AKcyA7O1F4DX0hR7J/vjqQAEh39N0l6s
KyaqO8bD0BT5UrtJDjdhuS6k+M1nZ2hmbVHqyTYYn6lXBGWP0cOmvYYPz2uThmbv/KT8RHB/P4DV
85ftG9RKn5ArGA79KWRpiOyj8RL7NZg2+Z9XHd3zjGq8YvLKryhmzEH/beO55tvs4ZTI/HV1aVNa
nLlZj345SU8mNiTkanw8yZT2B6IWy9lcDLrI0TGI4tcnkcghcwTdXEq6ZY/PbmLRiGvpPZBM7eNf
jzMjaiSRkEAGoREpF4Nr3cFR5JyetEU4LCel9HR4HFS9m44S+dXCBgoNbHvEmFxteXacBN0UqOXY
w1VxQ2IjbDB1+H5zRf1eEETdiv1dhbcxDOdOMyXYSIThoL5Pjn3unzs02E8vgw600x23W9eXT7Nk
vK9FavgIkdi0y8yYO8cTvl/M5HtlRzq+VaMp+gC2k0jlOJA5V1h4bgYCHdEiGcnSm2wiLYBwZNjq
MGgQnGLFOk6Ihesrpp0seLYALS9BuMRFi0o7kMtWzPojK6c08PymIe6wjs0t/s5bnKz9/BFjASIS
xIkC4vNcPs2sRsQVlEzkAmHLVo8uzEnjSShrqnmb/6lbahTdgJh1ihxYO2Ai/DzaMXON3vdWAv9Z
LJHTJxIXzdwixfFklEc4kXRnlFpTh0J1NtKOoUNoESOtH7pCEUd++FEtHg7XgcBUw6N7KNgY4E2I
M4v79MCIsVvFFgSFCxcl/WvRfYfHyrDN+BwEoNWF6cy/upgqrL3qmFG4fneOeXSa5OPisQVpqdMP
T/5HEOwcnntI8TAeRAEyO/14aZkouKrosJPt8AQ+C7F7Yyp316O1AwztuW6pYfM/2i1diu7j4ikD
M/JN4QNs2Q0P1+/XmLaeipeA0MhhwCcjAYwHfXqADnC7UAxBKklE43J+Lf2c/IvN7X7sTvf2AHSH
bpbKD07RWfqaFqFeXzBCDe1s8QkW5+MT2yH6tv14/Os1bdN8LsbS9YHQgf0OJXXzQgosdFhIb4Yr
O9At1STGqmQmng9Xyt22FvmBfUIt41hhTV40r/3zupmpDTgtQkeTbLizVewzxzGTY2X3NUgut8ns
acfRsQlIbW+ssvfySxwvOqxR8C2czCkL6MB0dbgVE9kP/8SojmpbfJ+ZCRLlLtnYz0k9qofq0iSX
0x91d24VW3xZ0b38qbupju5d4a3hkQiei3UErKapAqBCreHSwZlpJhUL8EFkhy/LgkPkhHuwYCrx
IjZqgtVnyMAoQfgo7y8rvCS9ZfecuzrzmJ22W/hngO8kdDo0MNaYHBn21X6+xA2qT5S1FuN1LsKG
ILjmW0SQnrjU+YNroeRuUoB9YNNgTreECBL/+Tgi0DfMsH8/4mPnLZACbzb46Un+6pyIEoXyYwb0
bAuZtTYd9wPSMCJuTRJ2+/TG8DP3Gs4HpdFUtsUdpqYz/XEDYzXlhGNF/5+kvqlm81l/YIi9jEDa
TfimYqaleI581S7SmBvZ6H3DmrFIyDVgEY+6P8HkXmH+Okw3uXAPj6OFJKfO3ntkS7/BN7mDex3r
EQNDhNFVKssWS8lryE0G2Z6/a7opt+3ACwBz2q6/XB1crGzVgFjNYTOfbYuxlLsU6xPJbfgOG+0a
mgyc0731JnDs8WvzBe3I9V+Fu++A/8uYeth5hzOylcLbqdJtgDtQZB9m6Cei0vM2uTX0U/RAhGQ4
PAlkYVp7ptwwLL3Fvlm6TyZWXNKGFVjYuNk+zMnQZl8Px9Pr6wjHS/shdqHk16Y+PwcG9m1Nz10L
xGCAGmurC8KFNC5blWfoW/mzMZEj5BZID2hFBIBQXH8z6D5ZjRJMzmowhPLo27pLrpyXg8xOuQKz
d0AuLVhbQBVEyb0b3ry7fznUC7bObZgyF2jFrg9rXu9itwVzkyYSlk+2AH9mnyXMtWNB06JCW3mQ
zjShVRkRijuNSK3gcrVfruggnKRAXNjgutEIUEJ58r+Yb0Gil+2jX0zTZRA8UgDabTcq57psSMmY
fhdCsRNjsO7yS5YrnOuxt6j5mP0KSo5zWqQoHEjcy16cBlmW5nSF5Mudjk0q6xN0dRkdn2ptpgeI
qGlvd/4X0YObs5fKc1v096K3kcDSEQBI6+bmPlTk6/z8Q7MGSc51TPB2jukoVUQY33v+5EhQ8EXL
xdsad0XYYmtnVSsTAHIa9i6Ik5t62y+Vnsi20pEgz5XqE3xACWlprNVxAuua5n/QsJCvGCjWz9CQ
mWpKC3bg6R6YkM9eCPxuudz2Lr4J8t2a2ixiaw5tS/CbDeDl8uccaQojSiccht4l4d5loIzDL30d
ejOUpd+EQ2OlsFG3YFHOgOE+QG+Zg63jBr6TN+HMiQkbFB7yjCMxE8mgHLp8Z87mzZIUnpvvTh12
aeogHQ6ygrVSChNEzI0dgJgkRMOYGa9JmdINVu5p4tzz+c349kX9B3U7b39Z4/0VIvqQmopP5aw9
K2Zv0LaD4WsVyc/MVe/fTNeFZ+7B/FCsp3+f1+lcc5Rf/2FWbjOAsqDHckznxeuHjgNCHo8l0B58
s8Ew3dbagfBHuY6+XXWD1khsn4Mo9eAx66vG4z3A4tPcZyya2HkGV8oWblZ1Q8QOTcGYISeHCGxG
X0MErGWcoImwFkDvORGWRjP2E5azDnU1MY/M5SgtWku6bHFpoj1Odo6W1SzUUDnFqYC8bT/zkYV3
IK/HF61Hf64UY2uT8zn2oQqdv0LBOjeP3KLTM3gUqm3TM/KKJjmAVBaDQhx2NpJ3hVqlCvG5uNoq
m7epL4APnw0F3626NRribi1gKbh5U/FRaT+L2Xe6TuQHBV84QxApi6CZJfr2eNsCaJVKAyMVeboh
/XO7WiTVcxlIFL66X4qg476ZFdbzuSV0/pC7A+BMAWi8wYoXJoQzWGSYrN4U7wxq/viUzP1/9BkE
zhEaOs/K7AjMeGgcVQpJW1vcUiA3MBflUVypsp3PtXmRV65AujjcNzVxqCBTwc5vTpui+ae6/xG4
Qb3prCU06tPj5nOMPcSjoC5d0RUL3UX0MvqpKB2obEEuCJgSSIOsd9zRqahmE+RegDu4aBgN0vtd
3RfqVXCdai0gvx41IuGwCHs+BnrxCtZ/2egC/9ltMxOr+tXQkamUI9ZOOfe80grR58Phz3OG307q
bqMaSvIK4vWCRdhbKq5E0jkrMii7aKQ1mzc20nK7z/3TxTV7JuC+zblelrhUveW2dejNRJnW/2jS
gr2caEk2WbogFolY0IinTFNfGrkHbVQuoBZK+vQbT6sKNOeW7tN6t/6xxhn1Eqh4xF5G8+oQbZI+
PIH2+xp8ymmH0vBfMWDsOcHV1kXVxU24rrs999Q8Z+ldxv7K2Hpw9vSPuqDuI4VMyPeuz+PxdDim
zEN9sJKCoYYWKi7bmq2cv1v9Cb625sh7laGa/flly3DMms781CI5wh+Sj80sVvIcyEEevqlCkucb
cexcvrVcWAYoIMO7kPhiC+eyVKkdQLNzi89fT0/mBnhB4LSJx/cax6jcggxnd+woyws7KVSGAB0d
VIGeN14pBkD4gvJXiznojtLpjsDxQ5MNX2WsoiJXvguqtYmZXNgq6XwvxT8Uv3dGcagVsz2OlVAd
jg8lNaeYhBDIdcqHqCQSNwkIJdU1dQSgC7cOeiuCLo26hKbhchULXUE1tG695+dV/VqLh90Jq8Zl
ibQfw4L9J+a6ZVR8GwYqWPQhwG4+LyRgv9eEqknPEp4g5bWEYo5Du9xeZHKxJnBC7xgobFY8BJx/
utG12cnV2YZFSIJOId8irFXP7HHQetY9xTbdMA0sP2tofw9zj+RKr0rW7k34nh9B+oN44+apTrPg
+0xl8dzJHIRgz1KVTSDDzW/4f07y8sUvvKT4RusFl+lmXYtgAw9gnmNywiWoa5nhwr9XZh1uxFTn
DksgHVvZ73A6H/IIu1NPxfBgQ6T1z1NhNspz5ynBuertxyaUtBIVpSRbSasAiCvEiZE/Lfuv1N6G
whv7X2vaJUIIDeOZU2iyy0CaOSrwAWHjL/HF8lVoSJDtHdJxT2pw/MF+Qo0+Goh3LIZsXv+Zcu2Q
nVo1ZuSvhhWjMSWPyxPBIKvAGy7p/PEN5Fb6AoBw8xAcBhAzqyptiwQqZrm53EGSFEomoukP+RHl
V2PSf9RbQqZWmSHMi7wilQ787q5R8iB5oITMYAn2hsDgk0EwyY9q6YcTB007aG6EfbQZJ4Fjnd1u
27WLxlJvTluLR6y5ZsiRauPb+RDb//9Aa9CsaERG2Q2vayrvwRl5DYybbydePvjth52vzkhE3t7a
2aMZ21gCNV6EElA933UIT1z4OEx1NErZJI7WtaWvIoX0qzA2Kd6GJuDX3wQO9Z49cgUsWD1ky0/M
5O/OSFFty563Do4XdHdKOINu/enjrmJttBfN/mhPyQCpYTGDHNlaIHkoeDKwSNK3y1yB2ZYviUOJ
mY6TkJMnYgv1+RK778goAswqroHlIOhrrx9i/atIYuKW/7I4fb/MY6ooF3CTmoAS9y5qyhtkBHNL
IFg2yQP1Rg8SbW5aSiTfdu3AVidKxT43xdAKyxpxtJ+GdN3PccZdpQMSRkAm6kMipdCU6bSdsUqy
tJm1Aavgl9u9d8XO3rC8Uk4asRglmB1TAQwaIInRsjVEuCyunrhgmvVRk7ZB5pB89P4K+uiL73/X
QhJMkr1AptcH7BnaCA+Pr+29GNzdl+lJOfsY9BGUnMEvI9gnRN7ON2QmE6ywp6NT7lumVtWFPzod
R777Wx9gDtfHRFqEBCcBLEIULoV2vqHA4AcBRZk672m/1V6G6kw+D0fBRA1PWrRKCiEDGRmHuPIA
s5Kq5VdTMgN1c1CrTSYRBmMqV4Fg6Mbn5Rt9fYKE/Kwq4fqbmeR69MVcEYPaInc7Ycr7qLzbCwXW
RqiPvS5ExWeRJktBpbkbwVTdmtR9pYwmXVq6va2W+qiJsH98DkCB1everhVn+5NrMrohQ9TXBshY
DZ8mF5GY68sS7LpEeCUEPsZSMZPhumeHPmQfnDrD/SkRHlFUBX55lV9DRZeFnsRAT2Es/tNeltjL
seQGvpAh5u5PKqaHIXq9UmN8Mt9J54U9c4G4mL+DDSp/o+l4ikWPe+3n7WE14BerWtun8E+9pGLw
VJgBxUPUl1fxXPC9BpnJ8LAB176FmNyKM2AKysReUfGO96p0zpVpL6Sy8dycv1xIfKauZ8qe3ZzX
3I35FmDNK8h4P4TOx7jr2N/mdWfmfksf4xvZEPVui8yST5QP77T6Ciyfn2E5BxygMHdB83kKXCou
ejsf482FQkWxm9j9rpuNz6+Gy9IzRlcY6aHLe+cHJ4CaEE1N7LAqwqYSJK8B7Gc2xAD6yjwYOb9f
8JCeWvKsIBGsyf65kGCdKldtAXC9cEEupaNgWgVDeqKsqb9XvjbzCVNO1xuPdvZ0B8MJgCKdBZU6
YfHmM1qjzzzZovHFwUshR6eYOkE5CnphcHUSeM8OOEr2lWxDY1obzkBCDMevIX2n1wdm95bLXMpE
JBAG2cMBT7EVbarS4ZO28t64YziatF9VUK5bAXzYOsQ6uCAnjOmg1OwhI7mueKs2Jz3MyYhV7IxE
nbX6OUnJxgwlaiSBPEp54SXFUTAWLUE+4ua5BfoIQXrzDR8/LLX6h1qdqjIp0Y4mGXu5f5vH/75+
ztqxmCPxXrFo1/GX8aT5R/gk0PcX2rK28ouqqJ+BMT+o8EAagvIsD07/HzHCC71gKIiYpBlegAdH
Of1+Ids/y8EMmTuPHV8caXETRbny+ug9EBiICOwes8RNt2U137FR+JGRPS545t2kncLdLSQSA+EG
+OxBs9d6tOu1Ian+gfIhrLFcXErxJqo3t+3riMAxR+dnOiDTjBPFBm8mgM3OvLYNEk7hjcgu2xqv
8SG4Sk01cxbYWL2JyZh4ceBXSWUCYV9gY+TOsB2zl8kx5Z68GXHHzEHb5sMumbyQe0gCMUJrWF+o
W5oGbWnPP3SnBDtShi41T97DLrcrlHXPJgN/qSGYr47j2O6WjMP4O0tV6GcSLkcKB9CIKoRktZXw
dlK4KEmEm2kfYrGPQr5P1z0f1I1kfobxUkHuO+UAAabIQhjCxbrn+8roiDMZsd8a23e79TAvUwpG
HPbaCgBAPy9pxfVZck32JHIpHeNDkBsqzALbjsNcMHypcKykxcbLCBssKqgI5tImhDugMflpeWZ9
Yr00yHEwvHDOlRY7V2KrsyXddrVXQYnIZ6+jHuGb6s0ylglXRhfTtiZkErKutYRmzvtPazTF9nUQ
N1q59LOsm5demsij9GYqSE5U8c5+vFnM73earQHpzLfBkKY/v1+eRYYg6xNOghw64Y7ew+RRQTKW
t8rB0ze15WCXhkWTK6KhPtkOtFUI1a2OImVdT6GvpV9vITqck8g+/gWC/XUD7Zn9LXhSzUSoNzWk
cxBd/6AkdRZzqGuSk37yN8cwDfOwi/3L3Ypihy9CxBeiIq2crSeeicRMxiGKU3oRT6Q033LAni4H
5CbWRPIotnOZXCZpqfctDtaXVQSG9idZqRXNh1PkgyKb0Py8JLkuqWMZadi5a4QanpDx3etT4pJy
TFG9Z6Vn4o+i0HAkcLFoQuie7gltfxsaCAgjnX9FWrv0mL1dWyoLS7hQn6QB3ZOKesyAEaldCceB
5HZ9RiDlI72ZclrNx6FH7m9r0DFnrwpc4LBbjUchXnSHz2qzOvLzrib6+bHwsY4sys8+ay1lQFQk
wQZq1C1U+cYMlSGOspr8jdbcrj10vKojZ2Ldf8kab4eMSVWSDxcOp3I/S6UpvmDii8CnS7Bm8bvw
rKILcPnnDi55cUyI1SX/LfxjV9s/Br1pDZWgtgWFx9SdxPqGR1cfl5t0nXDWOEyJe0CgALr6Zdy3
BlMbKH+wxX+DILmHLIaCfl3waqroQQr8esFTn+AtcZp+m0F6QURg7Wggf9sBoQeAX3Y52zNduaJL
jBIkX7zLzNz3YiOaPq34wmxzU5LtK98PFHIQhIv2kOZiE8uj7d8KXmp/IonPz1FXHDbfyQdFUvR5
jSd2JuxYHz5F3eXuuBjmRs4H9cvYse6W+PdFUjJtcW0XEyPkDJl1Fu3oLDsIJnBuXT6+w3oXSAff
HXUjlZUwOm2o3N06KGiKWKeC6vT9GqcctV9IjNoTnicj2PKli8hREIAmadS5SFbmDhMRxtEhAkLs
rJDLetNIaLZP/sNdIgrS3EAfnZaWa5CbxK73fUomUGb12QMwCeF/NWrSX9G4MoE6qQUpEesHYI7f
GR+HYDw0L1GzITSnIcj5el8EqMbEU1kpKZmGmKiIZCeBupLV7QaiSslimAKT/ZwS/ZRLbTj6Uvl2
Dyd+EJiMfI72W6aShpCvGPnysG0iqPBzU0Ahfggqtu6VSsn3eoZwfQuTxRLBelBLktUHBCPjB1a7
aKpMh43dUGjrhQrUoBb/xrGUrIIcnNwJlNkC2wXEEdD18Y5+sdWerfhoBlOSDL0iJ3eVhr3/1foV
/9RQ7+VWKvPpbRkWj6VWJB/OyTKWRApxK4mksc7L7egS528q98kFmyrTE0hLuFO6T+SXpgjCSIGl
X6CUxAZ21bUFCj5Fy96AqhC2vRYXgp9BO9dlkUJzCGhIlLlEYmLF9ONfAi/qlFhK6py3iD/DOOSf
bIdC/SZSwn1BD/iuo3Acm45XfHbbUeRc7mVmGT1hBe/lynYKLrfKlwfc+I36t1+h63Uqs/1MgHh3
lXNsMWp47UDqFYof40yhA/h6T+wOpkulYUQH5lkjIorsXnaSl0LgMeFmLhubIhC09kDxSLzVd8rx
W4r68jYUmebXPrzeANUiZ2zSp5YAjI3k7F18ci51O239Sg/7CN9GbpfavTcJMT81NaIBUjKCg2aT
jFrk+iMRCLwP2Sc92EYzPJgne+LSpym2a9r4QJ7+VGXyeh9xSDQ+cV+kns3UHiRgQSTQdgs/jcoL
x8fC6NqbLk1cveR2tTJ4T9wRypMjpMx/s/N0BULUCFYPAzrNGmqyOfXusInXoLb6fTUOIxHh20WY
lCyGlw2moAIQK0RLITCdW0GMbQI9G+K7FceOu2XoWL1xas5j7dWX4Ge2ZDhfnRPTZL6WoUDuYZ7s
MKQuy5b6KPur5F79N0oa5t8tv8MESoEPDLGs8qDpxupgDH3/vI33J1DjZqgDN+grXANYCSXVu+fa
/aQMUo9iJ0ee+vGXigZUf1izt0+ivkg9SCXpg9CqDs11Fg+wwzGhXdDwCG7b3bJn6ylDUCOFeCK/
x3e/uWFgjQ5KlTTpQst3nhT/5vtyUxlm4AFtqUhXq25WBjOTWyb2Om2XR07vcaHbS84Hkc97bNqZ
cN4FL65mhF1+9azAW4L0ECoFei+UKw2C7asxoqEgYXTJJzpzs13lGGq93Eo213BYn+D+Nndo48Fj
VAE7wRQL0bJhFKSu7xzC/80CBEbT3ilw1jPjCSpDYM8DuZZCTPPhva6UM3FhERQXpGgqzmKEETm5
b/ACrOdKt2zM4hec2zcc1DAWn/YbJtQvpidclBleRWXzrVjRIC+Ervy5SnVFrKM1rLj4C4SzjCxH
3CXh/N3LxyTRAWXXzXYAwukI0xEB4j8mm1qotmfc4dkGP+I+23v1LM8Tbv3Yq84GMui179WbJc/6
GXJfN7QDpdZYkLoR1ZMYX+2hFGVFIGPjcyow8OM3DeZ+Rm2tE3DB7j986y/8jGU/81CVNtVSpo5D
PlxGy85LSSPxVH99n46fWxbZHbN0WGshSgvLK/U4MDU5UHALG090ID7RFZhs8bNpMgT7a7MihYQs
TTK/D5oiI89VlvNbUlmN902dcksKAVS9JeR3NwQwwEs1PiZse94axrUsZKDr5o7v9mLpRvtGtz6Z
yIsnO6kmmn+jlZH6Mnx+Ap/wwIpJBlUotKrX03ZCnuu33oJOlvbYcaiaff9CWHcMZvSHOypjZLTs
eGi8qFwFJP/dtAAF0A3UprcvLKdws5sg69yxy7Zakr6M4bXtn9s15JhkO/IiEMnQE5Ntm4sepQMG
JG6CSk/jLM7NJ35kLLhlLBo+jidA4GJ/hYHyeyer6T1L02HvfVSGb3dVERmVho+KAyYwIwBTwuIA
7kcfSnXX6v5kiq2DfcZHccrnUnZ3R73IpN/TLjPH0km661I/wNadvEyc00X0ypyP9yq2tR5CaPoi
HjSt7pxArkXvQ6xW+hFrMyWyUfBzLBd2OQsJXrjCJNbr7+Bvxqt6upYeLN7yJnPjinJC+z4YJJ/A
yQs8mlIAxSdWyzAJ7+5I/xGC8X6Mlz4APXVIoEpdgrIMiyFXkm2UGK3u7S/RPcr+Cagm/6Dc3l1A
YGB/KtiURg6JpH6Auyt06ZsRdpyvHFa3I1bUEZ7DbovVg2Ya7iEiINc0F+iIaSqALn4UeQpi0reK
my+ODaRTMykSfoUOtS6vaHhltyh4PnMz8WB0dAY8qQYGBG+Z+KnxSDmy6XVPb9kX+CVHLcIjVWTj
bQhXArNZp/ezyTVRKBK1wGriPJlc1NbviWywyF+RFNwev1qU2jZh59lo9zLwrguTSeCzSDQBFXyb
U+DnthgWJkc6MIogRX8wwoglU7Zb7KS/UUXJngOz1pLMDiS/3td+Kxxnd+Rkva03pdpq6juXgUX8
Flk1plsKxT+aV58Rxw3GMvKhLq36tnlLk//DQLsvFzxTfJnLJ2uwlhPCsF//H693Uq56/xIuhzNK
6LVLY8ehJEqMdoBaWHU5jCcxb4jB4FM7zY7PTju+MUpG3OD7S32gXWfsj/alEFIKGKs4dO5bpDpU
U8NgZ7lC0g9JU8x8LVGLpP1pWDdhimXJnx41k6qRQ/w+vhDmw6nUNb7zGD8sm6IDSg6ZJUiwpIkX
QUSGi0ShgCOrBaAjqauF/SPCKARYsoG593QUEW5b31BTqtoGyPXOAOu5kRkk3cmM6JLd2GBERlN+
Z653j+5RRqVEjbTmEOEVcPD+oAyxqTwofZSgxNyhuDbkwN0Fe8n/Z13+E0IBwl3RVXpj8l60MFNs
46F3Y9/pX2Jmnrmz7/nivjA4sKnZPmlBallN0vu6KAA1fEGAX0lmdALHFnUA/yYGBQYxzoXy8PbR
8khSyjTRQnXqSNEswqgx/fYmi5UQ/BHPySYiD2WcmVi1estQxgZSk1rr6R4CVdtHazR1zfmXKAkA
zsoNtKyp5r1fI4aUR5w/9uCPoxH2TMp/khEgoMcDrVDetowimnuH60TGxvwL9tNOXKjuQ7uHzJ7m
3dLQsfwyeK9EpHwsjVZ+xugGGTptYS7orbak/QGJP7mAfxjsW83W5nqZYYsS5pMIj45E9saCt/uf
HEZdFAp31y4FcytlR46+Wa1zL27XQaG22fCVgSlMMsGbpTX0eyOdBxF0CEnAyUGpnMxXAO/Hk70c
kkBchUGbajAByJKoE6FiNgTfvYhyQH3wqyOgWr7DkMoMfUPIgUW4yQCFqtzINLRJ2ZcqCgwjf9p0
ezOLc8r8jex+e1hD1WtJRdzTfJan1tnczVVbJmW3qOzNi1/B9a7RUxg0ooCT2kJg3FwwqzLAgp2I
toxMdFs7Nv2oQl0SSIegAdQfki/UxWa3pGNjmETetUZu4bEcnCgnQcO1qkF6/IVZCAPSIGqEYXnE
QiDnox9FREu/lD73E+iX4L/8LDKK4ccIL4cuSu+Z/0+jscwXKvZsK6ORmv1k20rd7xgKxqaXYJC3
dzbrBDYti4y7Auf23taPkHveJbQHeB5/oppjeMbx5I9HE+kcGYof7yDeq6yf+6kRiFOaHckB6WDl
L45346RukOmu8CmU0O6vap5cvXL4KBLr/XoyQ496oRv2PsgWopagXLjLeaLjm+ltrQANzmRaB/U8
pP2McHYNbo6ri9CSJwO47MtGS5O/+7JG8833WTV8DlynIiWI32j7RN3LZ8/z+yWu/FCDe3F0UlXm
OQXcuTNxPn4p1FuzEzl2gk7zMpMI0dM6WEHVxT4PbdlGOKPQZoqrBuX6tfz5hmmVOw7VXQfw1vJd
4TvbwjiHZ6oHptSmq33XzYngxOpfbBW7l+l4iHpAntxQQt248lu5/ExIjS37d+cKD/GO/lhxaimC
KHjbiSOEzh4cE/yv//lYlZd6LdPU5r8mwdTXyp+4omzdOtT35KNjZz0VVZ3irVlOU0rB7EYu73nd
NujkzCmpxenEqfqDnkRbNe83uTvh2P9oi2p+CyPrYLxPViGC7DaV89tySNEE2w1+y5xoi5PqXjCc
JvQLjZAdu+ARGOCluKPMcWgN1rdKode840B1BVWzERrRjITxDD+4l7/TvrGG99h7vhu0yqkz8kvo
9B/clR0VeAvb6WxHLWg/SmDSVvT9ktfCqMfgApHwGaggfYOWE24LX1PXx9zb/fnIJCwRGkSP9UTr
PrdlqzCddDLFIBc6GCGUWt7W+MkHrBH+tJcfS0l4wHVTy3VTZX+RzsA2pdV074mstDGEr3ONOsyu
rxu0El2MGZ91FIilprA5+3F3YhISeu7kw2ZhwZURUwTYDx/nWGN1KWIhQXHDllGE+D2ydIO4g4/Q
LveUjkMJ3VajJ7/9yId2pmyRmxPmefr/VPGuCPjIQRo+NK9D776drpMU+OZGhpR9MrZSboIKYWM7
adLRvzbnKrR0aotNKLc+FdKM+mFGib8szVd2u1Rmz2fNdHk2Ot4+5tnJHENYw6+LMTtrHJ0eRdnz
rMIQFFwpCpmsQHzn5ln5CMWcMyiUI0FyY87hRItAVuU2ArNpjPa3bDr6YnNPVBBy+NASLv3DZXPC
uBHzlgPmgoWnHsj2krLzNhkqH89ME66/SLDxVxeVt6A1f2+iSjGm0EcdG+MhZ/I6b/QoLwd6ouhc
6IW3A1jhjZ60sZdpt6YVKhE52D2oysEE6EpFOgAsDIjHk5pKyDYtFW9d+Rm80i1vAmUl9IUNy2vy
EIJQEAz4LCZmMF6y+1TZshjHWpdkTm6M8yRoeUhx/rFJqgzCuairQDXOAcKcdMQXbcg7z4KvVKsP
Kiaxsq6qnMTa1Y8TmO+2jbBtXrRNp+G/jGc5FSAqHPw9ytf3aXnn6SncbxNi/plOlO/59t7O7l00
ayRQihTPEmBWhaUjOHRpCm7Gtq8qIgFgvSI7hMKX0ot18IwOfXa5kH2oUliUxaciax6S9pDk7xTo
YcSYjLXuYxnbTZRjMiTq2wieZDYxpcOQcBrG2Ulf3Wcp0svyubDZNr5RPhYorKjwD6AOK/sGlZ6P
yjGi5qY7I5qtuutoAxJSgbErkEP1wTBWWc/scFYsxP2YoOwOlcTEvKNeEithWP9rJ1k+5ba1HD5H
VdnANpYzSIDWEVa9Sh1PBAIA+wYP2edaKVq6pKvDa3iPM1B+x9OHYvauldob/umLkNlXxfcIg8RL
mmvzqVpq3jQ/QfRPdEUPOFEzUHBi6+GT4ybQ7reTT2n1VTuZHbQXhH/jAQ3yQMZC3HNDnri9H6nk
t97KXKP8+/GblvLfyOeDtzA79FxrM6lfB3SRsr2YjqDPgbAvTrKzVogPTeRFXbl7z+2QAGlxXb+K
Qf1Xatik9sMaU+viBPnybSSotPmJmm/qTwkmhHQbhMA0iZjj78tzdKsIHZpyadAf6je5yJMWjCa4
H7DYvoTgigAZhVY74VS4xXNSnQhiex5/Xl242nVcnakwMp3iSe43tPtcLCa5secMbcWUvJca99GG
/ZfqkkTNSS4RnSAGclakcHGlnSG0gM2gQ78YRMGryozIx1OBTKj9z6YEEYL+fJy6sZCTuSjefsNX
hDwYXRO5k0P8Uxc7DXS2tJbUEZ6y8KE+pCqzYBF4Hapuf9UzXaTuNWfW6jYEijwyvRqI2IJsTeib
54mUVui81fdeeLpguwvEKPG2YdTPvkgecALvn7k2yuxItqKK302WGBrcts7tMT4MVhenoHfq4R4e
myLkZxMs8RWQIpeVCGwCzWGWAIIUlDYYJ1IzlDMxZAU0mj5l6axfgbCYUmxWNRe2iIkeSve2bMyo
OCgrMPJfhM6GTXUcARFBSm1DNzvw3mHTKVfxjeSz40joosunkdPncS5KakOdfn6yS6adVLxTGEsm
aLt+PDI3IzFk+MbKJlPQIR/V2WGpTUvcc56nu/Vv+Q3hThPRiSvtu6Ka6Ixaz6LiXvLRHMCo1NWt
E5Ss31aUM+nOK9/ekDfAeTreqo6Xg4JFQ3j6dRg2fUM30lYWDilZUgaoQ9Df+YEC3ltCBbDld7Rk
a+JpnKFemq/Q9h80D3EUG73piEjjN4iFsyX0BSZVYWCxxjPvzh6iu7OnPggwPuSWpeQUPGnL4Exo
DtgejBL6eJmM0YAL8dCWtY8zbYlYlXzSRze9AQvLJ8CXqWA1mbb6A+er3S1bZuO+ry+kYackNbeL
gXuKIYxCkpt+xioKNT7yPrWG5CbDj2MyXus7WIB5dHwFgGA8wt1ExOBkOUJpnknCKTc7ylYUCoFg
Eq+qGPjXIZTczyNQIPQkOplRsNt57ko0fGhCd3yhW2A8P0IHv5xpQLrfUgiNkPPttPRiWEO3ml0R
By4s18Hsz13Uu/lHABhN5OEetzs1czxnslngos3dpum/EXWusP7qvrRrVKkZtAG4jSsGwzYfxBtc
1rmShLYFl3F0dCCsSW+vKknVKEnPrd+den+AjIiVKhXipzgJvzv90uGcI/FWOGc89drm699XLyM3
MN5vBFJK3U1jtUdaANawWkDB9xhKrS4VjD0o/lbeQwnMWDedoKlhko8bZncvldMlGR3O2kPrBaWS
sb/9FWfnxu8xwamA7cJzmJX184SQPd7Wf2SUA8fbHV2G1mjYaobnkHrnhkWnmUo2sX+tNv420mvm
hZr04zK//7ZzkDJUelt9L2cxHUsuWSl/OR0bss+mq5TlXasOFdBiN81rHrqZLPda1bhqN5IXLp98
87qX+Ew3pTz/7haqMu+0Azm7wkfD4TMmVYVpkQ+UUf3P/4eFvh821WsoMpAAJm7+dAgnlmd4kwlX
d1PjLl2HPnfFTrhquIpkJ2sCFoQwuBfb8S/jUI4nNgxEf1XkmWFhJW7VDzbPoWZ2Ou+jSJCjcczV
BPBEaTy+HR0YnpKOuC54EndhlhEh2j61K2e3doMHT/9/KsfI75PJGAO2BOwEvFOfcN3b9NMTSXO+
T0jYa2PerQ1jPlq5DOp5BirrzoR/LcQfEFC9D8G2aL1sHH5dopOcpwa2QSZ9+zAknoMa4XxLVoPi
E4bzn9qMYOce2ODNR8dhlSLTxGS4R7hGMRjS6V7P1CGGH4B91t8W0XdekDeCsVgqVdM0BzmQqB7a
so8r3Bw+W2R3PC2pv0+pLKyxfkf0t1D91k1nxENeCHevyI5jucprucWomPU8bD3Mx1Upk0/kr45O
wgKw7dlJCSm4jimHVBzMo1RmZ30vC3Hvl6J5wlI5GWXOX6fvI4x6B6pQKE2NPst4BPjfJuFFTF6t
AHs0TV2O6pdOQ6uYxBMjx494bGYWvteRyd/mPFT0dEUQtjlGptzPxLTjMwaHAg5Qzp2jvmYZa05o
Ravov8/7ziHaCDH4jJdceR0HVK/V652kG8iU3K7ZchW1zhI7vpvY3xx9eu1cdh0DfPlLWeWAXNhY
+um/DdFkMY3obIL+9djlMRBuiuUXry0U7BGaKaFLgVe1+CcgArscHlOVuCLfOQi2DLJ5N27jCwlc
Vbk1EMfKIAPLFY6L/0YATwAERs2Mavzo+bQ7nR3dH6q+XzV77EOscUemsH6uRUtrPq453g586zmV
+jfF9V2VTg9fE8w9pj6vLQAXhzQNu3VY2Z5NLUNP/lkxTqpcoVagHhWBzGXUHBAMnfTUVSB69FmW
a8f+GAzVtItXJJOiDqjvR78WoslWd7WGhxeDNhBJTMOgMK9+xGQuQ1D0qoldzXEtVeRB4TBdMx6L
wykPIYMMcym70z7vhteIxSuPUT5egnT4COBIXmCFHx/jWTpXaS1ZpzhBV7POpfQH/g4wWfqo6XIK
RtftsNqMdtogo0HaMmzfWMZNkznoLimFYNmUNVtPpgQh/agny3hgreavoJkxJGz6UTbIxMWN6Umx
HC8KiBexcrPJVBRpkCgwwC4WxQgJUjl3uXpFJPQEw9Ye4A8YEJsAhBW8LaGP5Xl8WW7BuvoIlQ4q
WfS+A3YRk6TPI2UKNrY2Hp6XNSfnlUlEUfw1zc/qJP5KFJ2lm+U2EVYki999wVq6QfmQtGmrpfdx
BHJcwgIHrUsSrIH0XGSJIIxuEY3ykOEIImoFkUMWOeI0fOQsChWfiOE8fJlkGlJdLv2vujCLqMHU
cenbLM9vsw3FahoDU4nIkkIsTAAHvaJ4/qStNSWgpbBpTR1F9JG4Yqu2iw/jCMkWzPXTixCGjaAi
W47+J3mMxhPP1vJBjgbn8vAbTkTA1QEAzviaoqnE7EypIUmRGO/Z1g2onNA3s7O0uSoCsA5AX3kH
DzlNBkhDkCklU6IcBmV3oKrDPGlr55mxckcs8b8+ZaifXJOHCHj8OR7q8krMq0kd1HaBs8zErJRN
bzbmSrKIEZFusuH8lAPmfeo5/yI4spd0iKURQkp+SEKkLdCtUsX0IpV7CR3PNEh0hD5EERvFTYxJ
hTcnHcict5sMJ6erbdSc0dnfbVyPP7/6vfvZpd/FjhCJ7l/Xg3ivX3PYifVGhA9HeL3lbhqpSg7O
T1L+JZqBVISq1biJd8hkiy4KeX2MvFCUytgoAI7u2A9LDpcGpQNuhrD6YR2kKppMCynh2nJ5KT8d
EyT90AfvUOt2JorQZtOZiNmZi5nYrfOONtCHSdffvH7MvAgUuVKToekAv1HCFTjwSfvQtJxrWTXl
IbGb/CY4vrYglaGPbHgXHqAYnllJPBUtb+dNDsPmvokbGtw5KycXtpFnoV/v8ltBVvDYper80qqm
W0dcTVZpQtkSBz1wsT+Qbr9HIrmF/gYPPh3Tq2XuF8qX8JUZ7LOuCioPaWOMB+eG399h0Si+Kg3S
YRAOt2yqpice8AvNsPNYmfoglMQICo5pOknaIAj6iKvxU0cn1p0T812WAFZsCOXq/OxfWhmWbxWP
pTUEWyVot0Qap1sf8lGdj4mp92XVh84pta6diQmAWXqEBCjkrP72GeZgyMMMot7n3jewThYculNq
6IUnILl37CkyQnFaUotMgRLigB5Bv+xO7Z00eOg92NRnoSYh7bQFDpSJ2dcpmQUhqTSqtFwEjibO
XvSMDHfwzEQT9Mgt46p33swdnhLt40Aghy3TZAcHcekAGCoh4Hy1wBlgF9lMtSRwPwxQ2d4GcOtB
p5bbLVPTmXcH9ympJXMpU96YE7gpPjiTUUtj8LRA923SOb2jnf9+I3ENeTFAhp+P53UOMafcrlgn
HVcrddBaTdZCi5+iDxIZjNwl1Ea7zDFi+K/h8UZZUZ6CJ+qaM48B2AtMHNU9TBwUNEh2NGMPAS7i
R9SEQ3RYX6XRG6sbHRN0Wrh4nhzu0Bq+jbUcSK0XNEBdWDSXL4Y/kjLnN+X/icWmiv+PCnHjKGRs
MWRmJnyi4/EAAK2vty4DLotZ+9dO2Apih6NhyqW541jc48eBf+W9M0rp4F8SKIic/TJY9SUvwfi1
s6qNYnP0uz1AWzmTG9+k+BxdBwlohu3sKlFscFiCZZ/pQGwaIoUp2+MRD3p0iLlu5UJWk3VqLac5
NKiSJ8ZeKISbIuxTE0biFAuXVp9mig7IJf0pLcsqCgt7rpxM0JhHeflLrX4873Wm4alUsMBHRtl7
GrUQum0y70rswCt8FcSxgFxvI5v1R5f4PCK6K7SptmWcNg1nenZRihc5l9ElMqwzM5tzDNX9bSlL
k6aWuaABCY1nM6T2HQE1Te5H9HKqq7piZrcBZEuhwi1ivrzEqiJMK+PwaVOeobL88x3Y+vkw8DE8
H2AUzQ35pX2HLkklBxZ3XC3cZv2gCSRG0+YJGxjl9eDr4K1wf/BEsQymxsixbt8F4VrM3wvLGH7z
sbwzLcnOZ1GDT4Nmad2eVvlk7ZIl99ds7Vl1WwAYzqbWtQqisfmzcd5ThDlmB8sumEm3hKlqa+bm
DEUIyYxGmzPr61v0S5I+6R1nNfVEa/gAFIKLH4H4ev2LcIKdmfACJcCQIXuH7ZKjsVMyzzNX9xCU
8vdBrIEMITI4hb3kL8GrrcE/ILX1pgpm2dBIAr1mffozdwovTMdcJ7W4E4bJ7A6hrKaVl+ANpWbc
4pEawrLcUbtSi+McuRrQXD2hMpnMosr/9b0nDrmap8q8+KzmMfV95BgPv14lf7VFtYIO1VkKUhDj
ZqJPHXruwUlxT2fzlv7LLI9F9Ql1micgr1oyPUAMAiO3gSScDjgPcl2dCcQj3GQCDtz+QS/amXmz
d/+rCr34PH4Re7a7bgYFYiZgB6W7QX/L3rUeS572x4L0EArxeUeXMzElQtqmSehxBscPSk7JgZMI
Da5WgZ7pSUq72tl5Vrn/MfgLf1dvRWD16h2gcUFZ7jYP7eJh3jeCyXXTVlq9qJHqQRBhPPpK02KH
iF27fPQbeDC63n9AEhq5ZcAlao6JJOSy2jTsW5YuIYFT+HyBWqvpBtk2k2qFpRZ6T8JA7x/4cL5P
/x+jaurO95SUTaCvNy3H6vd9ISRHkFNu9lAmfn2xq/IbaZerVRYiIEhY4+RBkJxPZb6G62Co4plh
O/G539dliJYV4W75ZQE3WoQaXRtV5Cmo2qmcZIWWFZ78k+Wa/YF01TBLcsTTWnd7jvPI9k9PVq7U
9nqq5H3SYjTO63R8KQd8VsKau5bVvdarS7PCItsEwISF04SEYsUWdMPTppxKC5pbkXmvKDn2lSql
elwnf8XU2Tv9tYeo9WL3U7wPRMTtN1HoLkVr/45OH8aoSgNA2IeGeTitFLV4klVlDW7jWZACBChP
MMFyaYWIHYo23jbxPNr8iV0c1XwzC1NqrZAiJ/0ZxvrX41bX90qqFK9nJI8wrMkF7NtsvsmCosZI
r2a/p1oI2LQ6xwinRTxH8iy57AyEcrJ4HIBg8ESbrTbvrP5fxEWkjKrlhG5ncKgASuYGHn81GNL3
W26XYgSpT8C81wyRG0CSIBx9yOKQvr3leenHtfJDKEbXCZUhOvLEz+4q5OzQ6OGRqiR/0M6KEYAc
EQEmInPQcV+8mdnw/zc3uh9/AcStrqTnhrzTsOOs04NLQW6oJeHsHAjCrnAsy8qm8iad96Z94W0W
xkTS0NDvSr2pDnRP9/tJ7bXowXXcoCPi7YdhySk40vkT7mR0kbga+pUaRyyxEobGeJAgOhYkPR+v
Q1gpVYj2HGLDcWHAvIjQKbzG5UqHp/ualbkGt3GZxX3S0G0CRu0+amkHqSpLiwQezKYBuiDDfV3o
xsQfdUd08SQ8XXwrFFL83mslwHiQCLqTuHhjeRsvwbBqCxrv0B+6rS4BLR8ZhNnvoSNdu2xCU8JJ
uoeflEx8VFM6fD/ODL1JEWB5yao3x/Nit3ttAk6f3h20bAtDaNbBdnYBQO0NKq2cduMEGD4hHAWP
9BSFEBHiMGZaRoJTuL1VoZ8C4StkN/dPvp0q6IHinhm1kxI1auMk/vlfAQkT35OMeFFEf1rOfyXQ
+1ah6w0PRhDmeDUyLPjZy4MsJTN4/dZ3I2gDqAfcgjy4CM9rz/l90z3GKOhNyFPmCpeZ+SfJffHo
2mNTNQWiquOxn+428CuVAD6EcLDsri3Xmf6ZDaR53nOT9MBlp2nQ4thh3vrSaxRCesZTDeAFCcB3
CjXcBmgvrc5J4S2saMng1EhNIAF4te1EYjdz10Lg6PfVF7NskLIyX914x+hKCmCl3mvMyWq9IQB4
B53yf0uJFi/bUsItNl0G9Osp/rgMN3K8UcikeiW1dNWwOb9TnWwNjrm1H8PIWcDlibExeNjtHlA2
BIwIJiBw+qnC0a3//JWWD3tz3xwuMN0jqwyUOcZEDRgZWmQLIsPyLILei+wdLhCS9/d7ueDazpRn
bGyOV5ZrMc5pm/3d1JCdO9EcwvUAkYDjBPmQCtx1Of5rdlqWwqpEV5Ux35D9woonbb7HQUTtlhNN
r3g/3KIc5bZmzknvsNAewgLApa4qK/5t46UKlfny3FGUOX+uoiX/HYBB7ONriKprN6j2030DdB2b
039rpgmg2IxJMiwX+rntsK1dVq+oF0pm+O0IaAmMgikzwH3JxKLdAKare65hEA69K+vs+btBaI4h
Bugxypml17gcb4EZnvTkbOCUVFOq1XN2HcKKOToJ+hpxL81bufmn2s2FmprAYN4sLEkxuNhxsaIv
VFKMc8tK1Pxm7I+aaJGGnaADaqOUbihwbYWMlzLCPxS0l0UMgV7RFbxxTkc/KEb0iwacFXIRedi3
sicPRYxAysg8J4xyFAedAiaB9yN6IHQxeZrrF9jhezjZKWee7KuVhA8uxXk3/UI1VNfrzuBN1TJI
U0Zq/pn+5H3JkU1lemlBjbpGmpqm+ajN6ivM/ushhCbJH7llPVvO02vhPsYgquyTegQONlAsXmkc
kiPN9Q+0c9BWLlNd9ec7BATNTMvjob+e/PKBl2ur9tldbmHzAW1/7e9N/yDXWOjy05ReIB4DK3uZ
QvN5eFADQNGsrMxhTWWsv4NcYLIJzhqEmVkFBs6IwAY9YTbu45ETfZxDCJE4A8rDdceze98K9uvF
rVLlBj+pZaHC4Gh97k/JWx0QP6nr3gOHUuJEJwb/H5JJeuCG5OfTaFLe8gPPGb3N+PePQ0hX6dAK
viwOHdH75wRhHe68t6jSpbCcWe0CCbzOLUETMtkV/zQ+8Hx9y4ZgmWMuAm+a5CkA4796FpFQHgfo
2S+p6KY0mULU63doAB2VTkudR8KgcR2+5lSHg772UGPpi53z+UVyKZ15FzTv4ucAQZRofPlSQ4Xj
hVMhgVGz5KNpPXxBwFr/wJM0Cm5ItE/NKyGr6r/B6lNMwahbZeafvLBjcTQzqohD6jHSKLO1x4kN
M0lzkWO4z1YwSdE+wCKQoYhTTt8CD0793+3lW+HWxeZ7a9tm6/9OGFhGAV94HowNQvmfUL3QjESK
SuUhskM4DUQRA0t86z5lMVNWpfKv7BiTpd31ModqMV3mvcxWK6Kw77OcLNY7sVaDlPinEJY+A9FT
SWdNzgH54Vk3g0terooxYGNfbV2j0lONA7V0REkiMvXGsKZWibtW3zABwin9LbdszPF12fVvpu9K
cKuHYXCTst/9aJ8Vvzhi7aocmVfZMDHCSCB3iXFDuaE0DIqCxjT4058/4kxz+1HA9gduHLTPDYaP
7QXIbvdiVO0le7wh8XR14liDemLdoZq5GWdxb5NQhhUgJpnrSjUNsP+tinu//JhiW/eqyJuKBCTs
NYHV3Uh0V+xCtwDy1xn/mSTzx+txpFvySikAxXqknx6X4OcG/bdXE/lvzbpBtAdL3bKAQpSpJ0Sw
3jncuchCd+yStVGWd3PKae9c3scPCLQCURdYhqXZmrPTOG7sQiryBJQ0aRbAlniB1qAxAEA1jA46
KWuVA3hB0n+9XJf/3gGTXIG/7qbExVNvL9ICoVihn9jZvKykV0aQbjGqkk6Jpm2WzKop6IJkidEN
lsmX3aPM+QXf25K+mXr8KySNR/RasFstFtTOL2qwDKsXKoIoAv5hP4G/mSEZSYTOv697i4us70jk
OYNIOrmCmOcyZNXUmFPAJMC96BW6MN1YgN9ITmkv8YG6ioxbQmUnkirLsWXBc5lNJxtGB8184tOs
tjCQK2/RmcRAnoxdqOPl5vXEUzGOFovYWQ/RqcRhWm2wGksH4CFndMz9HdwzTBCZF2mntcZ2g5PD
b/QaxaveNzmvkBFVMXS+SJbbopaqFydi46mMQqCsnK8K3rzZ+hM9nZOKEbpKtaE4QfNiM8XGTxln
T75BqeONXTe24agAMNMDwwJe8U6Vgf7ez2w7hDyQG6+4i82ikzTVnHrGaTodjPxzbTWMMLNrvCW1
G7V3fLI9CdLup2D/suIoby1/RJE2ZnkykRR5LFO5k+bqMdL3dOXUi773BdrqsqDT9XT0GqQIdhL7
7Gw5au7iYDiKfyP50a3Q0ZSdAhY4aN/sDlHTgzalu/TtSkSFvLidEbJevx+sWSTJ8R/y0+txwuV1
lpHnnYr48uMlJsXdLUD+jjM3XnBY4wp1JkknH3hvJRVhHnVl0MYR4MK6jBQcmzjbWkd+Arvsi21T
Hj0v7PqfPLCtZhUfO1gNNcQaAH6by21veqbt3XpALp8z1pP0ptCOq/PfW0fFSkJBjAkX9YpQkPQd
TGmxmUEpnuI3C7cEZhseMjWvB23pfazIa0a3izaObyn8eYfAn/VsB/IwMadtr38I63BxXYna7vk7
TzVZfODNe8TV8OnfEgENPqhk/JKKagXjJ16g/6PKAghXe7eSdV7+Z0AYLHEBK3BRP5Mfy/TGh+rJ
UWbCqxtFzpbnxB2WH2h72S8hGn9e7Hsqlr/N+mMERraBTouTm9y6Vy9vMWXia4aRsxPj8Gye+2aM
s/jsWeEcm9X+oLzC12NM8t9XV1ma4SRpQhO15BFNw0lPNeN0uMIerTzetIOnbqLf6GNqKLmCDv3G
ArdMr1HL/QeoUp1F6vkJZ2uc6OGk/imVf0LUWgGm3b49F4uIi0aSzYq5bgp5IfnGUpyPM9TymKZt
YNU+VINGU7ychyuBSSBTi9ddSbAC1MNQo5MoVYzY3sPc/xwAhtwAAADOZpGnomYbTbGGY6gD/VIG
v0fSqk5bZEYOCkuJbv91uVXNCVqIiMSyLFpWAofhdIt9MicR9ZkgfSgo+GQ5NotSh/Ujy1EqAJYs
2GR1G+rp156yv++1KDvBV5Ljw46eiVRrrDV4D06lBIVh6un3iZtWWtazI6RQB1GebuNV7QFvURiS
ek3BKL0fbqeLh3epfuCkiiBDX54oGAHAY9HS/SKHYC5dYJEBQzBU+bopKQZqauln8+3YZdc8eaBN
KGDh4kcvTR4PY7GAoDAYddN5AhS1/Nj8qOdwwCkWICUf/Ip6BjJZrUxTRi2kcOAfotpDPBTQdkVU
oBmuRiIFfgXEQ1q684hp9659Gx8XUzFIDXC7MPwpIi4qcz6cInlyGvYqE420PHIvLR57j+1/0cV0
R9FzsHNtD4mOmsa34Y78jK3/qbkmotCX4aypii4xhJn2E6gHy+S2LdcAh5oD5VYP0D3eg4+qcF8x
yy5Oqq5LjydVavnHCR9pmmBzfzuT4FQHGEqiIDRueEQDzmhprL6R9/dX+FxfUI3mwBTlSK7MSW3R
WUZuBzOKvbUO78wpyR5pYFvYJF8WxynWdqVOgw+/Ndi68q/zMfziHEWJgal1L6cVnCjl7AauuFmL
pLjn/ZswHd9VLlcmq892z4BMEh1eeev5j1E7xN+lb8hFShn96eHJn1cbdQh48QSTp6qUYsSnpt1S
bNeTURGBwT8v+mncpZHkjWUFSoFxmeAf0taqSrRtbQirAlqXaMZQvqrxSoV5BRIBkHiC5kJGCFnK
REqgvRIlOGMrhKwJyQlZWAV71U4CyPEdBl15pAjBhhqBcp2ex57UfDhVAdCI2/CAs0L2jLe5Dc9V
ZmI0S/FPYvYbyrXsoIDoPWV945BzU1qCt7mvt0QSJ0iJ/Ippcl7VPyBMi013oHqasPh8S+jFnDdy
70+yiGsFrCDxknRAnJPYZXaQilVhPw1klcEHkvnkghUyfMgtxjxVo/sMoaADu8cfBkekps3gihA9
aDTOoYobRii+dqXtABEMssAc7JJdef5HqRdvBhkbw/He643u5Ntpz/JhTV9PDvMKJ95EZfHKAgdS
jdzEwFyozf4s8jeOsnBEXWxW5dHQPgmSiLouI+V0l5ve6sLfmHELwxuysdS3ieEqZ3m+6LdqZq2k
x2HCorPZef9R/HcoLme64qz3qgfFSvzQ9tYwjl5rrGHSRP3TPYq4fhAWzxQxyMYj5FOYaDTEJRqR
z25newMhch/1F6iHFferzO4K16r1TNaUa42YVdIuoIdoWeDYIPumPkGAgDghyUFRMSJGZNY/7N4u
xOj1p1CyKfUbywZOOQ5fAJy/BpoaaS0d/59YNngoZiFsUjG9sb8g/7QoIjjjK+79nNZW67sBZ/1X
7nvjx4UJprLaOPLpGHUfpo8vtGPwg9vDLUUSRMnknpEhJqN25m7SKgvPGfScmGXX99m+589iCFYd
fxQs5ePwfPGgQy5djgyrUzIbztWA5MCSFjsHuINlBqOEd28ggZCtjzvaVF4hjQwaXYrv0mA0JT1y
Rxwo48x9xo1c/SJR9hMECPD1H+oOTmWEG7uProzte1RyAEccj4/Lp9OJboCD/ex7ZQ1rk+dUTuOI
eZ3Mc0Q5IiKNArdLt/Zc1A7ivM5TOvLthBSGhYLqhgRJbJdxYu7UgoI2FaZRpvAkXg3aGIBKCmph
VuzggUKJHT1MGTFkJsj4zIviBbMogbuRbvgGM2QAx/63QyMh0xwHG035DhLluJTvP4a5K+lSeE3S
/xgK+iOiBCy5gIF2v26n5jTec0y1sXWPHsmX37Pp8WlsCugUQePqqa/i2GyCMA62c00lqLbvN7Gi
j+o1muH2EfAPGkVhPa/nIKBE/wX95079785aXzDu5Qas2HaTgM9w4XOPCQkdmdCkQniMM5USH1xU
vIL/Vr/shlOvaPdktAlQBXcvfNw3XPoIRH8iFjLQJdwn6TxzlZww3QKSOWhoS7RRraKWxF79JplN
KH+uFLirh2Py7u2RwDVgdd2bDe5kYROFV0leqUftI9W4KDPCbqDOmO0dlYKdRu9/W7NjCc+M9+zM
YCjFTUhfFRoiMoNpEiBSp95k1N/qOIVd2JjFuO8GKa4PVkc5Ke5NE6Cxr2/8fqc5zWLrDejUhcTD
uahIDNgS4h/kSHQNaaemYaKKjPI28jBbdd4bh80LAIHAOV3ogZx3td31yjFHmbwbmziDDYjhF/iE
zcBCu3zZA0V4Xjk11IL4ZKM+Egpik8uq8LF3QecnUUI7Bib4+jJGH4XVHlklpVyaiUK/8x08ePoy
bY2qAp3N5E6Rt+5QBymbNOAlcxFgwkm2zGcZ9Ffv0Kr8+evmleO2hw9jaFsdpgd9UobdrlCOCGFs
7on+tBNMjOzrNMQUTeHmg36364I443UVzpLvvrFTs5UN0mI3b1G/GoXQUN3S1G9YhPN6rZy4xId4
diJ03sQFEJz0SZ1L1ieMtGf3MfrmfNcwzjuk1WWJHRzA9BDMT/avcWSTsRytODwukMIrtrwW2xmi
DKaGEJ9oyGOpedoCOpgoOfgsUu5f37FVgGRpcgwA1Pp+Tp1Bwu9CBdSqumwtfrWg/jf3aEjoCFbO
oMKFofA5pynDALTnJO9D6d1S9E7CmWvrk/3xfQOCMNQ3oRKNJAwRl3ACT7Nf4CR7frA9GnWt+5xj
te8lBivEJU/Hkv1MaNr6Q+5XrwqADUcfW19GHorm2wKM9I2eCdbsT2XJ/u9KN/2PSdSZ+VCa/r0V
z+YOzYf3/7nBgBflrosGrkJ3THzoXeqaM0l1UCaaDSBh1TM+fjII/wkuNPkOA+mMlxd02FBu3vZj
HYBRk1J/uAd+nk6VO4R2fN3ApB9LQcQC1j5AuiFfCr9RgR3MM3tQdvloU23qwdbYfU5RHtpONgUU
pVd5LOd8xMwZe64UmwkcbGqQiaNxnr/ytGDNjY3SAMZenpiK0RkIbYoGkOCkpfjbfQvKyyeDv5Rd
tTSwl/Bb29FtVBay+x5vBruHCkkOu0lK0SyXEHlxGH9rmlu7Mw8Cagdn6IEW2eUv8PjnC187erKX
l7hi6BLvdImQcyaIdjVq0e2nDCpV6ISlibTSd7SDTPA7dWzpRkVtrSQaOBPnmG17/S1W+u306GlF
z9kPlcPxeweWkhjaVXjT/zmEWDZmRxLvCrxPKE8RzGhVHTei1CTQqCDer6zCOcAriw/FSAW2h7/z
kn6JMTlzP+IcyS+NaFeRtd8/haF34+mcWS/UMiLc0s7xG4m/TOTjZjF/GFph1RZ3R1A2SfXNZBTc
ANRYElalQs1bzm3lTr5HzZI0ga1B398kxcWjj+0Ymv+iVY68tw8Vj873fmf4hcqES2o+BVnyFYAk
fksSLJOQsrahYb72bTMr41GsJdrBAxEQiTY2GmtQfJkUVk8zauD4Rio1oW/JHkAmSACbkCiYDMFS
kPUqHmQMN2SZBev6xAqheBc5QOdEcVx3Ldu2whrjxTwwXE9Bo6hZrx3f6XeyXt94TZl9BC2KoSTM
1olH9Za7dwolijFsdntT+SID1D3Yc9LFJ4/D/8YWsaaLeEgjyHjOFqEapGyruRo2uT4+BR4Rutg8
hqIlG94dXkuvqGvH9D62vUtBLof99+zO6Ba5sCI+5HYgUgJoV1yyL7Ae58V/T8PHJGHUVWIi9JZv
bBPoG9XXvsaCtkQkWAagb635sy+hLoFXEMs83CecQ4zJHJf4hPSjm+I8HMGGLIYrwbIEktNubI66
nA2RFjESiljeA4SC+kE+ud7JkExF4VVJiy2e6O4ug3QAVS59dQELBfcWV1LcFtcNh8Q2eqwJfkBZ
MXcUsW/zHKeq/DW+3H8ZRbK7rA9jCXLKvj273KNSiZLnfL5Q9v2aGHzf6QoXWzfyESyu9/RNPibI
J03yfKUk+GuZ35IOODTa03x1i0juIdIWH7n1IHe3xsAViw8FuZUL+dnZIjXPasIRytYHQDjt7gjd
QRtxQ5QKqSvSRM02Q7t026UmAt1zraNfpv+czYp4IMoCggCKzItb37ybGEQQ2oaK84GnUq9oPIBi
7Z8YA3Ul8eZ4gGLjhbAP4biTorM1PqzJ7Pnc75uunOIWt/oKLzLO92+zUHCmoeLIPQZEI1JDjr6s
MOdGLWU+SDV2MZYV9NnmemN1uhj/SKfoeFnSpOTdSiXFkZ75cBYFmyJBtzXLWjUnPYOmqvPG5GRh
HMkL9nvInPQvtuPBd/tZZeAlYmItQPoei8W3+cWdoRD5k0qePKgXjt1g5CmCZ8/DwYLfvjkxxB9u
bcCaNTaSo+WXWg3Vnvojw2ppVNW5w8A3N9WGm2Oc2kYAdO+mu3+VEQidOL8V3JWJHKL2Em4U1l5A
924isJt+h5yv7719NpBEP+a8WPaRk8JPp2dYM+sCn1bjS0h3vaUQvsKDvoXhgsF7Ez859QWWH83k
au/if/Opk4hyS0j+h/hlp+ZqpU5tNSQO/2UADvqhQaj/iqrDLdZ6WCRXhHdNGQDCG+WEipoolDlJ
0djZInCszBRfrBTX99c28XC6z7BfFwxkz1KFR9PHofsX6/RmpFavSUNTSfvd6m3yj61f2LO5JIJa
EeuzTOOBFTP3laLjC/Nt6UzamHnKme44p7mmqnNKCLA43ybZCQrkV6lpBvBTNv972OZyyQ5kPTAB
q/BAe3iIPvmbwIM6X2ijUbjcif6oaAzTaKbRxHa+m/x86Sp5n8/UD7mHJOnOZu/PMxKnY8M1bEJH
ySjmJKryRBY0KrzbDnVkwFr8L0WmFZs0ErvSHp9f1AnEpEPlp3J2AD/G/FltJZYQUB3CP+y+gHbd
zVVtL+kxb8kdhL1C0be5NtIz9MFWMiijFvsxR1SZWwQlQJ36YIL0JAjfVq4S1VFXC3zzHp4lC8x1
g3nfX1O7tTSmZKcwAZyNnCrBsKbIo0fShCyUg17sQDKpbiN03zZZZbvD5J0MPvo0moyLZvIcFtSG
qiZiMv1lsKmmkq6XvBBtxQi9iOK5TWurH3Egtax9xd7zSrxxkrTIHKQRD7BWmH0S3KibOBN1B+G6
bSaQzx3AVyEB+fu/ShFSEYQB7xG8EhQQcg7DWoHfJvJhoYC4YKIzoE1M3Q0n4SrijTT/GNKy6SfO
ssEMjbjv75avxejFg3YRvIjrXSTrge6LNXd28Io4uIhJN9PoP2mcs9s9ivlD0O7SwnhXhRkBIpyv
LHewrXaEZXOkNA9A+JRIa9Y9dJMBxZ9qhhGh2XXLh7168hK+6rbLJ/xK5wy5b1OtRhKw5tghmzY9
8jvu50d8/j8CSbYuPDBNUQKamEXyfzzPk5+qtty7YtQ7aEFsHBzFk7ygoF5U4fCBFWA6e3XF4ZSY
ee7BjOpY19RFBraJdsBIcNQRNvPtiLuWzs4xPBJfRtj1OpJnO8u9j6BhNcyRPl4TGwzLTidV+c9u
assBQxjTQKTNqAaABcHZbcrfkHN+D9h6KS3VywsToMzyHW7P6eD+C5wUR1SAvQxOcmQoEhmmY+B/
1KkisAjJz7wYNT0ENjJrXOkxqcKxval7aJN7tvRzf4JMTRUMVvvy6E55X6D3shljmVHrtj0WeZju
73i1UPtVaeMZU6d1YPjCINHzoCfJ/ocM1oMqX3ruJEf7SmfFzOXoFFBbuFaLJPvv9+yf3/Ci/TYd
Y1VhQE6AXJTCo1+LLRj9XUkqifV+ZbMwfE0/soiAagnT4UyrBibKriI8FT9tPUZwzcS4ghebcurY
kAxcW6lLVgSm6NcTY2WiPHGjJB2VnIh6JZlP5ZdDH7s2oRr8XCO2/TC/TZO53tgmOPFW49Ei+zda
ok/xJVTerokqonspKumCRr5aTg0YbzThbnGgGv6Xif4EdO8Nfs0P6PVq3b/yV5IJDQlAhgNpJ96U
FhfmVVsXES8BPAJTofrWcOKACArzAd1F+sSVi54WR1G2ZCKB1qcVct96rGbJgnlFS0gOgjwMlO5X
DKCRnPIvi6yQt0UjdG3UdXYr9ZoWANJogtaNI35LIXzmuyIdxqM7dMaqz9qWR1Z7Rxly3OV8xNHw
4iv3EgEqgpjrOxPlmBYZe+UL/oCUy0il3yHjSG5mfG4YAjf1aRn53KKhdzDexff1TuZsqIy5YBni
gC+TDDfCOcH06A2d9YtnPr6XUdQGRte4TF9wV2S931Wl+xbszQf+1dnJU63R/z1Xi3zVuHUP5BN8
dTz35Sl7rTEGuX0Gee8rxwDOPY2tdY1sCxyrdx9neEZ2m4PYz+SyeBHVHdKrJmlJcMm+G7/omMhK
6BotttHwh1rfK4moArml51X3qOJ6zdsudNl4uXForC6sr8ocjyoeKj/TVNVN8ViyYGCBYRw08+cb
yte1O4q5qTmm+e1Ml0155BmEwSiu1pHQendJKQ9U9m4r0klAcf869rEb/WvE7qAfPdRq/lzq2SL4
JNYY6+QanuH4DPibkDBShloASz0e3KLXow+k2fBX4awyTOlneD6m1Xpuqb+eUIYo9D675WUyoy5k
Hab6MNlHox3TPrnHr5W8RFCArecN/NdsBkAzvZyaShAHaArLzntTTd76u/wwwy2/5ysWJv3RBgEj
JrGk9BifMN+qu2/EqyqQkAYH3123rh2mXoYKtLovM/myI5NMJxWtZjE8gKqiaZ2HuaDqYTaMe+22
YZ6Z/2KKdn07p+Klf3azxmDUAyZJVoff3lTgutgLvC4PCHL5WhNmIKDWfrvkVHieldx4DPYI8BRx
wNtGhnM+ihuNizco5FaHPmfctdWoryaBEhhBv3ynZBf9s+M5aWuQ99wVT8VJTlL/keKaKyKA1NmT
HeAxF9I9vyA6w8VcwWf43O6QKrlLOEtpHa/bkJZsR+MiK/V39hTq0it9pf3U2dotAy8gex85n1pn
JoCwK29FfcQCjv/hFT2sac/qxGKykuRFz9jA3eeIwPDphgclq0GtGWX88jAIHpaPZLzU0MLJge57
otxy7K+dkNSrcz26bRy8n/zLr1Gr46/7El65wSc5xJIKUP+6CYyvCL5z91wlA6iJ5ca4qRGImTwm
coBSMNDvD03m3TyBxXdRI46D8i83lnR9MFEXHJJNvZtfQsxRyb9winjsSg/PUjb1y+G5TWkez/ks
bhqg74c4OgxY57UwTDchySkC1Kafc5OjF3HEPE8mIhCEy7338aZWsgBuQeTDcvyWV7Ahe7L/XFJK
jK6vRBBl4+1VETa4JWYTLWCNQtqtpMBBl5RJ1olFglHzTYShfgzIX55/OKWnSW3+RURXHTdY3aEM
XY19eKrtfgLPzIG0Sn9krNE/AI39A+BJg+hK1ZA6vyDNmQ1tJ0BqIZY3bKmwc5P3JV7WuB9GvIW/
WC17FNOEflnwCazGPgjc9OUAlI8H7UEmACzNsW51MV4u7pk1bET88KtGrjW4YDkd6/xjJKlAH7u8
YhpXBFT/phbiT6LRsdxtmIKVtpmfyylkyzuHXwz9UaW0AFOI1bMc2rIZBKYjjRZRbDEWowIf4nDQ
LBPRhWxXJanqGRyYBB0qc52MlFOi7UPv0BM3STpErHy0a50gHiLW7d4iXBhFMVz4A8xzAXOa5qIK
iJ2ZfTMnWlLODgnVZ1WSR3z7Gec2KV7FEeqNeAhxaFlM9Bf/6HHbplBNZSBLgIDnHl3H7g1U7WXR
Qow+Fz00P9HyfKRybSxxHaNaAw7ovvRKztS9JMuXKYmFDWN33/0o88j1nb+i3i5hR82zCeiRblEK
/DemH31WBTUAB+EvVUMp3QBAo23J+OMZVV4cuwjvQ3/HqAjORmXFMRC8/ETMscj8PJmcOeWFDBko
bkHw5SQHALGmr74wkEuzrkTs9NgPup74Ed/NHOh+Z5HIJykE6xh4bNSyTr7QLUTahCYv1sSNmKTc
M6OAmPSPAvzgi9L1LhCsC+g3lW3dgXsY+zoH1pprqcNUNeXKFO3x1v9WYs3WrZITQE+jLt+8ZdYm
JkuIW6JB9e278FuxeTMWoBruJrK1TJEyItew4cyrYdAejRU1zpuDzaCJlFTmW0QhVxeh4R/y6t/x
8te/vPrRw27KOv2JKnrg+rFncYqI1b9x/R/s0avIeu4/VBnq7g3KIUq1EdEbwz++lWMfXj6MH3ny
fUMylR1O3Y0wPfkLg4eR8YmiBsjzmliY0ps3neAva1c3SPahP0h+XLb3JkdFcP7oK27j+cndNR17
yrc26gXapDp54RDQ7Hn269twrOiMfOzhVE9PfFBDVI7TZjl1mavmJe5nwyVlZNKsDahFF8Jltkkj
UNaa+8aDq/wt/DnzBp3i1PgXr6+JX1VIATlgItJexOe8g30I6CvfYWJeNWxtSsMlHZE0ZLDcxwJk
GTdLtJJokz4D/NfiKJzn4Tuf9NZqMEOfe6FOijHwmDMJLFmvaMQAWtdD8T0N7MtnFcgyhqKZ/ITV
icZUSvUe1TfKAYFAbSC1x8LqSYeVVx2OrL0EbsZa/KSJGBftZBQZxjOJvdvNOFnXVskKXXdrjalR
wA7BvjMSn38ZG9CrbDi4tzufUi1pNwh2atRZn2qfZ8T/wOXJN8Oy3nJvPCiPIjCNPvjD2oI/tm41
fE3/Kr34qtpBx29+SyLSmg0w+Mxl8nCUx+qSWn+8SlY65oc24WXZqH2E9npt5EhTPnt5R6zMJbm6
24Z/m23SU5G+SM5EI68DwsdNPVkLoA+a+hu1q0WYSk7tOxK2wWyxU+hSn0UfY19QCVwOK2vVMj/N
JPe4+MatJlV3ClpuP+6PkJWihYfsxUIRwVvJnaIfHNcmsuIO6dNbyerK5FdbfNnZMx0wYKf68EmL
FujMyaLjSh/cILWoi9QJH8joKs29U5+485DbE2ITVog6wFmInaUAYsbi6rjyKesAexvVlhO4KHvY
vMTwVNd0ExzifjLrSoAIwtW/xwda9aXn7c/hZRltIUOqmGyggMwGmjk7gw0CXq9g+lFmtTKSrHIQ
OuzdA+FLs3uLc6+U3ANFiJTXeyfZeUZrQXOAm8lBqxYKPsuTtJDE+B5Y6tDZEWpH0at0QEGU83EX
wd7pnJ/Eds8sSgiKEAMxvmRBxXXSpnnrr6nYvKRH0rsVPILttUl2eyRw+lcsvzG2751kgrKHg017
2UeHDNr0LF5rZe9NGdqEq4ztqAAVg/hU5FoMukT2XkTi8C/4f+McfMAW2IZCXrFGEDZXXNay+0im
8xh3WIYyj9wLMsJ/lrr1FEcvZshgE8lyGNi2uf+TVvMYMobfUsWHrWS9nsrocOCrbSOJRAqW6kQI
u2M6bzdDGIEA/i4d/SJ5c53dIKAgWdtc0fA96L2PIPx2NFQuuC9lLuD19k0PQ8Qv943xqjib+BQs
8A8OTzQ24irTJhOeDv9vWDikogivJ7irSsJaMCY+lRh8A/j3TjjgJkag7CSsuWedY+zAkowEutMQ
vnexk+aRqX/y+9mjadg9/IIvMsiMmPZ1n/GyJeKKsCAHPCQxEDZjOGYg+n39MOPN7hxQa16drYRD
aiFx2BLujFm56dmawY7W8RJ0qrIYS44ScTx5uzaaBcEJZSkPSlTIEnYZFPNb7rRPE5HdesDDPFFc
rWgLDdsckkYkSe4JLLWsGQMSxovvf4L5RMeHfohcbWdOr+Vf+KglSW2ZiZdMR2y67JBFB7eYSlef
ncMfXxC++RlJ37fondzrlx7rtKrQ1xTh8I6/8xkLpbjo3iiwQL7ntjbmYR9P5fkaM29zj+3NDgpp
7w+LwyfxgVA3n27RgHzKf/Us8ytuYt8WRywAvmyiAush30Sn9KDSBfuMF9/qFAwm8JPSVTrQLgb2
+0yJSrYyeF/zYTu4/nfneSkHV5suy2wDduB2dy/PQzbzzrNq7oCfFYcuol3STTuj460JBpL78R10
wPz8i6ElkKI7nZ8e+ODQm13hz1FVmmH+/t3wVOB4oxnKwFZ9BJu5VXDAeQaOVqE9JR9cNZfVqyzQ
Rndl+WuUKgJ1YGf7EZGA4tdvrmNMXGO7+SvW+1rhci+sa/P9/H/3ch81EHcuI1RwTKMdjyRT4aXN
8U+Tgt/WKQxyz23YMr08MNv5Wdy0amndh7My/2b1LnRwXMssSo1qjEJ2lw1knbMy2NhhPNco1hFH
0w8lw+9zvYuYw3YviOUUHHLwxdpqlOANF0X/N7i3rfE21VsheMsKzwc9XSefG18q26rFRSGbUOu/
+PKXn++oDr/puFXXop9eqmfS3svUCXu64dc9VGvSwJETDpQ4lzv5G+AmpH/z7TudZe/fgQTtafWZ
wq1+g/3nmPYXtawR4V2J6ui+WIWaDrNqxFSKqihYo4AYUPDrtCOehR/JwTVHABGV11FoWZUNUve3
DVEHcEKXP4WZZpM2KDhEwI7tsTSf+xjKs/KNImTs4cre/HOaf2887Kid840DgRxotQEaugPDXSmc
YZ72JyRjjsJvVCK7RgDtja5pzRVHOS1olrp+4Ns5P4gIP51d5sPih1L/v/i1dePnJ/ZQxHnimYSI
inwjmqITg7pRRnfSSiyjkbg2stLwsU0BZQxwa/g0x8AcOasodw4Fu0/cqKXS6ePwVPVecsfay7yb
hMB3tZ1/BgHOhA3IgeAFZoLTmii2T5QQCOoqEqD7oJBrtd1b3eTQEXRIt4VvJMYz/42hNEmDSQ4x
e+HOGW7w15AbPzdh+IY5ajHf5uV0xW2t+WbmKJOSLVPxsWhSHlEA7XKRuI2bwi8sGj3wwN1NANPz
JLdpP0DyDeZj82ciACC1ucIQMQK4ByiaKIhmRIdQkok61Zw0ZOPBu2U1DaAQRFG929nJyIrg8M5t
wjNCEWVobxfQpJ0zNqPgGH2/d/2cpjayBdTadgjbsH4bOih2MAIt6f49W8mrqzxlPGa4ddHYvm51
YsZ6NRvdpXhSrHkLx57l4ZSrgOU62vapckceaCGHW5Qh/KmjETqE/lFKZ9DIm/d+3vYELtkj3XkX
Q/x8GjvOahVkHjTadDAfEM1IVhpOKtcLQ3FrzsJlFUiyqaqQul9uCIMAzE8NpicFct0glbwULPR6
m0jsKYgE9AyQtpEre9pakG0vOoxTCQVXzmObYUD5B3vh+TVUWh8nLJDO85pvNh18nhcVXCOo8JqU
+uuxrecwb8JPDT03xcbjw/WStm7iajsEakx20xJ/vj0frREh7VpANl6JLS8DE14B1JMEiwKHeUbM
o8vmVVi6oEZOWAse1fUuUJu+YQ0tC0ehSZgnCofT/BpwU45xJhUXh//R5H1onmsJ0gSNaCkZOaf9
lXPaJ2dDbHCSKvlDbK6yJTClldabIRjTlgiEJoB8YMMzWpxgEEguBSeR87KVC2wZP3Z+cZfgHggS
u2P+em+KN22apjCa0fVKtKb6TbsHNOBMqkbIL9/rsb2I4q1k3uG3bwFT9yHWN3+f1OeqdbfCYK5O
b/9GmAJyZHLl1HDBWYfTEeCol2zIpyeN0UFBeGl3fIy06d3pmftuarDfrnbHtq7J01dMsXG9T6i7
tWZuB4YJqWGloRfCKHdH9O2VcDO/8HMUDVDe+8X4zeRF14gjE1Y5KXgeeYBkDsPv1k8KKO5rpLPI
t4hr8mgJ4QTWfH+iRI+dHagP1DSBJmwSRtvO7HJZLjkYyfi8xPXM7AjgNOaMoAhBcv/qFBtdG0Fk
CgBeYgjZakcmMjB275C+McbFANFvLEKToCgWk6G23PriqFYbvFxRvMqPaSC1WA9Sql1zEco62Lm9
i06XmrJgV8L70PZpTFWNkDehRLMH5llRY4xXKOlc8VWdLR2npdb8WSPzWGlRq1/JfL6BX+ZCtwEj
YQsDpn4HJcvKRUbmaMLIhDqjZZT0uUJLtfng7za4a4GeB/o70I40t8zZPQppmlhwrZSa8yRV8Ifq
3p0dVSRb7Zaq+Sazi5iQoJXu33WBLGx8gnjE5OTC+U9xFdo5VuRXZ8PH6k5lCCzmSV5ABmiJC7RR
ndDI6ExM48uoNxCmXyqPPmEtiH4oB2z75HIdjMLBUMGbehl3nKfPpIWZTPIQoTXjh+LAI7PVHvNe
JfG3RLFOepghhYlD2t5SQ5+9H7r5/JaBKzqKdhrCr19pfPNFudNesyA7Wd+GlN3TrEnfTmaHRKVk
qAMKr396prwCYFRawSacf620+9k1N0r2TDfENOrg02kUiXN0AUCF8iJl0OPZIW+jwu0n8q9HRayv
AnsqniXYv0kLC1OfIzqS1hIqihMeLmH6K6WYa4X7xq/qrilhnnWWwh54vjhZgDQJh7aUyB6nWngx
Bfh5uXMVErFleYkbWyvirbjhYrXxY1vEh6oDgrAbzGPT9Q6XuKKq8z+slv+3X40xkNwDTjUj+g/X
qLCzKHCNRSUG0Jlqj3sleR52Mdh9cpAtp/Jy9aMNyTVyyniZdb5jZRg17FC/iEZmZbhXZpupvI9L
NTQKzWKSzI7J2LQWVORidz5UySqeWUvBkC6a+I3A9Bh1j2hN3rJ2fP3jF8MvrSjNKST1e4hI4Xtc
NFIrV9M+EraXHoYrcM/lX7uE9sebP2fwrRyqZm5IpFLSzsG98I66QhVr94zb4gqEC8GXL0IZ9KCh
wC0IkxVucl5J0t0kI7KqW7V4Ui6ZLnMd7uDLIz9dWhdi/X9lJFZv1MT94zGEjMHndAI4UfjcmvIb
vZ7Og7QG6bzcWhgWnpw1CbbTBzCXHW6CNE3/L4clT1a9WiU34jrk1X6l8+ABYs17urzxQVWOB7f+
1ZBboafBOwVQok4bQgZQ821ztuSdB2eoyrHyiZ0fzHmq1gHXmOOc/5ZmG3WBRSmUaDcIyofDayup
UwVAXB1rSxO2vDSKcWos/ivTLLVD7+pkHCjhlWi/Yq9/7XWZMpapVRYmevNTpsZVGGfbHv2xFR9b
Z9YX/tNcZJBUzMMozhs9++inV8iK+MwMe7XsWL7vuk+q2kUx87795u2PefSVe+Mi9ba8TQpDdYA+
4J9Gq2x3pTrav/dWvzpKw9FkCSnHDFEcjR5hpshUfk/NBcgiZRcWwLxL6J9Fs7WOFN/QvY1u1OI7
9cjniywAuPv3ah+7zazbkuKtq06EDP2xIWcZKdoNsduKumoJ8vvLTi1/xtHf0coSUxCacMaFPmDx
nFoBBv+FKe/QpkOHWnKxav/bj96h062qevzDSp6jsS5MxBaP55UFYz5oteILbzyVYxe3Q03TFn3A
fWq15fga6rpLpiX2cAmzWPc2fxRND19nTm4Yt9AR4MjhEF94coz+6ly5LEIA4rTB9HFSij8UZyFw
rXRvZzlstctXQrN+n30rtK80F/gX/GsR3bST8p5+6+qGbberus+hP0stP+bXRKvBZ9ecs2/sYYa2
Qy++1G8zO9PZV5QpGZ6QiJu/kuoEu96co/foQccVuPCtgJ5a/8iCVbEdcztYpTIHQlZxYV3aSDJN
oehxb7OlIIuGVCyyUn7EWiLhA/a4GQcHusqgsnJjKlYcIlnfsBWfSDP+2Zfzh6sDYFIaxeGGjKbx
sU/jyt4Fb8QLfC2zqBMaP0wlBB0SfLPUI9mGPpkr8zgxw68PztgWQ6hqD+GCVbWGYqs8tVfYx9ZL
g8mDo6CpVGuWKVieAfG/odoJueGhHy4485qiTVNQRJrZ5WMl+Qur8X42YKXDjDIJ77ZdiH0MO1GI
KysFRur0Di1B/Xfse+u79wKWbj+761Js4Z1vZrx0gqiLIMG07yUfjz/P1hayDmFe5NElqyy9qIc6
2JLCQ0yoqtWK6KcuBIIA9a2TpIti0GucPfy67PxGGBZiQONRfknZ9SZKGKyvM6G8bscC1lofqDH3
FsCL5A9JqaR145rMcE4u+9ZLBFu6mnDjPnG/OV5ugK8JgWwgRb7AbSPVXc//ulu0ZbJCeUmiez10
rrn9y3yZYqmX3GEWWvYA8wpYWIpPPE+gyu+0lay3C3+EjQqct1IZzPO6elDUaE4R/zmsbteKQUiB
hl9Qf78P0pH6lP7rxnRI6deJBwsK9CnwVnBsxeOm5cubb/zulAYCuCTm8WeiwnCee7rpfoqs6ADp
Q8asl6a8Dpsqkfa4EeNcpfc5HJDlJm7GJjaAww7n6a6/lJPm2UO+dYyAWjHmAC0y/uMTnyxhrpOF
dQTRn7VDmaMyBF6PYCL/lZse5VKVacg7feZwYpsthIhZSYXMcA6s3x+PX7MzKkX8Dkj3bKN57Uce
fPJkN3fONimBzFX+XNW6EYHA1wuQmZXHJ36Z/B+OzEBI8VJq9XEzY7l4kh0K0WxPmoeb5Dn3N6E/
NM1mfu1QruL67nBNApgnxyVnAWe3ib6AXMDWMO1KdTImiDwg6gxeXNI8ng/R3JYXV6Z/Pw1bLczq
GUh35uY7PMr3MwOQfHGPvgBSLawCtd5pNCPI74Kc9uW+vP46KueCO4nOAnhRtZzQy3g4cAkQSRDK
jDFqJlPmQP+4iezNFYPVpVZUi0E0CTRjqyLQQ2nZ0Xo8b+pVITq6REMOMgMQAhoOyvG+JY2VO5mK
3m58c8efcdN4fC4Fys2u/70ZmSsNoc+NZh+RB8JsmGJB5RZ9amjux+7vW0+d0ijgiJfYnjGJGmjn
1muy44EaKnfjbNzjNpgJNrkmxlHZmbzaVcQ4tCOO6nKRiHpTuLhkrCO8KPGi6rwTTG7lKTe85iYB
3qQq0VZNSfb1B6iR9FM+r/5XdaifB7r08sPAccTDE8MnpkGR1Z2WSP1zP0mVVJB6S2RhguUZJzmL
fmsPCOe84sIR8/SVbS95HS5lg13bLATyWiSmuuOkxDFaqQCkKOsJ3JVowuFh0lD9hZCZVTMxiwYE
sWCfpslKoqwurdXjwNVkbWASs0z6ehs7WKbGkHlJAY+vGYpduR6ymbSRnHk18iywbvmfYwKWvIYU
F+jyL6Gt0/jR7lZVBcQL3UWPpNCeiujLCJBv25HnzylhwDAqgu/U7Ap3fMkOAFM9K7fOySsBEBRv
U7KPNzOEw6VZIZzc/c33R1ftyD8iXwF7SO8DIEOU6NUsl8c+UdUY0kSYPbzqmap/CKvt1s9WoAZd
rUPe94Wz8xNs8lHzIz/oRKTBio+LpqNZnzrcOHdXRr9GetTif2oakot9sDbCWO/GZ48j7nwUGlpw
wUmkx0fzPuqVnDrQbxe/NiMC1j55PV/1sGVV6EmktYjiRhlCSDdm8lohBiDYza15BwvWgc0lSCfD
OCnTMS7d9oOyZK3j6oOUseFgI5ALKH+lDiqBdxvhRUQDWalU7yEYHd/SdH/G1h0//YrU9mrKmnip
/2zRP/Mr5PD3X10pcxXtYLbkS70Gt1bC0jr/OTyMyhw2Ub+DcCjMx3QV8pQKHIHdpAAwjd36KO+K
c7EA34v+9dN+3Lp7eD0k0bqt6Vqx1+vLz+IHQce8PDz0KHJyWzkTq4Rj83eFw+ZNTS47YgEheYEU
DOs2yfR9qAqVXqNLNBInBTllGMV5NdTU3uJssNf928gwFgrp+V2luGOw1AqUKzYEsBaQmE7PH23W
vZ/ARrrs/kMxQRni5lEFRFuG5UKcLFN4K8frX3brEME70DFOcmD4p5y4KSnSx9sRyDSq9R/WeTZq
gMVFEtueVeMIK3QxnBbCTNMAZu33PdMJuyIykw5e4eWGZWbFYPL4CcCCMr1I/eHY08mTmJaKmafX
c2b+xXIozKcdz29BPkuiV9lvu0F5F22ktMDo+b0kihPfpgFqIZ06ZA7Fex3kgF88XZkuWo2exmoS
H4Zj+gQgFta/u1r3LpfqJUV+a5553ipmvnIadwDMMdsy79sIav7W81tIn1HZp2u94cFPO08Cloh0
ghhm5TgkiSN6RHH1lWSbmyWAb3Y/nMtkr3i4VjrKiVljq1cl2aoY1tbe1NeG+KZjDo5MP6EqWCKy
B06e3FIL129uUvoqxHyrX48+iyjfjQpZQebSva0352rRVJVQViAAp+aa4JcXZrCD3CiyB/QQWXjY
jyJ+K7FXQinSIgazG1iKT1h7xS5xRAL15jLErTnFFLPPYfIr1wxJm7In7CvD0jPpx5raL/xpT7P2
6WSaQF+5Oou/t1J9qBfL2wkeONKMnQVNK8zyxFu2PvexMSdyiTC+XfMCtRkeMMbqNHfXvjwnwiI3
rkX2jQRbjr/m4Pngv4NRsbWWgkIOjFBtAcna3XSHxvfdXjO7jWx4NMITin5/as5zBx29zyTPxQ9t
3F7PGfyVI+JiThnTO3Bm64/Qwe3eCXWgtCwMjxKVFBHJdHR4UI6TytjyBfYRBSMXKHR6SAgCV9b+
4nHKFCB8ya2Hv0uMGvheBvJ4n2jPseLUW28m6iChP/f3aCx6pgo5EZnTF7RuS6JjabvICkvun2PT
LPSMTCgVGQ5Y2JCjX1dy1tdQtbp6H64ol41a2kNTlIvcIgmKheL/U69E7erhre+CREoqGcUWxMgM
sjOWXBEJ+IgQXnGgXHQvknOXYaeN2C9lCjei5nkbqk4F3U7956kIvVxZtCZ+Z7jzGH/UwRMng9OP
aJk+XIAUyPzMiNyI7us4rqumoCKiH2lGQHnwPLWvTs4IKxf/gnOMAGBbFZ4xYoX28JFuc9XZu16j
dHhLiWbOA4odiVOWIkgLDz8PDZkm80JIALHZ26e4LeEZ0X3m0sepO5Ln6zR1TOLdKUVIGTUOKEZ9
zBlpfJ3yV1+ix2NMovgf210ARmUj2qyw8tvXIKgHcMbw+V9xZGql431mIJB+MC5KzNhz/VWXJVkK
Si6ZTCTeopspWYbEl/i6yeyIZ8NPf/Cn4ZPt11IS+58W+QW7OqEgVgdVroNhjsfEvxP3/jPrmYR7
xVMQTq2zO5JTI3f9+YvRh/1rLNKTngGW6C29Xaap8eZw+K1YHCuoJjrTBbvTkABw1wSklFmMb0F1
fp432+MrrIz7LDzVlX8GBdfGVf9/kvVE8d1wiYZtI00KMRA9KdhObA9cwjEiwMYHpo5CLpZPHQLv
ySm5bkfXPXnI3lSKzX55prs2Kcb7J/ThJjQEiXEA0/DQcsltCuTVpF/0MmrhZr3Df2NAehyIcYaQ
SZP5bo8mNMsH2VF6LutD9lbiR3wAUyd9c5m+72/jR78zPkX/+EDTfS/fDGUbFEaojrcD3orn85Tb
z3FsMnBsveC96FMdizaS9aVy5yPOrkNMPHUOGKVsm5MIHYza61vGsZBlKq7e6KO2Ubv52pNCFNnt
GxtNsBZwtBujam8qVfR+ss1J1Z1bh0mqmBN0CVKxujOpqjgUajWplkH4sqvl5+V93UKnK1KlB5pT
VlQS5MYyj5lEjgi0CEIx44Zebz2FEtZO+an9hxFUpHrJL0ZurCWyOXUq2NZaIOCjO1UYsrXAIIyB
QYXlcOVUCAtgK40QOHko4WHO/BgGp3MZK3r2mj4GoR7bJxcvPStW5K5uPVSEEWeBV7a8/OqWVfxv
mljn7lWTIkuKiLOxDfgt88lR8id7jTerFRRt7TbtS12JL1uzu+9QjZ1iOTVgeF7jmEhFK6I3k3E/
DkGl1KnS4YSmvZO+NP7S0ZCJEr3XDStDdjDsSmTsQ8nIN9X0XlFMuZ3b0uuXmknFmBYoUIdHkuRW
b1t5EewILlKDlQHuOZ1a3y/P1Fr4oY0tTa/siImcgTxN/f78ImVjLoQUTBouV1fClb7i/lr3o00/
nGmdXA7OGImyf5qY9gAP3+Vunp+cOczqrOWM0j40bfjNyudXR0b5J8kJbyTMDWi5rkIFlUwHJLM3
mbBQ+8xy+WH4+A+OHRn4gBHOoEz4VLheWsoZEmFmDbqt1DemHBD2ZWDfBbisQP19ebmMkE99X1rG
mPamATTPTrCTdvONwMKeBnjvRlwfi72aHWAP+aL5kJRCsVr0iaGFacTe06GV3ZRANk9pZYvdFpDB
oCrylsaMEeAzQDdMn2Yh3aLXxaRCVlh3nI+Nw4Q7Mvi6ZBAAeJL5g2EF3sKWaL/M4AzjZAEdGJLE
GWqsCh2Q6XKvASf1Q5943Krg9dWMLUZoCaysGBOFOksDWjlvsl/zHUH+KXPvBHd/+PXe2XlHEj8O
dCtp4b51kyiknmTP2xf1AoBcZp8/6ehf3Po4MzSc1hTXe7YyTmrFV69jtMsNQhYMuDrB5VXwvNop
gHon0oWecBZq25W0aY4Pt5UYM7wquO5RrfESh2mVj7PJcBd5QdryRngjCYCFZ7mfyCuW4WX/GdYD
+N5S7cuCalEddS9/hm6CrNtiklx79Cao6QqprAjgkQZq4FYTcsYpUQxSl9XLA6bnPe3l7PPlXel/
PL9ZdVExWl1B7J2upAcNv0EX5wzyVjgefwWH29mha/qLb4/XHnVDBAtL/JbQkGwd3Gj8R92j2v05
yTUiE3DtAwqYxBZ7BUuEf31omo4Yzei5LxE8EWbt6m9jbeh2l3HSmynd3IOM20CVNTttqZQLu8E7
DWSDbmScBerFZTs+dhRxvoZ6J+MvaAezZK13RVgRjtt9RtfW5uwGz1CWXN4CZoN5b4jsMP0XnbEv
a2aapmn9HbhpYKfA/NircqRNHeyxg0QVClcKYX45CTqrUBqxzsbNhqMgAWmDPt2JUOKldwNONTaq
FgJwaoKwbp+EEME7wsBGeVKY8RZa4q2Xs0mhcNyMG/xt+12xpZ/5+aYp49a+X2dSH00su03Q0aIx
YWcNDbXBL+OvflBGJLGWSne/Kw4r7PDSf66Wkh+VrioFBGrNxF1iQ+vht1Elj++jO19bR6vwSXq0
byIat3wu+aj+O0DUMAV3RcPj7ZRpY/eh82Fnfu9pHCjVgNRUutpjLp93CrnqmAF85e1sO8eM9jcb
qhHrLCtIrGM7wU0X8u1dyVPk24o+QV4tZAQHqswrXykm/yWIy/+8eAXDhMcSZ9G2roOVbFs52mk9
a33MJX7hDJfdKrWyuJbDk0WUxui5/g3EQbQonRP6HGjxDXycom3xE1m+cPnqQ3qhCaHW7JbBSrwY
YlERmcz+mNglXm3Ib4kMu9az+F6xbRYbhjga0JMJDA80nGu6Rb6hJp1g5nZPU1WS/UnCctx55y03
F5yaagkrrNX2Rz1D5r/3uqU1KTTqhtFvsqW/KTN/GgyME8BSaptVPMnTc+kj81Eb/JDn+SCxu+71
C3+1aomBArBy97MsqUQDS6WD9vh1V2vRsC2BP1469hvv8mjWYtlY5Vi84FISzrKCXgX7I0/Q8Xx0
oZOtLX1jejMRsLGal9aHyxdpdCS9SMxISnY/yBQ27oQjgJuzl2vvqvbCVOvRyxJ918o7c5bdvqdR
Ft2ML/FrkD21cY5imBB9+ejI6+DLGxwBtzVEUvWvjyji8L0/9zX7eX0lUQ/NWDHJe+nXlO53OYL6
IT7ZCcki2uRbyaS2lOLI3PUKWuYW3bhT46liIz2n7yWWgeinn4hM1arkQuOoAL3JAhYwZlZj8A6+
CgiBcHpCxnp+iJWUR9+ij/RJ4XJhbfR9Two0vrZW2Q31vJ6849BXjsCDACMUda5eHbD5UG26aT7x
bGnqKtr6RrPXBaK5eDWxCRhZjJni8GtlAZLssQAz9MeEccWbqUrfMYhneEm/eSPyjvlMR1I3cJbS
rIVCEsAN2Up5x3Ea/Knxx6BKs+mHp2M2oL3OBJ1a7eGTo64BgQuyyFOX/dcy6xxE6J75lALAMGs0
U5+f+8GvVg3kcs9A6xszRpgskxzLyvKH2dx0t9yTAZvR8Rp4n7HvTjxDULjXyXTplSAd223KHCim
CVLF5BTYd/7Uz66Nk1+kdKvR49z7i/s42D2umEASMn74OayzFgVLPFXqKTEYobnJkaxCrz6Va519
dZYEgqMHH1ahIkXxJQgWQijJiC3/7WmZNg6No/7CSEaem6xIcGskthmicWvyFfaB66I6ibLf5Z3u
ENmx8wn+gOdTY9aPHPkw3kdxu1n1hkq1AEww4nqu4hpLOdFN5meu8WLZ0spC41LqEjzkv3bAcFAU
q7Q8hdmlAVUqWuZCcQWVd2brFZYfGO4wsVHcUDGiteuWWBlG21GD847DlogQIPliVbMv0XR/5Ml6
RBlIOurXrLJJNPckJCIw72Ov/PLI2TMnf9ZyyLJv8mPYsJt0R4Eeo2QKsW2n8yYmMFN3A7Qu/lhi
hNcHsmM981K9fvbOaBt6YS6A8dFizqmBQIUd0atYm02Y+MlgMZOx0jWPlhSpwGpPKi2pSDj/+ov+
BO2IDrywfnnLCxX+Ob/m6OglnzWmqYdcv1odS73pHpwWssNk/DSp4Bfg4YCnf7wKH+EUyQaau/IW
QdR3VBYwVz3LiBsr/owlwk/xwhymolqsjdCi5b5vT7cXBpDLvfoz09qSgc4s3Qt26tGPqOCpX+YE
6V6VigkJ/EQB9+izFU1Gy+VFDY6XnexK+9UH6yHApTtVkUNVsMm5ZxCg8K7u4ef9cubSKt7Ayh/g
jmx0WB6TIxP46X1F7/gSTZSOtG1HR2hLYTxNdE6Oxpbtfum/LCusEekFc5H9m0Pp3x9HhF2PDIoi
z9j5OEijLBr1iBjlDRTYV+r+nfaIQ2jFvWgFtQ389TbSDvezgPZaF/HVIExY+Onze5t32c6mxUuz
QWHNLN+1GK1F9G1pcnSM048B2xj9IEHtKO429PijeO60XufFcNK4WGwsZZZL9jZncLgUuLZ8aWKL
yFjqfjHYpTsQZAYCR74yzKEp5NJSC6OcutjCakwHDZF16GYV9Y0UAOcbllzMh5Xzen+xPo0h3Dar
LbBWoOJ0XX3fPeCLX66xc7IVJw60T66lDVjHrSZlupahY5ytpzoWbSUcuHa2Us/b2DcZacsj3k5i
AqTUcT8S9i44Au6+dlsv/2+c2GZOFus4kCszQhrgbb2uJmoui7Nz5RlI5Ib3df/X0e5tG4V0dUHf
xSypZvBQDzQRcj3bw6fJVrgKL4Rl4ZPlQlFUzrJ2oz0q3oweJqVBUSHfsyrVrTXDcFLE94KXJwxX
jUYfxhmZCpAiAQvrd1+KvwKjPbK+xp8cU2pGMcv4aA1jRaLDJdAzn+tIwmqxd9UJCLgJsfkuxxj8
Dy37sGUrOY4xvRRXAxzDB6m7/jMNYktiLgxjRhIdeF7+4l+tqbDKUM9qJEXUozX3NR8ykeJDgnOU
SbqirXWEbsXPBnZvCpyE8JXUIWPIuX5dkquq0LnnbcqXdNjwpgi1iLU/og6aIYA6CYO5ZPaXBYhp
JEOn1y8RDNmIWKtWDvCIm6ZO6yf6hJ5sCUs6G6ScXYkuFM9dZAo5M6caxT8laydmiXL9Sr5hJfp7
7fKxOAkfAmG+2VFmg51qQZ27E+RYhWc2EVL7LCNUaZaC9w8cXCB3pRUDwrQRUjn4pqrTL2LPy6Q+
7X351OWyfYU05cbFsJtJAMvqh1XykuPnfyl+0kSaUFm2dzi5f2Ubyv2W0NoGpvSjFEsW55R4JXEE
IwF0q8R+YAGlv4eNhJiD4voOEu5muUFmugXrRXrkec3Rgt071F15/RWACvdOkkxjg2We/FSzT50H
rDDEgQzesxwXUWI+ddaThrSHkK69CKk6WgcZqsBzzhHeDENB9QgC5ZnU7ZqYqCKNCu0RfqJ8867N
QkB0ZC1jKDcK3YN5W7uwaUBSASgNRyXQqkfX9WgPx/HbUXybS9FOEqI3EO9oDsmbLLW1Atl7re+I
ugo3/Fk8Z6A8nv7fizNWvexgEd46fLZ/UV6Dncrtsg62V8R8ijJONyiUsIVz8CxPVqoyUdVnLWys
V6hRaM1KstMqpAp+WeQG/tXMI++zngtv0DHGLm7VlCOz7uyer8jBYaIRgonQby6HnOcCxA9qcRAs
0fzUsdDx/f1lxcMvZV8gSX3tjdEDgjXS8Z50zFzdZOP/rYmeSaFlRuGeNlnA0Ys0KL2WTFqFABZ0
3DHpwExNUMMLiYdCR47jJSDdE13N9X3nmB3aqiyoqQVxDwuY46FtdzcjlmIXdtRmSAlXHg4wX5dK
h+jkJL6JJ8HB/TexVfSRVIsakzbgSnId3BAE3PEzrBhMv4MXWAbn519Uhz4qf/dWIm8BamhdPkvo
DAx6D3Ooj3r48q54fdWC5hzC6H9tbbaBBQXujFm0AbZw2lKEyK3zFGqdNioDt45kLs4DORDWUCim
1Nul0DsFPxtghmNM/azWdn4f5Uqd8VQvdwEZdBqgRNkBNom9P4zMraQjLzLlDz1WNEv+tzMPebDA
TVBlwk5gZMJv2mco04dOPzrKJvb/9Gt8YqUyfBcqGHN450Q2Dpzk4y/EkjOpMR1U6LgCVnrqK60S
GXmR7iDijginZRwwMDvRJXwbA9giqHdyfPne47lqpFGcAOz5uq8xAQHjmn3dK0dLUw2zaUuxzZt/
amRbKKpreb+goa0/wr3Ow/uYoYvtKl8Nu00FxKb9vUXOBNO/PCtitSxDjf3owAbC/JD/ncNK+bUV
hovt7jw4MzRc1fMGYCzRo+ZjHJUfI5bNSEacuPh8QCoZqiKZr4gn0tRj1XwQ2A33x87Z7QeyjeX8
dZ+eF6fHjvxzI6QfAJX7t1SzxZ9joLsFVBDLg2qGuVTYn8R3F706dFp4mHxecVESiW5V1oWtubaS
G5IMZQMQHnijZ4RTzXARlKpSkdPTMY/mi0G/txpI+xBxZqKhQBFOsBt6PN76HraaUiWE8s2gvtVj
nML2u/SlFtr5nYo/Lq0D509r9MykoI44siA8gRCNWEVCFPuB0UM5FWEMhKTt2lwvcP6sYV0M0TdQ
89ik1cBekknxTkUHCdaCZV9tMS+lwsDuFXl+buMvTC+BoLMRmLJo4umaxhFStRZT8LnqUayGTP9r
JQ58uEGdV1/bDLNcpmQvIA+zf67mQMXG6rsxMeeMcMJ91vI0VZcf4io+H/CwizTRR0mdvrZ9Rw+Q
iVlhZ1JhchHX1sTaDdfmpPPjiu0xrk61sPDZDIogvqt8zbycpCfrZ4T+L3cHNUTY+KNZvcOrZhq6
7Etp0VAjeoU8ygcz7RvL51OdD2OEj3gSiHchgwDcPQQAwuf4CKq0D0kN73OEe9Iw1+hv82UCANHu
uX+mOy7bv44Vc5Z+cteaDhD0rXBU53tfX+Oes+A52sznqp6VH0JyRekZX0RTI9ar/hZ5H6JIKmVV
Kb4kYLNrek3AkwvNSobRJp9EspiRUJjbLZETtqdiN9vUa5VtdwOm8QyriFv8YT7A8l1tM6MznxLZ
ro96uzNF0SOw8jMAFQYbWebFaW2EmnI+jY4xXC8A0ZT1/U6g6Kjgym4QEi8tehRko0qosPByskIr
iqjQqlE9AfC9Z/E5tPNOw/VRX/Q0muOio+P9B1xF9FNYRwV9pXyKAOFHhqLeSO0HfAHjWglhB99n
RGbmWEJpbLXzk/uEPso9oqfJ9yegu1Afcq+OdxXvsSUfYnvuqxYB/OKIzrEo6EaWwoSPcAJnOOU8
mOM22tWdEVlqkBJq0rHdZxLG3Q5eRnlm5hD4/gA3wDfT8FqBOXNUkZVWee8Ekoiw1YNZdRdf9Nqn
i5wbSi0mCJjHQ8A2HtaPxVU5iyJcgjEQYExICsqrz1RNuQa7gFw9HPvkMZpkc/ueidcOfPbaaQ7D
F7nOH348k07zCjh2i9BnMeSnIkYzQwkTQLNWtDYH6IV/Yh0QxpvXwCP1CGyTKzv9727dLbKvubDa
BbHk/l1Kmeoj+VvWhhVArjasGrg/AOyn8UwEzY1UA9N6H8e3gS/OBhQTmJgQpvFlrpzwA6ubFve0
a6QzUEL+CHt0sOmYIO0LHRxmtlGMRld6Tk1KmcW6AC5my/xq4lRxU1DCun/GYzQcnjl4ey8Z+Bmp
bPj/UQBNtAFROX9OdhHV06n8wmvA8Ahn58rnZ5yvFu/zguiHX74vE81barLMWadlF60UehLwAfm4
e10XTncGxiPc39WG/sNsybvHg8RurYz6kL7SYeM6nMr0Ej1fPgRGn7YBswmw/cdlr4K0XNHqxj1d
M64CTG0hprA+6GxyY7qRF9gKsx50mqQDIJ5LFaka6/l1UiNY0zKhCEp2HUwotZK2M7teLAOdTOXT
FA6UYlpxn5tyauWqjP1gwKTwwhuKxjcaXyw6c9AchzPsF4OkRVYOQE8yijadbJuxx2y5D2SfZrwV
b/idhPSX7l8BnfEk4QFFdIFyfUC9JF9v21tfZWLVJi1EoH0HJjht3tomVrabGhgbI8H6UlRPo2bq
l6T/K4NSOSp/V3UnBXTcIj7FcoBQ1NVMdsLg8CYsoVfkTiMt1P0dJmhnuos1AGKGFtY2RHhkd0U8
97n98kOZrYDyw62i3OLUYdH7L4rBuJQVopXful74Zsm+r9RJBhNnYJUvJ1U7Jk/D96sdOaa4xqa4
84Td1nqqvfXyZ9CZR1Tm3m3QspCz3Pzv+y6UIo9dyVgc1K2v/E++vwqsmyOZTWKaTCqpHZjGEH3u
ZwHY2MStia/FPPdUPlsKufymCnbjGYUepF25H6HicMGXwDM6cJzpbBlF3UG2+cb7BfaqIK2rbVtZ
fymtJ4hfyrJ7xXwtk8ceGwep5yKFn/HdkUDMCb9KJv2VfDvNwkYDEaKCv8Uv8FfhGs95knH6jWpW
0mAhB3sJqYjAUSSBdNYikXkn/MqXu4GXkSNUx4gLBkS3/w/sXoC0DWeU3Mncght7UzgHfKzbhyFE
+fW2Uo/2Hin2qhq3TSgMVMzKN9S4PozxbCa9jF2k3DFqxk9Twa8prFGq4kpW+us/azymXjvuefvx
Iqo2GuvKnZ1UkpomX35ZaMaCIyN6OFOmH9hN4OxgwFzGXsghfU6IHIUOQ/dc49MoLTcWm/RtADw6
hpPdG0CrdnegOd4WZNuDY9oV7tDyW8Bk16e9695nshUMJKhdWAkRhDJFpHTouj5rlekmKZD6zZnc
A3GRhp0Wv/8PtVjFOaWhzwTTXxpDZHI3eI8Qx6zJa1om8btrpcaHmYsfqezdXNB/8Mm429Bgl1HX
3pkn8vGOvycB7RzRm3CDosyQaIEEki8xkb8DozYn7xMkauNI5eGdw+zPrBKME2cw6asDAbQSWOc9
52PC9CEKddYbUn9LtHkFygDIVrtHhvh99rl4cU0UDjvMpjt7D5E+cHKaeQnVlYp3VP6dCim3NCEx
TvuSSPTPOpc/S/OtkrB6T5uGIZTKcuyHSU98dDLYcgvxX9FI5YZqaG8qhGxQODifMQ53dpP2pTOH
bRnSTmZuysmSX5XdoWYvS2p1qA/1Q1DpDUgP5GycojNjJpO8ecs3Yai2yCbNKiMZk+Vn9XIbPxEF
mc7yBbJ4tuG1qR+i7WJ9iwP36mEAdbhU9qBmCTsL3dgUv2ZjJcS1cGftVC4D4OqyqLef7AX8L6YL
wF8y3Oe0vFYr6bJuyh98+wy3MLKnpYoe2wCsXC6ahNTiOfe7YQLxsTKwj0zEJe1qKVnbJSwvJcwp
n40lGZPNG2cggfqywjiBSz9qkwWxOsSPLC0TNXrigOQI51jLz0FecgkVLcUZcK9Z0Op6I4jF+0Z6
OX+FHiRRl+LlniHscXoGNjrZix3a6CyghjuWjjq3j6mksg25aErMcSo/biW4+TP6n5HYN7nNnGDx
8SVz0ra70EYUw6cSz10GuIsC+wmAKkuhKFdm7WjNdNjI63x2BnF0knJT8zuxqIFDMvG2mXX3KxS1
9AOsTP1iIq/MYIpcuJkUbVtnGhl/OvzCGqFb+zRss7aPv9x7zA29dfeAVSWP01UErGRqmzALXF8T
szmJ1b29emW+yPU0ooB/e1QRDFd8yTWfbt5dbKOUmuEu4vjvx+QLcy4FNE3/HGgAWii0S6p/c9GR
GLHZvrsGsvXEz+PpztSmSMc3qPJAMVIm9sG/HP6iElYf1UrnqDf4nelY1ZcQIi2BbSpfK//yQL0Q
Ww9MIYlQ0lm2fw97MEHUvos+8XbxgTgPuq5EDk6sseCGTq/bPQb3FFJ5gtWsvjNgrfxtcJXcUP/p
+nrGSSP23ilgW+APCsdyANQNS0u6V79+etLEc/cePDM48GfIYfnIrrsZrwvwNJ03Ls7k47D3moGh
nRbPHkPFBAeqIUNrRyiP7h5T11gOwMRfk1UjaLHHzvsEfCMYLRM6Z7RY1fd8u6iovduJImfuMhqT
SPChesdURh8cJXh2Slub59H4fj0R1cTqL5hCzgURGSorsHjEAkki1thwToCKj7zlfAtPcaz06tnB
vrp9XhRhkfwjHEhzv+Wfs0xw7Qwt+sDE8NFpseMax/iuH7Vhc6x2eivegVRO+b8y57nx+Wm+6v6K
RncI/jbhxKtWapv7ffatxKQ5vnTqPmKiLJG7LLov3Bq63h5pRsGxcyMTcOoyaGTA6BTpBvFQPCUn
L/yqUcO5dvF9PeW6ze+22vrTM0X76+P5gFmeZLwzHS/5obCbtapcWmSiO/uzN26tWpO77OY6TwC/
0aSJWNdeu6RL/KMxhq64qk29bb+1ZLPoCnvFGRLmvcETs2E/nAsNZl7kDUCotlJarOglmcXqdnvi
hnUVxbBrQ5A1P0jBBvuS8Pldb29xNN8QwnkfTV+bn8KS0ZrvXrVuJ4blgj0IdE+8YOUjSGmyUSTZ
VxQUSm2uz/l9EsPaahYNZR6zjPw6C3RbRQmrnjnPEpnG6JmtQkqY+b0D/tToyPMdMSylwozbkYhk
bXVKAFPDWrYKVJPJ9WXf8r7VrNYbgRZhE1rA2gJ/49fTYYgt2G72N9fPpJhpEarn8psp3InFfqvB
/Fz25HL7Wk+0Ym9nEfN4VYRP9NKWHOsf/uDEfPjcELXV+ZWHdVdpNCMTcma7O9thA44mixplaNAU
TONN8ip1nwFyPnrNoLkZgE161njm+QDP/8+0TWhfPDi+t5h2+xQxt8TQPIq3At+VwDIC1eWSEpsl
WbVIqE8GB1pFzR52VHjdcgzdLf8kMpjdqoHkCHjFEPuhOVlatBWHKBwJtYXu2PG1gsu1TG0zSGTY
fMgfGwjhFBZ3s9HFQUAtIHWjhRnYqyo3udFMxeKifRFEp5qZH+5Cc2O0uTMMnQfqujdS+u88/8by
S1779YvrChgeUIUgmGNJgIwJmGXNeClCVlrNCxnRRHFZbTTMYyuvbGEeh2pWnW2Xb5gCT/yvL14m
iu8NI/QBPujcVWS324uCEvFPZuysxu9De6HEzu5agWp2W98EAdbLUUxpNPwsf2OBDnmLksL01i7F
buGzXMEPWbD2p2QvmDP/EfrnQnRbQf5JzZ6JHWI7p2G5jbmfFyGmI4ccnSpby7CkQKZ1vwI6z1vJ
gVYiPM2lRHGJz7FyPZXu1GoOruF49X+w1uRv4h4GwMaFScFsXExHSPKsfmhmyTM7918or7nemdGl
qs+q8nQYay+xmaqEBOwjDYl1i+sEnaEUmFyUz5udVHbcf2fnQxiKKP60BqNci5XG5Qjc1R/mVkCH
6GDIyC9YamHyK6GpB2L9zxsBs7Rns+B9WBJnqwCezKGRNTJRx4ks3uqxl2iuJAjgDbpstiRcBzBp
7Hbtlg5/tut0XDyK4rCACdAu/PdDjJqkhcLxpM3xzcWE5etPcXxg8l5nKnHeKc1z/AD8jmb9jlV6
yeaTnAZB6808kzpm1OpSNF0LPMiD2Jb8F84FjRoJoyKKrtz1blf3ugeBrub0Xusw7TS499e45mk3
eddD5qaNx5AdQw5tc51XAsOQd8xCIG1gnnRpHF9Sgu1tBNZ5zHD6iG5NppwjHfBShOnCAUmJacvt
Lbqx3NAdgxE8XliTytRLoHUqI9KTn4D8z/G0R5eSoVJPe6EelqB/84Aj5oYC0WM2h2B0x4rMFG3s
24+Jvqr1lhNvMQ6Wp2qk8YA3RSBT96uOk8N0x2ERgus7XfVbU0BgV1ojRoMFXKxTr174Pg7yyK2O
Sx3nEDdIy0XoLtcIUCyo+emf1+e6EiRUwB2ubyrcrUH8r3f5B7DMp7Ak92WfFhVOZLpOSmmCyGB5
UXNsWiy/WqmY04KDATOGhVQv+q1jz2i9cjWTn1pZPhSkcnsdKmpzw2pMdOwPo8JtX0ia+VLCurLg
dvoEd/tBruksYSe1jWHm5DLuPhqs18GdCXC1bzw6y7Iooe0LEnB3lahorT+FJm/+W1YtSgcTzzym
r/I2Z1Q1/0b4H/qFZ/UiH3nt6Yg5YUi4KB0NLnZtINWas8iNqDoe5b0tZBVhOi5AENdEuvF5xF88
dnbCQXbJHGqU1T9CotN8MrbGpQeTEDOWM0n0of2ikrb0RhEotfPT759mhD4AowyPKLgdWoUIbfIP
LMaRnZzCEW6n2ySP7lRJXivMwo/oLdwAc6KaR5cT037ZVswvGmTmW9MM+2zsdMzvfZN5QT6CtuTj
A03hT/A9oBdie/eCEZbUrty4r1xKFvj5ANuJ1VwSooeTyY7F5ck+VRCIANma+ef6kwGyiviK/XpT
VI0Vkbp3TqefYRoQNP28YhReIyEayYNNtQXP9Xqh6Dz922pv05J9Yx6n9W/R4dhot2HBn1nS79B2
HiHfkBX2UhLzkFBDyl6wnepO0fQnIRvkRl7FZ+MFfv6TnGMpjLttac909+GL0P4kdpRiJ+gsvJcu
7R14vm3evzS+vRPlLJ3runGUDNjF6dzwbhF5R++grOVJwZdVgi5J1e2ZITYhhN7lWdde/uMyQWti
IjAYu2Y2F+DJxt7EzTWmh0Dfysy9Kh4ECVyzr+UDFRwYCg6vAofl14iLZRlDyDwaMH0shHL6oYsg
wYFy+nalbjnxJx5mgCCP4Vu48iYyo/qESw8+9PlkIczusCT4ly/LazUKibL/WVAm52HYT9pzZCUQ
j4/h4OiRdG8Cb5tXA1ZzH9QI2/1WFBIe7QcDfobcJHxM/+P0vD6gkb85rJrIfsVGr7vPiTVEsYSb
X9LeRKAPh9KyILh/lQFP1wR8/U5lq8f27p8VhyQE3MDT58fyQabmy0TO17HnjsxQp5y+FewJjsU/
+pumuhNZT5O726rbqcL/3VfChXb9puxwxBvxdinldbIWnEU+ebdbtKnwsdfqbAkNYhjRhQCancOd
aP6IvR3dBKImxyog7v35Rm9k0ClNSAZzeT3eTvKU8Dl18mWFeamAh/meZAVOPuHdyL6PVlq6Q9ec
x3OdZXM9xH6R0QI8j7s0aaZ9H39xmQNWiTjkLZhfiHuqX5SeC98dLlTXe5mhCTWZMDV/9a/GxZF0
gdtt40w/vzEWUCEbKXNJdrzrquU8HesuDUbzXasOWH0mAqfe5p6oV0WLWjimVcwdBiiRZ5XKzWVc
x/WvTBTqmq0TRQHJOb3I47H2St/ENM0gp5BqFYpSDyWaj85Zjgr4xTIL8SijxUpSDdaPabh1u2P9
Nwp2X3xkNCXCeKT+ZNLcFiy9A4g8OVMsDPFxrM8wKL9FVtBPiEQCONo1Nj1K5+if7IhyDTssVxRs
cmSSIRpmYhT34Cw1gnicJZ4XYVz4SZmIpQFVNfc/Vj9nllxg6H3K4pM1161MD/10hc/XQh1plZTO
qlibgei8YO3XyOSZ3nIoQnnOVnYpifbMPDjTG8q0as3BAoUF5Fe/jJnz3VokXZ/ng6QDjUZkqcyB
Tz/ILSq0KBAziZetqsE3NGc6+ubOEQDmcKZ2dLJDXtHfWLYeQXKrnZ9Pb/UV381cUOXWLo3E1gyH
m7AsBN+l6pCNV3GjB/twAivVk75YHz6kJh7lBbwuuh0eixl3IqII2tkOqqhpcOIFWi2ZlFRmtGJW
RcEF9rrDcsmCqmuv8Cj8ou5knFLHkuUH8GOKNo/cpbMGH4XFTU5kwcUaPUlQT/NvT0NYuHX4J9oA
W1xyJV9Jn+5eI6DmLNiYBCoLVfxee9ogwzKLFps9jev6c++FavaAeNiHDlrgCcahLFa5yYGcoBHt
UEOQl/IguqiE+g0GXZ47ExTRY58Vf+o4L5yXwOjTSufRFfosljeqBTl4hgAnE6v7p+mk9g6mQH7F
LZnG5hgWIGT9JtpTM4ntohYUAfOz6GHCs8zZV5Ww2qrE3TrceCKWmJfr4NUlNoBgN1P8VmDvfT8Z
kDf/kBspM3qOzzYNwMAPePDg2H0WXWozK6NJXV9Hsy5YpW1p7mG5mC9TISVNPDQT03sHJ92ENary
RlGdyN4Or+eMX/Kx+thCdwpfBy7n7EKQmhEGscVwwzBSasG1Y1rwRw4U3ctnGnp9goScLzFsOPJD
AqF/Jkw2otbhkuP9yLA3bHQcskgVzFvKxJ/gr/FEy/KMzY0mJ1LRC6q3wt6e+MNtPXi4vOAutw3c
3TSo3yFJSKfwpLb4DjljKdRM4EmT1+j+SQOwKPqf9Hozjmr2MYz9dvBaKMMttErO79djrjUlwyYW
oRi63rbJti1jrMzLQxSagZNprn2K2dFZ8mz9v8mMyGXmUutICApuU4HyseYcXBxpSvnS/KXJIiDC
MLs6X/y5PA70wIgBLb3QECOIKWR3zs2oELGiwAM0HfULggFL7HtzP2tCQZrQk1eu5mfVCYiGQQPp
V9GRxnCnmstiWLo1tCgSVkN31LKsp+1/PLHkDGY8VapDcgSefQjRcstUjWrzSU8wJbYqU1bHh6L5
54s0homPuV0odfyrTLBqm84kgu6Y03JNWYz2tZYsbVXGLEM+BRj66BFfLOCcbobrMKMCYMaXnf0m
lfYFeVj1nW+Q9aE7Hwm3ASr8mG9T61Yhll1xlcc/OfR6JnOQuVqbI9AD5ek3ca0OqrTeDQRffpj2
T2kE9rEdODj/+0S+4wsxn49sFoxwvDMddl94FJKQYVibSyStBc5ZX5sICScKYQqk0ccPEOkMbZ44
YAkeFpzp00U3Hwm6Rtry24mX1b0jJHEjxeHvERK7JQ7PmY4WKCpkdXT/rCNravHZKRl/NF9QywKc
lkfoth6ipHk6QPFI8VQ4SzxbolrAauo3UmSwodlNqNf00RcsD8tSfcl1sq4GmTX+cgIyAoftvyK9
Q8zVpAzBLuQfJi/fgWD+ZHXLhlp1Q+vwsiYwTibiyJ+lIkTgGo6ZZsUlJvBLQN7G1LmM43lDwKho
DnrOdcYPEXaCbX7vAIT5GJyoMEuj6HjMmLkgJBU3M93nExLjqrnlweerFG0QmEEB+LnS6LBn6/ME
rtt+qUgsF/IYRhQTHnOObVMW1CCkw+hjJuRboA027lbZ/kYk3kE4LHzgrRLJmLCrgiPyRYJoQoQz
5x+tCxEceSFQ64BYdov7OrACBS/TxDE8LtiHqDVovOjNvmkqdAKP92+LtFGlX/z8fFSPv4EsSwFZ
DKioos1bLTGwcZzhjsrz0wNlHid3LE3UiEs2Csao0qGrXJjTQwdSra8lEvHeF84D/DgbT/TRAk/d
1QXoK0nHuRQektg4fJxacMxcPDxEAVw1rmytgbt8JfyK15pqVTh/kR9kYFSp1xT8FJZqMWtI+P1U
1F+XEfRV0/gUtIceGAOmhrSUwqO1DQpbI+I+SGcTkJuWCxvvBDTo0xNbLMuaUTl88AXaFSsZ+9Qw
ACleS4qNL3CTruArLFMoxVUY6uBZ/slcMzP51Bk0yfMSRdxMc6Cl6HKh+mjKgvnPteN62MyPCxri
cBWIq15j6pzEEplAbglUbNqSzhH+dU9j2gzhk5DWrp42uvOuPWB2v6Yn44BIzMGCDvLlzBGGZZge
+Mdm6+UwhIEPEP4a9PuAGn7nXNxWrD42ITVmDAlW4zuscFb0ecGnG9m3twPz3kjDgBRfDcaAEMgf
b+yHFs6KIXq2ojYuuVLYg+2cxoBhBDxAvrTsBiQFiykspRkwkLv2FfEXSotFj2MM1IetzQs1BtbS
qoxCneOrrD0sjsW93rdq/NydnPzBSGtRTZstTqnWYBuZJLQCuiGUZhJla0hN5LT6eXgtMwOti2K3
Ey2CwLxAyM9RDwJDmnnNur6lPrI64PpsMCrbi3IG8ahduNihlN8pmEN8570gJEMzTUI3pahXQvTH
6E6wke6Lyjc1OVhD/yvyRvU5Zy9TrT8H77U+1bF5iZFKJZAY+BuM+3iSLhflG5FxvqA5dDf9MEZ+
ye5BzobpNsUogT8qElVfxUnHfMqxTXJ6/rlC5Ozkg55q0N5JEMRomlv1ZpgD1ZiI4F+/m7mWHERd
Vt8UcS4nFIhmR5zoJ2HPEqZDjRp754ddEP6e3SQnBA+SN7RbyfLvxQDsG1R21cItcLMOghZu7Xkp
Z9aKWRTufC/pXbYl8ye09WCASKwrOQfUtp6NkYZp6qyFSKWIfvgF3DxmJK34no+fY+edEw9/6WbF
yZuxxWvrlkLIe1wEkuoOFDqxzB/DNFapjqQzXJOoSfKyM/oOfbGPK0c+DN6TAf8rjaXtiyutaPoB
0kGpR3NhYswacEiUx9JBqP/r/OeBc9BPieo7gC2epD0eYBdE6FPppIBsvJb6yRcXbZ3ULOUtKsks
3QfNX2PqCIqnm3twubNPt1+wz0aKL+rv7Oh67jW1wy8t/4YMo2KG7xBF1HdpprJS5/w8PxGLeWIy
tZinxdEsqNAJW3HQO/CF6htG16MRzzm49bRN/SXdwTJwtdGD6nCS+VJW3s22utAw0i/SWK5Mj8o8
kvIJPh9wqc7coxLzRmQyfHcmzeGvsJi/hK03x56aeibVfaKYFP+gsROzwAIzILWo4g6VmWJYwsUj
YjupyQ1r+jyFKpGZayxnxw03GBLpers1/p7rrYP0YcyvApEqoSZg+jedUUkPakXVrp6zlkf9Fbzp
afbgT0aSRkuBNJoYlc5vLYacLwFP8FwrwIWw5OUpgriB29nrJZ+au6Z49Rc7vpzlmh6YPObTb2o0
f0pUtIEdEzkcDGMW5j3STXc6AbWeuOic7KcvS72WOj9xBrBqtwP94W1cxsiT/z7P2GPdv02sTW7j
DqCbGuGx10s+fowLiocr/MCyuBdYSnWGpQKIDa0f20iSnDb9VgmRdTH9Z65CDKWLqCw/N5tnRhcM
DtZdDn8vbDMZzyGvAe9i29tTrKpEx9I4VuSk0FZJCYDiD4QnaW/nJBh49WcKW0jbsCMryQjdt2WX
kjItrvAg9O0mFB9MtlonKhvIrB64vGjVdik8cA3AWyQGL6pbc6gMgQAlSn+EGdwCm0Vk4CMuQO5H
wXgVPhY4KQN+Z+WAQCPOrI923xMyuV3E363kadjFNZLQ/q4BoaVVMaMO1Ov0dNzZEuFWQXnEySFK
0bvRUZZHlaOBdJ3Mb4pM7RA/ZnbRI9fU3+tuVBesv0unlbAPemlOMJIrEHGPgM7dSxUaMU5Tk5ZV
lSMEZhdxuHVu0cAixeu0bkWgg0LVgD58Bxx6JyOBkxSZ3ysuWF/i+zoYSc7XDVQqb5IujEx9hrdk
Un+VS0gnI5L/6mdNEYfBNZu3C7kqIih74iH43PT7SkvBv0HyRQJ3GGWPFSSPBJar97NUnD7WvtsR
xCI1wsJsQ9kI1M6Fn5Kx3ApNigBUAdp6eeu/Asar2Msme5OTEoakU3FvUUeGZ55lc24bxtiVhlrL
JdL+VnDpN/fbOTYt/sNfHSHRdenjZJaqeOVkm9YqbNACfJGD+MpTt2hRw5/VY5okrjK1hdLgW1Wr
rzkbumSHyEcaHzmcUt+SDZZ4cKT4lYlY3UVbCMf+y8HPSqtcUo9/P5cn0UTCG6/VCefsAnEqDPcf
s1Zuqr/1yBVD0a1Brq7OS7qDLPNqJ/m5P30D6RgeyqBfjZmcVLjvYtZuXcur2v/He9htFq/LDDUY
WOsb8Yi4id0Z/K2/xy+diPWE05nDWq5zJ6kyDrYwEOKIcsW1bCShaSdDqz2alevucJbwY8LOW6Ji
Iz0mgd7tXl4LNH5qeQrUCQQhrJKLmgpRPUwJJY0dQGpWrGyPIkH5lUmfKM8WPXS2akJzZfB1ir1k
QoCwVV8GAS3LsAouX/2BbwC+hoQc6plz3kv25E5//ntnk7nGhQ7Ksi+iGpgvWK4gVJCGm7xuZDLF
0Gg5mJdclo65uWbmgfgGELYlERKmSvN9IsbwuTEIsbc0LyU2YDpOYlOO2dM+rN1/XRkVygCaSzwQ
2CKQS+7wFp41Jl6Q12vfoetd3hBk5FmzRDYJiTRHDhDpQnhumSjLa09Z/4Ed3azQv0guqjcIj1YK
xbm3RsXBG2CN8EFdhCw5tH+FTRiBTnzUwVKdZMnMTvoiKrVl8S+TdJqTGOAmfL0R8jF5ZSJ2U85w
n168rKWmUtAKgoZJWbZBIa+tbuqU84zo3imBJFQ4pPKkjc9IcoKdDoN6uWgIXT7JFgqeBnxQczf/
1SKBacYntxwrgRVlPtHxr/PYGBdU4Sp/rDwFh6Q2jA1dglR/4kX9p2OFwKaqOYrdAh6BiyTDFiUx
SDOUVzGw1bDV6bGL1IA97by5f7NjzFo+SZaE83oPzQHLjI7/++owz12tQZGXxNFHkV0oNqlEXts0
9YBcL65iih77dYacegrvgmyo77VQW2jlln2KDGBwPDG60wNKo41dqa1GvM6FRObEYYizdcD6YjuZ
g6oO4GuEm8skulzSZZZl4FD1rpb3e0K5q+s8fQhEemeq6+izk6y5hquyJd6UXsCaazI/zusMc7QW
qv9mJEJNNpLKQCH/xGlpp2QG7t1EkPGxH2rrMEgUXazFOT74YeeqZaLw5UkZEDwzof3VRCrhk6qk
E7hMcblR1ZPdJ2nYY/TVMeXzrPm0xCf6XIa9BGjQnfIykYbNSQuS/MvZ0MWuQRyBHWnoNjHEbpF1
SzAMCO+XWmXx8sjMclAEIQem/IJoN6q6uCtG9hXyES6WlV0xvgiXABI5u6P6hNwSV9TrVHQPSO9p
3szy6hwPuT59tIIyRLPig2w2E3Gy4y40xvcal3cGfGod+wPVlarh+hFVxPK99obOny6hizghrgZG
j/18F3sZdpi2BewyV2BJKTkdpZJJJsjGoK/5iCZ68Xo86dU7Ds/WaTruqTOzHEfPftivHAuhRKxG
LPymoOfHLryadSxKywdh54EYHPhWAzJC6qIMs6xTTwI9RxbeuUbsVVsM81T5fHa26Y5Zkvya21N6
dFId69FPyRiSS7bLo2b2UYZmgw3/bggDKlqIt+6rXJmGHW2tyaB8Rvaa5GWL/6ZzsYqP4sADnNru
D8wCTjKDs/Ls/ImC/uV1FBlluL5dpko3sileNP/5Mh14MUj3DnGbY6eYEqyZCJya4mCVbtqx3YqK
FLTNUu8yz46EbMMPIKHydgMUlJlR2kYJ+apCCLHinQ0W5HU/iteNCyFs44xaRyF69ye16vWs2wzt
o59xcVt4OrSwtKH9LLz9vl2y5FCZgp5ea+kHoI49aFGeVNU77ribhiRt9q6fkYnBr3huWtfeV4GB
wTSUNZyAKPKjjGwcdNRNHCLMADL6K/xZedbzceUSpb9iQtnSoUWX3gkuRkgQfIjbow5yHOP2pLPM
9jW0kvjQC3CC/7V3Q3JGf4Q6Sb1AxR/ttEO3r/heH7lC562v1TJ5J29Z1f3Qey3nwxbGgW5Tx6tJ
XvO1kYjPa+VXadvM1VbEz4yG4nQ5WjRCZfnRNKFWGbsBMOqOCl/69t7Oa/YjqAVlXes/+u8h5PZ7
nTY1x5+zixWsgVnjF2EoF+pp4UkkPY7OWecmJpRTw7DDfqFXo2HaoQEVJFOjE6B0w3eK1zApC2HH
WVZmJD2OiQM58k3WjaEIOH7PhizWVC2HVc/3nYmmI0i4SkIFHt3IHo0UkjTHgsg06Fpf65fdcRl6
J35i1p5x6CjOwW5xphTXLzu2NpYU0CXxTzhb3e2+plwuIoNDLSCD5sCEDM+ibkp7sgYKfnjiqyvX
P/DBx+SV+IPVQBqwtsaMAE+7w0D3hAzUpold+0IBM01e+3NCJ7gF3+tqgmx0TrEK1hE1o5p9IRn5
2T6+s6cVI+GCmBNrq7Lz6YXqWJIEQ6UE7RFNtXhlWVXXVKe8Ycwd1mROniOGo0aS3LalIG1tKXUu
xetwwbBLZWU0jtLj54oxTIL4WsGOO6xk4hyC0bq6l162X4S/ON97SYFHaxXvGxrsvtUsNb9FtAkU
HcbK2C9B8zVCNr9KKA0J0C4pWlee1vBEpooD4kuuYxnKtPKFpIiHEuvNhnGNJiB3zM9rO7ynxHFd
OxoiKMV2+9U1iusGXUKOY97EtBvdQVf8Y7tGB/hD18nmJNwPFs4+aa2N7aNXgtlln/Pnsgfr1tYz
8nI4EIokoarRqu7CCukJtIHtH6gHNYCObp+JPjIOWgQDpf6tpMDVZcUNcIm/gfdBobp4apjIbpWS
QKBdZghiMWzdBJ4KnFFMiyI4JGi0h+7bIPdfiUpx4sSSx8V0vx87pgRtyhvJG/OiaNt4wrzNEgLn
//IP+q35+G8AcuWZxVv3Ij4il4LP5O10Lm8cKuiOOJqDLhuQSu4EVzQd75lm4Ox/PUlFrSPzXjHl
f/CTnc+loXKYfP7dNgXImJ7sUFweSoUs8VVNJfEpo9qaSirV1Z2g15AArQ07k+xux23jvU9FbvcM
TC1BbWUSaRcyiFVkyAnoucLsjQkJ1nkxpnyIJtJzETyayZXYhDMTuunwPOdIOuzngwua9245PC/r
f/RH0x8Cr//kMk9dowBPyaljnUs61LGfpGRc4jpL0PJ4e7hAWQyasJP4/9CDivJZcF0T1GDO7Jxx
7pqSE6hvhdSeQ0L8A8WCU7F1cbcvWXduvJOhEtb7J7NP5eILs+3pjfDSjanlHH2xUX7dFgan1sT/
/kqGHmbDqmOlgqPl+x2UYn7PqxoUg0bNgJnzFnz9GFay065QElAow7l5FPrlMR6MorRy6JnmQCJ0
BY3JUyWEdFuS7WT+mrGs5GYKjradNd3OpBHjf+XdyVrS0uP95MOxlEId2AXh63ZPGPbuKzSZBs3u
+B7M7YKLLmX7pxbTkHS4phbqdeJtsRH2REbAsUbsX5KM2gb7vaahfJu7K3/994tgMTnrdgwMZPYb
YKjXOORTwjJ/HPM9GTjJTUttFCQkjbnL9jt0xwWQ88C4+e7Xd7Quq2oNC2Jm96XwLq3/y2Di+4sT
UB8ijTp4ykvxr0upCLQ3TV417X5o7fw+YP5DGD2M6YkdRG7Vom7oDRzX/6EjE/xfQ0RNut/ufqoR
3mWVNSo/iKozHDd1Urm359EMoGZEvSPYn5O9s+5pX2Ab/yjA7aWV6RGMGmd2/S9vlOm4OD/a5BAn
evUAUDXWu3Q8LK0etwHsH0gBhGEl/MX8ZRLuYiwIkJFctH54756SfJBCLFJNfxb4KT+pRdr/3HPX
yBCM7HKQbMGgZog/bVNco0QSSN2VDcleqmHkKwg6t3EWTDXoFjK/Um6QmAZuz8UHWxpPCc6/n95G
YKAjcWiRo6Aj7X0Qgy7t+iR+dOSwao4mUpIXrRGr+RJ3meBUlYZzGPDUZYVBH4DXnOb0xv7egyUn
9dMdN8WTBywX6S3gbmizzlswaRxQV5rBtNHXXgcxZpxajlgOs1bAN84UzfC9qN4J3kFXYAHtKyNy
SAnEmaoPb74BeHHl/IQHjb/XlId84IcTU3dqxiAltFKP5VbMNqV95N6vX2EfujXKTeg2wPQok4cg
DfSGpDHmrZunuyJnrQaQtXQuYVbwZ0D9zPFcGFX+2lXHyKmP1FOVAKJN5JXI4hgGlIkQZfSYAGED
4IBSYXxTtn31FpdpnytURc9T9KfhALmmq8uXblYdImqjNFmJeRUXHSbMNtQmrE3YNi53yRSxPFXY
+3irgBLJr79PmJL2MotkYFCpu/3++xv2tqaiAakb88wv7/o4x0yzO5L/BPCeXmNkBN9Fo/4UvjXV
iRzIs2SopKSbxI/utS1TmnzwgtgW4rxwsl4q0hv/lPOSLpYtYFPN31fF+BCul4JiF+cEE0AdSryS
uVGWP4ulufKHLnuW0RnlH5Ne9stE3xQsPwl48JTbX4O3VAdQYNBRaTx2UVG5U2N/ucaQfw45R2ZZ
Y/11qDKEIf1xLBebhRhirvsfbegich8zXGmUmSXpopaE+AR9CcEkRqiNfAJKvUGGPrvKHIvTLLlR
AXgwSdkuO0WaCG/7P6RghCJ2DXWfKJ+OdhP2Y4Z877a8IYm+TWIpHHzwOYLohwljXMEgAsRUYoo7
vxSPw9PXQ6xL/qMr2ryt5d4BTdCdmfv2AAgqjIiXfXltH6kGUWcLICf6kqr2OpNRfTHdJUVOKPWs
9ImXPnkZOsIIOUjSwdDbs9UKDq19SZjvr0q3MTEMCkSAgcTGu+A/drlZXP8Z+Q+RBcAge9R4DDjy
ZrGEjrk+TyPSsPfmwZaj15eTc9GUhbvyNk39H5PZMTU3bMhv75vc769XdYXwcK0HSkU9zhbkS2f8
pTefefdRCrufbpfJy/B3LG6w5yPE/OpjxozUSayw3i9Fit38dC0TKJRk/A4pLAFC2UvoOne9ClNt
Hzi13QAdGDVWlKstEd/q6rD8mcqa0Um7nQBaVy/aF5BGeHkWXj1LLE3QIGOKQW7kZa6VUBNxxk/l
SVtp0fWamZb+sFNfJAlNxJ1jt6GhAPjGrUXjLZcIAtyZp0QKVobJ+FicqKIRO2SzJxWZSBMlFOAr
14V5FY+/Wpz6JyCBhEFbv7SK7W40TssS1peVmbQoQ0WwKAm65/p3BT5TLcPD7uPNovrpUawmBHbr
skII9Z8ITEIuJTdc7IiOHl9rCpH6dTxHaaDjOU9pSHh2ezk/47J0uomAYx96FolhVBOYfUhc/3s1
/YZ4HRkRUQ69NHXCfdbrA5uuM5BUa0oksBmukKt+vBqBtSi/Zr0RQgoq1NDpsaBpOSyiL9dZZAUn
JJy5GSh3Pe51RVK+oItANyi2KLxX5WZBi4/6XVuXeOBElKStu4BmPSxKhVyldf4Jgpq8wJ14fxAx
5/hzITA+kWXzufdhglUtpMDpdcF5lOCEMcQo7REvyaIHCQuxKnzg4qSHuUZI9atQyTOA9lnOq0sE
LtR19hjwqDM7wD/6o/e8QPlLv4iWyTye9qZ1rdEzWe+oFxDqgmg19YCjtIMvQsq/pqkVNYmfMMCg
RavCXVr5CYg9TdPGZt+RV2RJRyBwFrg6cFn93KUEePVTI1NSF6OFiEWthPfpcO7zZdsT2DSfa43/
xgC7dgc+0GwdYZvC6zJQBfUlLpoA986Vgl2Fn8brstxMEpA+umWkCA09xjjdlDgNwx2WYo6WFtrx
i17s3toKtUBVHlFuGhOXFdRIADzUGkdvHBfCEhFQFMZXVX23992J611E5b1ZP4Y4zQagjK83E/xC
vtr42AW4VAE4xqCpYFniboWYrZC2lf5UkiBcj72pD+gmTyubxOxhcPlrfRbfHytdsGN1/RrLnv/I
NDPZwsLNYp/RiMXeYOGBR0nKcB8qc7hp9hjRxdKfNVzhvV52FityH2IiET5uTfvqk/drYLT5fYD9
+UF7VrsbUGC3TZMgj/N7YcgeXHm3HM4LQ6MVcP4XqwvsuJuDWt/nJ5stXK0sAR7Qx634Ck3PTdFJ
yXKE+6fQdFZGTLs29ekG8ezornBLNd/Z3uFgbBp62rMKqfcBmf+4LT1+uticA1u5PaIN/E15d5sz
sepWZ3Xk9ywFAPRV3tLlg6Lu2A/Rta8C2F9LBh2O8Ynn7rA4hgSf3mcD5esLfvY0AV9dQCHBa4L0
tfl/NxUTpvKS5X+lrALLwazKGDcQSB/vjePnzZbY2J6IAlFjU4f5KcMt8b5Kv3Oncg7eim9wWuXw
loHg5dz4tXbYeU355EJrrC1eOl6w+ZKHZE5pIhrJc00SAMhVr+OxVQCSkr7SKRUOqLvX4dvrsPsT
8TupaLYeI8N0oI8OlH5k5tGlC/rs+VeoKu8H5PMaDJFHW350X3jPdLWxY4V48RSVMnGaa2J+bLSc
51E9js5LPQZsOox7t1vEGsyVRtGQ3SFFOy/cPvAWOxVVS2xHCZvNcBIE2r4NA65XKjkD7AlHFVVA
tAn5A7R5aWwiwvbYybBmNwXLIi0PZfSG0WLUEUJbofjmMqJn/A6UBMSm3Ba0EIkDan/gEfrUP81N
DjEJYxNjcKfRReKN47DvQKOg3g3s1al0ArYHTjmXlxKlAUJAMb/T/mOS3JXj3csnOkuwiPO0Qt+a
DajU0gbSKSJKPqcznKn21jan8m6p9cu44vuZpViVGiwr48lHcKnI6anEzfVAutiCJRv7Zb1rlUVf
n/Cu8B3elDIa+nfl3EzmfTACyOORgfMqDxVayogu++2v2YzdrBozaa5Mfp+AiqIG3MUAW6Gjdrbt
lewNmAsyBSpef7GazrmV1Gb+VV7oBu80Hm1nxYX0pO0MxBpzL20zeYzkipcEO4sGDriKkoXYCi7Q
BgexeQxZtKx55pn37/t3M5pp6mDgdyDJjf5BnZo1QWVwY6DN1ZLhFmwoW8A5UnTN/qdoeUdrPBCK
KlWPGX51laepyabVcNue/5qcC/ZageXr5p73c6u2QKMJBiBS7Zpe0+5YHueYvCGrAHlBZ0ZN/2nK
U6VIiAl6HHCbjmNF7/C1Xq5JtFzXsmz3exSr/GLPxg3M9WQwtc6ZmL0OWk4cF3TgcDhUHfE6xIwa
bSWZf+6BY0BRK5DAHCWe98Qr5YQtp3GBVqC89Vfj/N2Hnfb04RV2zJ8Md4q+MN1VDOBed7j7QWrh
7UwqRfPb8C8dPKAg/mJt5nLm1tMjRJxUX3TFyt/kVmHxRZ/oTQ7bVPwuxSJcDnyAbhCItKn2Mn33
jaucdQTbUXnI7a1aH+bXIsdnN7UHvSNDpeObwl/2buCRhCW6CcNEOCVu8DrZPLKVpXxFvrNZdHe4
APqURtXmvRnQeg8Iy0GzlAXx+2YcTs0yV/N2m5MAnv8nkWIbJLkB77vSADcliwRvt+NPrSC8R0GV
AGh8KAvM/daRYk8IE0TweMCKo4g5O9sNGbQEgAILN1KBLl1wZRCSsVOsfN00wXlFmWMzKicjnQsd
x85i1R6sCrom4S9gZ+1NWRABb7JMhVPd/CtfTGe0yDmeY0LEqPMsNTmY/38MPl9OQcZeY3vIaYIt
zYfqDnPp7l6r8c7guhFT504lzqB4sAdToRcNdAHcBfu8seIvJLB1Ob0bXaDRTD4xQVILIRX8uIvX
uPGuV0XOSABC0n1Kh2GP+D37TkDyBGT4CRFxJQUrdWLDMk44MIFR0jFdxiBvo24JEwBz9n/ZtKyM
Si00YThMi1+Hb0KnOUolZw4/u4DxJPGjopghMTJJRoZoEsFpUZNhkBASxMDrPZPUCXHFxZSVLXjZ
Is1EzJCzjZolwNGPW56HcpktOue73exHZ85M0QWCK0JkCiH5N9755tkqBTWiMLBo8fV7b4Gl2wrR
wx4nhAhSXMBuDpb75xecX37THCzY9PkqrdgUR1F4g+/Kc5XxHOxs67xtLmtGuDmhwOGUixPDgkc7
wrEoX4T7wekHIsSSOhNdpDv5hk1lANLV7qxA3SBkc9S0RmLbosjOq0pXUIOEnxjU1PdAnLF8SX08
uAGzZWn126LoTIY4o8BC5fhM8nXhJ7PSEpy1zbB3Ekg3SYPE1Qb5/s+QWi98OtsV5s/ZB8TT44pm
Y45LRhtgFDK8w0WXEBGpz/pTU3nvvyIeoGuoeu+Hklk/cQ4bIQOR+VVr0JcCOEiVnRrrogiyGHdt
7vHtn21RqQJ9ErYuKsGjcvTm+KxxuCyfDUasSstibOfKRak6L1yetli8liQ/tcU+/pYs2iHF3d7N
CJTLzigg1beYpUwHl/KcGW/YMuLyBoQJ+R68Y7G1uznaM/7QipthTnJlj1puKzmMoU/BKfJsdcca
MFfr6NHpeurhw3eAU35sQ+1mHL3T4trxszGqn9u8WClVIEeULJnhPG6iApMuSGk49iYUA0AaLA0T
SIo5HJcdTzino8oJIF8BCbKnOgZ8tL8veZxf20Pk8mwD1z0tBGSRlFRbCqJztIXy4doa52fJZz2n
ve9Q17N7es46AtqUya9yU0ge1zhGDCrFcUjHAvXpLMW9AeOScJlJYd6iU8OkpQooYW7GnZAvA5sJ
XEmIyyrU1PSLWFnCCY+nYFrKCdn5kG7wP953arUFNQK9fGrORJP9diYg2gqXR1YrmigGx6Vw05oA
q8oIkaLQZJSCwnvXQXl4h28/fKKbY/c09vlpxcOO1v/ZA/F3gBbY5kmtri748uXXTxsbUBOk1Qe7
/t09SXiyVxjOTtMafxR+zaComlLDjKRknzIQcFDH3UYdaRFSpUanS1RvH17hBEMjauxinoAjAArs
8WP4NjgNl87WZcQD4nxjaIR2CZ01ODGSJ+Y7npCAmW0xIMMagJccF1QHA8hD41ppZ/c3ebiD5UVw
89IyucrOdgfKVRt//ISwPZTeRVrrg/nJEuSrz755BqaiBGwx+3eAPp7hQbSKbmjfuu1uK/qQi84v
m4Hnbxlg/JGtG02yDu+TQtDDqKoGtakDf14SkOFOSzSy+Zs83Eo8K1mrMJNSf+DMD2+EJPJpdF6r
DysdCaspPbwD+dWExYLKVQxMTzCa5Tx7OKjdEDKQeOUmPE4uG24ctOBicC/0rmK3trt7EB1S6BQG
Wuc1XjuxYTBVNgIbJFzx//6CPiRZc9z2hEcX4YRqu0eBUtvSrq7GV9YI88RgxHR5Gxa1jYrXaKKN
sDgmL8dK4YkGSLEhMYSGcRz3QKmUOfQQn9oXnIioZGxqeh+jMgSfoa+GNv6Oza7Y4zGMHc1eVNdI
briKWQkUerh+XmnTzH0z4mKEBohLq0bdUIcvh4kLYLxBFoIXtvP5DNk/VCalqERiqYLh8UoRY5nT
9Yyi5XUQkkOSt6sc8Mi67O/GuXIPnhh5VmATZZ6iyF4q/sJBb+NJVjEHzIYbs0VOtKR1El9H6JQ1
EDIyvRa6xZyvXMqgpWMxJOJMzKj8EXB3NN+8i+AE+7hauA2ZYDbN0mLK9dTwogo0olC1OgWMqWfB
MvETMIZsnG1ycCOSbK9eM+d+L+2gOVI2dHVoAuNJ8QaVKud6ydn1TzD0ZxQohR547HTG9a3nXFXl
y5U+AEm0mswDuWSWMbT1ws+PkpifbNV5IEgykoOY/GxCK9uFf4qD2xP/k4YyBctwQWk/A9olHeLI
XbWa3p3GwcMVmVSvk+1+8RYrEIxeyy3JyiYzS4vERNfGsfxsXylreGeaTN6bzBoxel0aDrJAN74G
faqo+tQm0fhdAFgw3am41b1oYnF6gw+aLiBN3+OK3k6KQWhqFObJwtH+MOzbPbyvm2kXKvaPIrJw
vxm8XIjOstkNZ03U5qMxVOgQ/Axt0vqO9XCBcTARfG5v9BCdep162jxaku9TqEtD1lmLVaX+vBWr
DnbSphYOEIA5n2b99Zd3pT1QmrPQDC60P8q3PVhsnjahKLi0neSVQtrC0m9YZMOp752va0KEY7Ld
SOsi2r61DC5qki3PuX90kURHZsZ9JixCFkXK6WqWmNSHnitsMiUfbetIb9GlKlNF3dO3W5QiIbT5
WAW+OJF+BmQc0EO2OkmbWuMB6u3FZVqCwT/j0XiuHM/ErbQMsGgHwqFNGWcnzeuLM0QTwTiRDv47
wT9AuqJKJaX0WJGYRbdl5yfoQnvF1lxiRTW76ZSxpMUxWxuZMMQSPDIuWG87A5yk+F3oo5aHfR0V
tOo9kHHMqegq2tMytRfFScngBDhBgaKCDFoUI4l4SApz7TmUVxFUoh3PDQNrC+r5rIM6YookT9W7
w2vomGIxj/o9bklevRZ6CyhdMTvxVic/pSGNg54nakXna0B370BH/w5cpR9l0rt8sWFPc8ieCBNk
8rPGH44mVScdE8BQ6i7ZwxkGyVMlwCRPVqB++vAhxaFQULuuOqFSVKrtP4Mck0DAiUGhNqeO+FHS
SovaXwvQzL6wjrfb3MR2NPRdfHAf6T1WKxBSX5fdwRxvSvrWT7BjjboCCFz/9apX4XoPvySmvRur
dfgsfXKsXZoE0+y90Xb+LFw1863DDren2y7efdC23uE8o/EZwL5KNlWEtv2cXMdtTl2hjc6vp7gH
0mKjew+79LQw727y4BW3lq6Im3jw2DKpxP9IWxcJvB9sTEt82pm8m0PQaROHfhX/mhspNKKl6sTK
JbOpbkxnWUeT+Q23CMCIdiXycMgLY6kMQBhOUFS4mQMdSRtW4q6D4IReKJPNXwNTtcvo9j5PaZQK
q7uHDIaBifBdYnijbDCZW0E4JHHOQ6o+pAFz/HM1dh5Jd/jVbAc2URwxuDfFpkW0z9ZiL3zgUiqs
PeOzMZOwhP4r0twwG054xZpMf72nolkwG+//xWMYyOc0v9R/mMRcuWIw+/USK7L6qFvqFOQDx5NA
RNUcWF79Os8PqrdQu4rfkhz5LpuWX5yWAbSyJ8lteG83KHJf35e1KFWXD3vFK72DUSjGtiNZsIxY
8RElpVJahDImTyofs6Byjz/29sChw9gWNLOGVeZPR+L8Zzqf6rZwDicGG9k0sHNqm6iv8qriJRYj
7ElWPnISF/zDF2BYBYa05NNImLUQVXC5fUlcogyMWE3Kt5J5+1zKTByOe+32bJFm7W7nEEI3kgsM
7JONEl/G+zvwejHfab4dSV6OgpW9RPGjwNJUSzPraYjhoOu7tsXYLTU7IifwA4QZoTAOE65qxpIj
Bw7T18nrXlmg/tC5F7I2TJ2FpHAB/rQ2lvIiSPYFp08XGc/qKUPIw6HeAf5DmrmbO0FoMiAG7wK7
0lY2NQYPzXfwKk8nocFh7MBmzJGvDgpnVNAY1qmJnoRDIPTefVwRQUu5PgztZR471Bi+Yty1SOIr
VXTqgU6c1cZZfl/vRVxzSUN7mFzRv5Sd1a98/MVMCRNkhHAunlhS3Y82FdYdQjcv0Rp6hZcNGW/1
08jrS7trGjrmuQwSVq3R6m/Ge6d5X+nQjv5b1Q2as3fBfOZZhUDfu2soyQ8wJuDmQ8xIEOUdHgjb
HfN0HKbIBJwm1gUISmaVGDkTvN5lmQ8zevKTJQ4PKqTarFoEtA6O6AAGTdDsHov0KcGSoKgMhLYi
LQ5u0+M1awbsSynspO0osLgtNsGMQL+GCumYWlhlOMw/FAk/XqC7cSChQOX037CnafX0Pd8YQ7h8
A9GN45deVisQLQYsJL3YU65hDMcMOpEJ+qfDjEMW21dLLaL88bsKCVL2swyGPt08eIUnRHsi7a2x
CHe3U/9KbzDRx0kojCmLKZV0SwjJ5/GLumbpNoin6CylqdYc6biIXZVeqXNvPgQTk5K0PRy/YAR7
+CEQ4J2F20TB2uRXwkoUwf+SAR2izVf92dFfn7nsmZd5ryLaslNNC2/sU5e3O79IaJb0ymnvITfg
97IF5osKTIUo1zJe8nKYx7j6RPfgKC+ZL9NM9dqgI/LFNmuQFW02inl07HkxSCHojRSbfu6+m0q6
Ifb7RARCBh0q/QyPHsMUAjAVSPfntPGojBES55pX5SvoPpTZmwRjJeAQ0e0ZtR8aLSm0zEPMWvWD
WdZ2H82ML7CNQ0AfjtOibrPvZR7uYulptkxCHxUOnWCVTT4W8TqrYBxkQ7fWYPZTkHdCcbCD06V2
8iKH2kDXgYdwdtVHh/7qoxKDXs17yeNHuxD/Okw4CFIPQkLdVeNvR54R1ivRhEZR5h5D1QOUJzBA
eP7bNPjR5TevBdCLLLn4mhkbEju1Q6dYLqsDEYnDXhoLoHcOxR7diIMCFGJNKP+e6wIcxD8unLst
wOdu8/LU5w7FjpeogkQ6vJAJfKYCuXXWj5JBEH114gAwI5bxEutc7s+zcJBVsU0yGjiLwR2IeRcv
LataDtgdpkCe5Jhgt7832yHsyGMQH1wdxbRv/8rCqGEZZBK+kFfMH6GaFM8H5qdGydGdqF33i+g1
JT1mJMqiDlKXT9D40P2I1be0WfcHAr2v8AnC4Sbtt5KCgeVomIvegAcX083Jk4IJ2f1kTra1DUrK
bHBrja5Q4YBrC8pABqn/XoiGIemuc7Ygj9bAO0u6G9x2M3e4rwvnqsXW+iv37wZ+FwRD7+4ib2Bm
Q/furuQMttKkmxCU5xAotdbw4nXDEnvcjwsImdJJhOnoi1kM7hhPoK0hJVx2zegSJqO+PO2gxKEm
Udol+pmjF/TwFBWPddVH/l0xzDRtJTGVELV5RZA6/Ft6AOUCMt0Bo+xHKmQBOqW/dJPPqCKEMYgS
oOt008j+S64i2iO+ZCI7hSTGgGUIz1RLz8bqlP2ebd+YNYtUeU6E00GvjXB7sAMFrWHRHnMQ64DL
1C9ZBVfQ0r/sizqjdY+s+vP+GP55DYCfayAHTsy2x60S63gmMkOsd8jIpG/5XRvBcIcjthULvbCC
jChQLNd4iAr37oPXFK+lNJLLni2Xq6TB6hFf4pJdbS2mLJvuM4X03aFVuopB825WeDZ4SvG0O0fH
P1wyxV06/GbkcVgjOLgkqIsSF4XPw1hslozwhB0QzTOe2HZSC+nGVM1YtH/3JIX8jB8nz89L8/zP
WgNIIUBChcON+6U3FujuIvUQWMYht+yEoGbY0Igte2VhBcNa4DOurN/GWyTwth41EiB7pVEWA0bV
NQjt4a9IlQS/iNPxhIS0X0hVC4g+cSekcjR4lfocrR9NBZlgNLM+RcDli9r1m/qyX1cSkarBYyu4
avgkzNgwH8UblfmLYAEmYwWvrK7bsvzc1Acji1uDfKDGKJ0tOf4UEzXJvKR7ht4Yjy3sIRypsRIL
n0kAltuK6xILRSgydlqomXPKJpjCp8Z4yII6vYJc1CKJX2jJpEj5+QUbkDhgLGO+YkvCRk4N+iHU
tgy30QkxDLfEzwmPYFZAo2CO8tMDTSnN4XbdJdFGOjKMffVBRnzrikhzA94cumUMw2pjWtZ0tVv2
YbPkUCdpbSmskl/bdpCB74RcR6Bw4rPPcku2VBZoIDZe3RB/u1zDBhjSCRq17i79GtN0QbdRov3B
8WHvdKwYNDLTLG33+wGAcf8ztX/SzUj6v7dRZlYfVvWbdKMT9ei8uSbC14z+zKSuXFu4dsoHcZwe
IEr1hNCTdqbh4f9jQ9dfxeAQ/1AhE/XTO9yV+Xa8lFoeJOhemL0wcj8hIW9vlgT4xUV/8CBY+L3u
IuROdcFhL1BahVkyrs/4bXNbAocXjjbo0Snp5sFAywUVklZ/1szJl/O/N2TM/ZSt9q1SFww9odf2
Zy0nFjmYW2QmML9hmIparg7HiRcZTay88zgSAJNF5aC6ybsetLHm9CKyc8D8433MC/bd3QtW+ySA
YrGNm+He1cfMXxD5y7Bz67XSaiREV+jo59TSxxmttj3TOV3YxPlToHOLMvLDjwnGJMqDtLjCgUMt
BVzXpMcvs/YNtma3XQuwAuMhbaFx8ssWVi9q7fnt0E2gV3iV98AsV6PogG1ZakN4B/BSA4sRPX9v
9A338ETWhHtGW3+mLEYHZf+mUGco5k1XlMUKv8fNpT+PEIy/Az2khfxocdTZSXyES73PA4QmdFnB
8QACwA4XOeTBBCz6bN+l155NgJSKcqSDbd4RC16nddjHu3xeG7AjTcv7gxf75xtstl12ZB0m/lsk
g6w3o8drsoOPbpgNjPsghKajccnZrOY10hVyEGPlJBJF6RFSSwcuG1z5W5PzcRGtIIavGhdNtqK/
teVmqSFShdyUqL3+eBaXKHUY3XnQiUJAzp8sGpXlXoOsCbDNjtKLTMbsxqSTWpq4dePTY8iUJVxC
XXSykmNryeqpeappqVZGXpsIfjl6KYvp8z1gLblKR5XYuP2qttQvqcgHC6DAFn8v9nch3w4RUhTA
3keOMxVW2wCPxcALoAtI4g0jhdzefmssaRoseRs0CsL66+WHiVXe9GHgJzdVGR+GHdkA3uwu28Qv
/91dwljmstumJCmNFR+2Bcyb02bHa+LXvt2FWREtwa/0lwbKvB0KeIUkcG3uRBbTzis6aOylrDVs
eQ5xWxdwYTr7z4GGEjJEAiuw5MpUyJBocn/yWOXWAPSQe8alGppgruhLsYF2yOj1mvG2mE5BWNsY
yN+IxNUFD2dpnZptfir4C9z68YVI6CdsSRIPdUZpTqwUD8EUpYLckDsTisizD5zmJbfRNmsBpRVW
hxHpauJnlJ3IwSn4+YKY34bWhuJuS6K6DDPiIKRBhRO3FQpqlDbck0yVvggV7Syxv5K2kEC3gaZJ
4i3O0EnbuReUQSfzsJF7Tf/8KyybqKj6ucLfF1PtuBSrOz67xRyg+r4EWWcJkKJnugz4Zlch6A3a
rhX/X0/epBD0v6BBwWJGMcwYB0KbSPCYABYHvJDsQY1LL/fbMRVSO2FbjdkA3uJZY0inCwJJivTL
7wCyOxZdRF0DA/QAKzsiCiuAN5wkXYkLFn5RNkbo53l+b9jiX3RpIjDljP0jHFxcpmenOSmoKSfp
eG6mU5rQ/ipvo/9ioEcTTpuoqKwhpdAmQ6SW8475LZ5BjTfZk3VOARvMAtw36F9TVPfsvmnNf6lc
68zthTlObG37b0Tk9gXuF2IzYuKyDixBozcdUxRyvx1DNgY6HGgeR10ka7tcjmD7QxKw1O6of5dJ
/I3v43UNuzVrGkzOiFGeQ3aW1rC6LHVxQoL7cnAgnvCsg+PprMjhRd0zSdQrbOLjnQ9Bnnh5FLFj
nLFzPezzt1byQIMdJMvpI55dZAl4TpSOZjN8OBV7Kxr3PXFQhP3zWQQgzh8bDZOQZi2SW7RRSk9e
tLhE4gPdGcs1gJhID7yxnUpsTwzq1qgyv9RKJMlg5/90V6DomCqJ7/0bwR0UbvHWo6YAs4FqkRMx
c6+7ejIIj1c5SXO356SoUwFZnzupNBdWJY/aEKlyOwCc9XcarBO5Vzo1NOtpe+F66W0FK0JCY/qS
/akneWr8aJ+nLmhRCRIc+H4InFYlrg24rX7d5CIZqQyNLDody5/gMGvj2vRqEbuoZvKlrlKiog9l
+xbYQLlKxl2XXVXMAsXijrI+GejfaEPbJFo3GNhuacnfkr3mtmy1LNGo8/zqy2hVsRFb3amk/agz
sxEFNi0M4nXyKPAjRqOwwSVmqbXezzaqdzURX4K9SnE2wACLaXFNeIy3Gni4ej7cawDew77iFoFY
b3NM7qIh8SvLKnvntzQsXwGiR2L3KUrWdJLcC2DVWBx/cL4bJ0bl2zqPQ59CoKS70PSO51DuChwp
rZMGIuStschXYfSYmtBc8rIqlF3cTzB6Ag+TgLhOr5Ic4k+J2cAA8MFBoL+Xnhf7nh3bv5WdKD4R
DMbTo0Ih/ZtOPNhtaMisSjg8T/P7E0AdoV+VKCaI6TJGArGXCryzfgBUvaju0/8EICkxl+Jj8RBb
BYkCnLVMktrAUHblavMZkhdGYvC04Ihvdc4m6on47dyWEsbFYb22jizUAB9NlcP2SKuykKVepmtZ
829KXarMWa7C+NdmWfsFdtxJvRMjHgQRXZk7XkNgZ/aQC63Ls4zTq2UL3StMmcqZVGOu2AHw+jY2
+L/hjRK/H++4QUJVc8Z+7CckUvRgCj2URbRFnK66m/Q7dJr3fDTm/2sY1Bs9Us8yg8wHcXY8D5nU
LCNRtrWlE4J9OEAfe9HbzzTdyJRbYduSHpiskoQlbvI5kFUQpP4p6Nl38BhPAVU+v7YWSJkzZq9t
4atmw8afPXKJppYEbt2eJILTa/jek0G4D9etzqHDchf+FJdONr7YzXdactakbNzYK5w2w2VjdqbW
qUyo0bB5af5G37CSnHdPf5MH9205Cm/eXuFUs74OgjoGm726bSNPECSKtP+g21K/7HXRjb9IsoDy
GD+xhv5jgFmGJvvn/jK6xr/Xh7+VF12Hn+3u8vAyljaPRUrV23pduuK+KtkyKqErlj2XKNDGn6cb
WEFHAi6w5BSlMSUCkgcadHJLhpTx4yIX0lS46WUL4QOzn+5TRbMJOldgp/sT9Q1UfYE4Sm6GkdLs
QQWHU4J3Dcv9EsUv3Y3U5MHIePI/KOJPegCFQjVyT0bbKciCr1tSrKXdQHBGroQPaDfoI4QRxO2A
3O+RWzPHeofwpORDjVBlt+EFpzspdChtGgqSNX1/TPJ8f59btmNXVNsHwKXT+k/K32k12NJL4Uuy
rm4wyMxxQlFfJ1J9GnEECjt953CMyIXTjpL0xqnFekKTW6iMb4J1U1qzOD3rPPUfc58gsUQoE5Uw
j1pn9fSV2/6S8hidzi1mxCCV2rfV4U1zP504vgqTgSL+b3YJKzMNkAbY5Mr4ZWt/tsG8fGFHXCxh
VRy4pL4/hgKv7KD+YQi06VD75hhBme4L3bv9BBy5kr172uNvSviyj2gbNHYlM1pj6VulWE45eIxY
JSFa03ML5533B9nx/8JcFcMHjXqx53/LCGIjt0TIawH1n+BA1hbbARNmbDZlOnBMi9p95ekAE9Yf
48n/JanL2cg4wkXvhdoy+SKIW+1bxc8tV9Z99AdJSogVxD4Aqt3DgEeIhA8UUgWqfssTJ7io9niQ
goV8zjtpdLHd1/WEGdFj3GQeWUpmzll7bCuTCbM55gO3pDq4TKJRKNj7kFm+39G4DyZR0WNc8dhn
xWxrJ+rMHZ1vh4SnKaEZLT0Vpa77TBSdbpayKsZw/5Zos67jpnspJYNF5Z0cgdAESQ63zwOlY8dc
qBW094yPojqNyicf8MR+LAtdpOadxjJXldeTtDptPX73p/3JG7QB+peQ6HRSpTVntNyZIpz7uIDj
/L8Zp+hHDm2QcWGtXqnAfRl5nufKeWT1O5AjojAz+awy0QkYDghTknk2vDQo9tdiCD6SDG+S4zxZ
h03x5092pDnNJhdwxVs3R+VPOAYbEH2rEYeLoVEze6avaZs1nBkR2jcce1mPcKFijesvrsaKhmjW
NrkngOmviSyIRN0eWrEBCemxo2ztBnYiD1YwUynhFRNioVrRLA/xQzW+5Hp2ZwWeBwEAPy1sLIo9
wKrWTY5x0yNVrmkNQ74w9CFUY/YALlysn47rSxGeC3A4MxFImIb6QOOVHuxgWDF9qQQzVVvesfp6
pAE2vwD7wu+liXXIA4YG5IJtq96/mRMKQPe2l/KeHdJb0pY2dRcBhMjyy/I8/eGVznb9S6KB7xa/
XS4MJtvYN2+IVeUuwMXFZSWquCSDq9rb5ijwZXIu1AW/uYa9BdWT7QRBfwhv0ydKPd3EuN81Hm/T
fN4nT0qo7u8F0Stxu4l5xZWq7aZrD2C2NVcM80VKvPpT+qt9JUFoVAIivVqsB5YnJS4UbHiI/c6Z
7Ec68LMHcAClg4Dn7t2EZRVv9qoMOFfBel4zgyJWojNpMDbE07v1W+4sxNvRGPDR32bNm5l46gt4
7TW+3cMASFsuM1SZRbuefcPY8jN4t1QjIBNWAmxsxpYeFc6i40BKjuc5zGwvTTpO59qR9cNOE31T
+xhzNiTCiYCYFqJdEx/0JjlQXW1naXI6xA11mCOP9/vacPIaBb7WbHzrG93An8FvZMVR3TTVZiHK
pA3d+a2GbGNxyz3AVw01iso8n6B1YGgeRQOyVFLafNNg+cE2/Hunlctl2lUGYLUjqP1mIiKwqppc
vSFw9/iz6TXcpLkFtBRj0/lLliHql6CWQJqspcXUtM5nhMeXMyYanunMYrggB5/ObuKLaN6qRCTq
AaNTdz0LKuWyOyds63axx9RuG5c9IIZbAHe8GJXRqTZUk/r/DWjrJKgGetewyvOFI/f+BM3TlHTN
u5//qraPE7eF7owGwOipRCH/3jGyuMLoYkcq2P+tKvaZv12rrmIYdIJj/stLhWDYmNcBJItQ1GZ2
lY7HAR7Pbtl5+81FI4watw6qCgqfwdCGyUvAfkjpTQ8Y1TEXkEY26Qyfum5Q5LkqZqetH63LuBnX
icPA/gRrp1tQCoekKYqE5W8z5A0507D5Nj1GahiQf7YvO8wnhEb/v7gfoFPEYSOuZ1htNPXEbgLx
QDYel1cl2KBC+it9rQi/tjVehvN+ZxrYeG+UKJDfy+VDN2PZVfTZfQACS0YMF8ow0Wl70f38MjwD
SRJ0IsaQYxwkYoxcztd9Fium0JXRxJMx27muYVD0ew57px1SiPrsZ+hjklarwy4Ec4zPEwRnDp1v
VjMYTM855MY+hDINAfbdod9Z9U4PGJLq9igvR50rPyU/YgGtUtzDn26it3kQBdlPKmpIuzp+sDfe
FiDV4WBccrKPYeorXmmAeHFWnFO/Ut0ktFw7RjcArFV/jdApOb+CXRPXNxzqOnmiSFepYP1jfHVc
EN2DAJKCiXl7/leBmK99mBUGnV4L12dpe7yeIBH5chb8eT2sZmn5q2KOAu0wkNCbcYDEmoxBocoH
MEEjXNnAkJZ1z7psiCL6lJVjcbSYCxzHSB6B6ybjgU1Tz3QXaN5peJviEpGRnlbG604NwhbPZMAz
JYT47dvWIc+5X1duhJRK9/PWsLWmR2iBqj8pcVcn6INts9+Idv1Pu00zC0WrJNEWpDsZq2ql3a36
SJBv840WNU10wKd5Y9xvwkchpNSqGmSJ4hAHM/CTT+apcC90n1nPmAif/EBUufPdwURKxtb4ZmA3
Rw6tjDTh3z4rCvzqqUM4uq/uTgBficlLuhIpLply0MVwnJUGC4qZk+39WVPrSa7wyPfkpIT1awLX
DvNtrF833TEDN8LNR8Ms+9s4QkIMdMZvoJg0ExwBEyt6EQiMVxPwJIS80m1c0sOryDA3ej3CxXKf
+NkD+wzRVMcVj9R3uOha0eo0OnxfOmX3Kg4Gw8wgyFCHdp9XAXpPluRCMk/wa6lud36+k1JjORqB
cGr0TZEzRL2I0+dEt0cB75KuJ/1aXdCxjKchq6uERzrj8NMN1eGaqjN3loqgLFxwZTNQMhE8uff1
qfBZloeUe5WcbNUL6Nrn6XqsM8y6cxXk3vsgn1sy1+jxZy+ZCrUN+CEmiq1eYPe3dA/7wOxd9DKp
vno9T7f7K9U6ZqJ+5axh9HauAypZtxjZHrKRA/pqFLkYSW6V0HfeeqfWFCfqN+ij96/O2lnR38v9
GEXX37rAcPEt3Af01+1SSLIbVobG1k/kY/ALEngB6GFNzNgsGzOCxs6p/PqXWDXAWS9CHfkTWRRq
IMj1uf941CmJ+KARjn5pLx9J+2BionbtysgP8393uwoluInW9x6FEZx0LHaGnPw8JTeEalVToihT
5z8PXxWm5dfv8NrbO6jB1vetG0aqb5m24S0cVZUgFORTY5BfgpZNam120+gwx3D3r+IWgRya3U/w
KHVFfGRCwTM3uozYCHiAVbiPi0uTN7e/GXPAV/TExTkeS6/9onmG64g9IRSMZaFNWjGDdvl4Vt26
KlsQ04Ebaz+5Dav3qRheZvY1+bV2sgSYrw25XDXWVMvghkmu1uMIpg9j6O8KXW/VG2XQWcAXUREU
WhMqhpy4Bneq2tb3YxMnTgmUNPUKa2OPFl1t9iLKQ0nR0zs8JLlUs51eeRUfuJ2y1/j3uLuTq6P3
pb/p4iVg8yVnG8I5c+P97+zDSF4LYpkdwzhWfZD64LdTy9m1uiddZmLly7KXsh2MGj+pIjxij4Pb
qEkYwqz/ROXmIDiMTTC0iXJTR43n00Hf4giDul8u17XpkeryRFLajKaRAjjU3RPiHwm2AWGPsfOR
kP/+isCaBY7pGdcwS31J64u1Gelc4/ZFPOkB7qCRoeOVIxBBx4hCrMjTmaCMipTK1uXmNN4IyYMe
4yY3YFQidxWycIRQlNabMlw+vsE9O+wQGWwah2KYBIME2kCGrQH1TkaQuu6oaeI9bf85DJ8+UIxj
hXFnXTpRgqXijUUWo8Siqmc+JBwCTAD7JF1m27/6IhfsipjLFa82E80eDL6tGPYmwDVIZpzCectq
njPidTiWyqjXvZhZ1zfgYI7riadlVfusqsttGIE+2+f5N5JiV8u68y1pSD42tHA/v61FK1nNbKZY
C4k5uGZAnjazyCc8mSXkFlBSbDF/vEpIusna7YLUdWFb4ifcgqAtGKM2A/nYb78ex3WRMO1WEe+M
8+fNcCYXwappDJYZ2f4VGm/dXFm4hSIFe+6efa4zzXoGjPGwa71NC/v094EgOtDrreskcl+cLu0I
Q2DujJv7PekU9UBv8B45cyRY2odJ8otXx+OyFXZsKyXr5ypNTbcBTlrvfR77x9a0XqeHAOGFzVBM
p7CEtz1JdL4QmLR7o2F16hdb32Odhlb90Xd1fU4hOB4vGfPz0CUdpTCVvYMPTkVjSE9ieRJfkXoN
6NVBsdUApuxNy5+QJwDGfJFM44wACxzcZf/FnbA00j/tlzCLfmLNjiy2DPu1Q/rf9pk+tPAVFQFh
2u2UfD2Ep1Uq2r/lDUPunaOsVescMsF5RRixQauV9e8pgOiC9MOyWsULBbKTlfjCfncWH4v3qZCw
qqd74XonQ4qhelgHBGPGhD96MIiYejkDGR/v5ehyzl5T4A5jtICiv8hUGT0lIl3hesZWAOkSzkYN
d5uGpc/gqtbj8CgcKppAGxX8L0kucVvxNVQSO7nopsz5RQUTdI8gOFJQMuJ+g4S+j03QvCGMa+RI
Rp3t94AmInjaGDHqc0XeCHdAkrbxuvgbnnfmcm1RG2jHC0ntHKBk5VTjORG0SDP+1EFoiwYmv0st
B9B0uQksySXapCv+xEtHFIHDxsfS4pBt9PpL1n6aDomgse3Amk0LlXdKhq4AohKZ7f3EFuL/IXAt
JtfvnT1zL3v6TQk3dxNt2MjvX35XoukAGq6N718aepHVSxHrQMJU+V36sG7xGT3085ks4MMyi2fV
6s3AkOzSgl581FyY6hxOdSGE/ZB5SItFntQESsR2iBea9tn1CTwqobZUb7OojEMRGtwmg2Pt5wpK
gKEBh+pigyXq7Yu139FWjuKGC3wuPjIZFjTE1eYjuzuD1I47yci2ZxnWRwbXP5EAGUarrj1w0I2X
+yrqErXYoSmpFy7HxrOIbuTCBCeqyQAOzWXOEdIh8AgiW3PzsO4zZtVm74KiSZXnwBD6vRGZO2XV
FgDs+Nk9RSZNvbPa0WK8lQcoYV9jzNtt+NH95UJBl2ZD0Y8ihyMCT+LGeVnxYAgb1IzugKZ3gsLM
/8UHpVJCwK0VVQsmEv+gUFE2ZjJVi0+zJoTuJdZ9XvS7DOJF6tyuVlwuBL5HBiah09sg/Th0o8TU
DUBUu53BzcLZh8i2dlxc01TnU2tGSILyHjJhujjNfJB+r4Cee4cuw60M6YbZfdSvb7sX6m+UFnZl
YKCYxofSby4ExUwCd8j5cDHRLLwehhFddhn7elmiBGb8htK1xzlxLSIBDuAByw9oFutK2j6JBBAz
+IZ/gf0I0OdKErLEyMQTjFvl1Cl593F++rzuOdZ9lXmVM9dsy7/22FMaCCIYW48nCRfrndNqn2iI
4PfdQw16pZVsvJ16WiNmP5qYQiIm4NyUXgmWTrkwwDmMP48O6FLfnYCkIC08ecgsneSrVwE9ThMl
wJM+qoCoaG+nm8WQD/VC9GtjhwNauaNep0FBqzUvPOq2N8OJ+56xvek1dT6CyXj5+EaoxAr7e+88
Te4npMbRizKbUpehuhGH9HkhYf6dFJyb5VuvR6Km44FAhtBCq0fM03fjkibGZB/F3jSQci4kSmHQ
UMIqmrlt6SdsSYu/1e+SCM4zKh5Kkq1e4WSyUdJEbFJvJLEJ3Lqqk8qcMlYD2BZrj0G7dNRlA5zf
2pvsfR2s7A2tEo+2jjJESeOxP5a2Ke4ytfGDq3GMoL7jx9xvsaW4ugm9K6cPwNHza1lrxLIF4Rh6
WEAQQRBwr6UEqH/HxWsJsl8pnGl1BD7gAErK5o3MfQGlxvXb2NCjxIzb1sMzNzL8a28jZ+Oc6cB9
BSgdUCZjJW+7TkEPrYIxc+q/PIp9Ia/hKIK1826SpYQV13BhGpzQkUKrCURBkPHDsrUMTMcuC0u3
n2dJ3m3Xl5Aw5WavR88MiueR3m6M4Zv/atoAPPIgzjX+Xy1+iqAt2KI466U7bqidO6+FL0FN8rpa
NXG8iYd9On7YACS+f3jzXMtrdwkNvWje7Be78YEgv9faSnToMiDSV8JiGOcktoXRdVklpnPXALJC
lcSLHLP/HN/C8JMw81u3zXoIIXaCxosBZTNds1u6dPyzq27ZZGtgxSp2qDZPMauTFLnZdFfTjgm6
XH7QjYUmDcCCPpiWRu4Rnmk/+/QFlFWZcP+AHXfN+OJYpzEFJsrZun5IG2oQJu/38X8uR7GSTqnG
1lUt56iWh8+SUszyBg3f3zDqAePiieyI82RlTwqY4InT0wzAAX4A4+KwljLE8vRFIlbGy0ZhWHWs
NPh3CHN7dBcfp4DBp2MIPmzQJpZvpuZqnGi4JmPF9sk+tAZb8ZXEyczvHb1OQu4P30TLfaxMGxWA
iMz8yMQ+DLz7lzgOZoyO6MBD9HK2x8is35X88mFeof7j7iBBgJtfg7lF0WzSwbHczm/2Hyhl31pu
bmCosaW0NColxGmSLxORJ38l1uwyBkwIkF9VT9iM7mbSLW02k+VyPvgm/rILMRYtV3fCbaGerfV+
bbUUIi08bpUsFVLsypkJj19YChkfykOxXAqd8S3yEey4E9SgwnOwJX9prURHXX6HsG8XeK3xc8QZ
K532QNqJ7NBBwJokaI+yr3SBLVaJkLAZxf2zpcRoMMN9uAeeIOUJddj9ZvBVcZkJH+F6wEtfJLCz
l/IGZB8Yg3cCZD0K0vPqY4lxx+gD2SoXgkTdvR9byEbXCzh8WXmhtgD++lWleFsMsLcr9NPzpiIn
HggF59leHPJgljH9xHHZUF4KLUGDoMScvQUOabzoP0Knv3rsWVOJMNttHOFsGkmSthId08Bkr35q
05TIhj+NLakDSQjgaYRfCnOOOCea3YR7TCIE7nyVXlFVjo1EmE+c1kikC6XF/+dkws3biq61Ox9h
y771x/mW19gszz5lvCI4m150UwXspBrDGRdBf5sAUcci5y9244uA8eY4Gh/xbsQqUpao/gW5RVJw
jGCp/4raNWfiM8vUdgNS9VtLVAzK/fIzlxusnCQ/SMNV4CjtosdzDXxf1WdgqhU6kvbYKJjT/cDp
AHKdSByGXv151Fb3I8aFhRipywRLcnhoiYj+cgIpKNYTPx+YNGn7204TzQ++dtQwuyD74Fbgl5h9
a7Lgm4YNQ0vR63NPczLI8T5fwqk/m5w71nPK8uypmRztjtHvLLtevrCpUssE4BgRLck/QabKn/lk
nT2QWeH7TqMh0lIVLNLtcWKQ5/lDmvUo6IDu8zNoKUdRpeWu9/fpWsgln/tzGFFMtgvcHyXkQNnG
X341RnviyEcPK7+f1OjzvYtRMwBT30lYkObAC6J1mh+r1UFS626KJVA5EX7Abs5hnqy1uPDxlRNt
ChkLPIBlwv7C/G3rHXU8A1ddEk9W1pM8o0n4KO6RJCbgBAIFCvhm8iM3WMdEyA1kbRPIgAMZrVfl
vCC1LZfQasqUvMTvQFuMKwsweNw5wEWHvZsIKC6ABWDVihCiYzJ6/3ymh4mhtzt3a5Z4jGUwMZTV
ahCVPDjwBPzeWuzIt67f1QbaaoN7YdBd4Qn329gbtgM53T/BuA2jxPedSXYQdyrxjuRFi/XtXCiX
IAEOTT/vbLpr8QU4OxUj0A9BUYNeG0nZZKjKgLqN+ZZ8/X0czmr7XsOaheMALsdcHu4oe5fgzs6p
uCHO1vZCuCdUhO2udxzG/55JZaVy0Tdl/6HBlYmUx27Q8oHCLYRKpQsXDcR7gL4p4LRYH5qk4kPh
argMZF6lJQil0R02wvb4Lup2VkMd87BghwC0MwdX7bZqqyLJDBmktPCKXwBIIvDshSbq+V/OQ5+E
vZiSZggwJYgk3OPUeluhkUNZ7VCTadhVHumb7fHbBGAspq4yXb01FlJYL6HzkBPSZlcpJ/n2ej7L
e36GWw5GsP4CYCjsc1Mhup2ellbQeMvmpccffjUzF2SinYqTdQl8be3y4oVmPsdpQGa9+gehLCRX
eoa4A/IMzRSajretqp+nuXE1xCvzcxyEAhGL7ZSH2GmDvQC/RkZdWL16Lf/oUkR1sgQjoGSSctOl
X2pevQwD85YTKZIlJKut/IpDIAKaFQvoGYklvUAOUEK5J6FkwC9LUCfdudh9k7IGsnz2Kh2Pz7Cr
0mHJ69KrpvujzNi8ax37EjcmjPKVJ0Wv1y8saQ/qfmEZOYQPXOcrTaX5ekcXJ+/dfJsXB1bwIsgi
SuyuOIQgBJabJYHkdnG1KYbJJvnDqtdUi0rN2dD8R6Se52P1KSGKCj1LChHs94eO0pL+8lro52Kz
mr9zuYPVv49R/hM0Pu2qkA/5O+6nD96ncrSCVgwzK6zpFSW29oqDTvtk7vEkjpBJV0sOTIZ4b8+4
vXYuML9qpnRqC9Y/5CF3YncuW3wDCPQdD0GHDJExVBEwREsRxzvyl+hKcNvknZHxfj5sFq4FpbGb
HDk5tbd5wWJHpAF/IED86JkiCRlwvmvvgepmQqFlczpRmRt5D6NqBXK9L7G5DHb3QlY8ykAaPvrR
kYxGCnEuCPlxX1UvFgLbMcF3hwixrQzeV/xrGHtR2UnoZXOeQG5rEkCtvGd/7sKxdoqXvkxG5eGS
C9u7bWpgacFBT0VtAdzpCA2vIsIo/gAiirESQy18cCI8wHZSEJFOPGPiTytXED22wmWALxMf5+E6
Z+xl/zrNQJjR/f7j+0t/g2MFx3X1VTzqtx4QrMDgecx9X6f0FQIA4RbwkF+7wabQqT9/F8kpxYrS
IW10Ov40nBDSB/xBs51WP+T3VkcziTzkygsLiGhLWZSaF19LmtbxgefR1MpzFmOEyx7F9OvOZfoU
rMaYIiAqjIXd/NoRyWRKldTu2IYirKyZWOGB5+mF0dGZYGnqwmUo8kn6m3WfoZNuTwfTXOKgLblM
zDmuQgNAw72L7K2OCiuhwhdxHzcjzCmprfbCU5rVlOpklPyD8ALbF2f2OdaJ83Dfiyq9b4faRSe1
qWO0ZSvTJiw+vfXxCuoCskHethEIXpy9bd3XIsL4kgcdhLGVN9Xk1ZY2+hxXWFndATPxrkLITzHP
vYCX4M1EcdHBZlzPO9PyxdN4PHxmt/V8C2Uxf4rG+/sMvLRE+QGE4jGeiBYr7ECcGxcTbVd6YOEh
288Ai6D1EPv9Y16qcqweY3ECKbmDowYYs2gYW0+tTnKLTJ9wpzEaLcCvbPm3QnxwP+0GUM0GRyYa
OeamvQ1FLuMds/jkCZsP8LIpmvBbAFjeRj36QrIU3kBRxQtZplFmjqpO15alWPhmtjuVDshBpsKy
bIkaNJGFE0DqE1XsH/sbgRCHc/URkwiTYSwcQGOTtxzdp8tZzaN4EQk1/G511NJXN2T0XCd5zUJ4
9x/ewaWA+A0gQ+oKYs0WF1auPz8Guldd+A6z3SjII9sqoiJSVEXXMihHkwkX+ydDfCr1OfWew/yr
B2MFEULngQ2DyKHjH/cT2DilN6PkR6358AIZUZldlSzDCAiTlb7Bt+VZs4kHHlc/hcrqm4p9Y7VM
rwLNMLBLyLbvHikpp1QERIeGK9ULfQxj6wrgKPR+zt72O6w1hKFSUSpLAKt6MDXaFYRQWLLIQsJP
6+oMG5OzuA3KrqZx1D6O0xNWTkR/7+ll//27UV6jwgenxfj64qUM1xy5QB5PUaEsDzXJX8iDWU/W
q+ac+MuXzKTUM23WkHglVfN9SO1N5O5iCXX/IspfEl25F+8bobnDar6l3hZhWuuXCv11+5HPAF3D
zrqg83ruD6vNXmimTJd4yKRPKp+Os+CJCRWKtzj+iThhnXF1pSqTRZWiU5SptgNvf/Lh/TyoGxAq
ffXoQ9V5AoRDIxBdCBDdGeW6ASAXN38Ra0HC4GCz4tTuSDqxOA3TiK+GF4F9Oxg97v5E1KzQAP9S
aPkFqfHRG/us48ZbqDKQcHYU/L+73fyN2SUpZxuDQ7fpxBuUoey8kbzi/R/DUi/LrFFOfSDoUT3l
6nLoalA2O8V5ShtxHjUbCc2cngiAmJWhxRG4PHZEYXjOqbYRUvegXfYqsHJegzO5diZettp1VFHX
BF8IAOs4yO3nFAoYfkzCb7KgyzKFN/4u87vd7V0zmgT9bIo+grQwQCW5mb7EJbaTtXYTaQW5dYRF
YmXpfsxofu9ItSo8idwZECn1nlWnMPhrHA/Xyod16WOjXHUnfnAxTwHbpJJsoI0yS9z0zmfXYSWg
gdKskmroFp4queRcd+pd3QVD4HNK4jZYlWOV/zG8g7geYNUaShVfyi6GdNlrFbWLC1PTsEnLwf0R
qCBIsUFVVLwQtEAuNNe/90HQmRFIDBybNK4yjfgyI236Xf8Sz6DGKDs4nxofpS/IgkxtwPQz6EWR
9YfHZs3Fzpw7iWJFSeNz0830ABA7RCvs6UseCfuULKxFvxEL8ZdwwixFRA967B15mgmpOCaOEQKX
lkqTJ7PNV6M1z46J/lDCjhcZWe0WEKLBkK7nQHctODUHRIgUJ6PDTijpfmG1rEKCVnNSEI1YBXP9
IvWq3hfBjDd0MvSC8Ld7RMa4N6PrJflj5rO18/c5jvJKMveb/B/n/kbnHRihMv6vSVpvkqICe3hS
qJVo2LK02xVJ5c8oUfQAi6N+ojVJXFye+uhKMYAaZBFRwJ/DZiLLd2S0M4JRFXQL19PsbmQ88CCI
GCqaixm8jY2kzL5WyiBHWU4FQEpVquOMcM+KUw9argcburqjqmG9yYdJ3mU4i9J/qV05Xs6mEV+Q
xgFhIm9CevFyNKFMqY1M3QHhC2OK7pwrHuw0itq9Aw4nIOatEAFA5Hl46K6X5g5dVV15LfyGVndd
csxqgqKZ4jP0ECG6f3z6H2d1Jctn1gGWIqtqSLOuOlZTGVVkllEjgmh9VDD5Rc7G+1zR53SLuikG
B0j0CBrQOiImABw+y74NBipl5HJArpp12oux7f+mhpiad+v6cO5Ks5uwgJuo7gKf/c3T8D9x5ZLX
JfF9iiV4MLiOMP+V4S2TbN7JJX2R9ghLGYclp1LHnJ7eFTpLgFml8fOD0SgSDpD1mIW9zh/t91jZ
x1VQQjvMrBpAcQlIyCoEiZBpMhLRZONjmzYsrgHDDk6oDqwqYqiQVXcXZSvxDB/3l0YDFJWhWgp/
TrdULH07OEAQ9M2L1hvR8Ygtx01QO4iKGb6AQS+AwgT40RAjwF7JjOE9XhPmKyrCz04k8NsJSwZb
GhtNZGCkt3XybDrPke4fT69/2pggPA4ZXPcPLSlOYxMwlTN3J851rkEVVm0x2cwZCCqvb59FYTLw
5TalPOYISLwv3crJ28mDH1b7dW4Fo1AFo4vdO3mesPU+FFkOD2D8Nlu1G0gQ3KQpmnR8QNurSxxB
QITaR4yyCqjXPworTmrschq2SQUJQc69lVY2VDWcahPUkQjg+F6swPQDDxjzEv6SvrOs2JevDh/L
nRlRQJr0EfXW92mztTYgp1UpXdOfKV7kWTdESenSzzquE9EypH8QzVVvU0nSAsKalfzTt4DqyU5K
tCowMM6hXSFHTuUuN+fghN2TzJwGw+pnmt5Q7zh/m/wYNOzjk8Yozq+ndGvM9KCf4czEtam9GZ64
zem57BK6qFEh/D7+p8wxUg5ch4/H5aJbDVBkI5vdO/7EWKvkVrouhJyikUs4BYpsqgziqRKk30v9
64SCv8KF1wbjzCL7djrTMP9ceoMQ42Y3tAs1QGQ2EKtz1by0JXINgAfACL8ithTWH5YNvtW4egSK
nSzN38Y5Y/Z4OfmuU+3QjntYphSIyf+pxDu3Rg3qCIuaiCu8Jkod4tYNwoQqDmbRy2rrTmY/1wjx
LgKY4OCqX2sJeGgkLO9iDVKk1irSW9bzN63N8QDkx6IwpacKiyB/a/7ZnkdV6vEXnR+m7mReaEW3
QJ8AsViAuhjCX5lfmx2Edwy9OQ+eaUGt5H13vd9oTJgWwOgnekfeO4IU19gduUkDBLjg0ZyrYIWa
411xfAzklLMVP5GmkMgQzDwjzkKLYDc0Rgz1ehx03j9HadEnVIMcapBnp9VyLa+DTK7Mm2GxPYSZ
dEN8NRKFG94VyM9wfiClmVZqJzZMlIA74FEhHlH2UwufnBvpMFxC6PNDIf+VQGigDYyAx+xVSI9H
bS7q3/0XcU7aViaj3xyxl0TWzORtmoFckgs4rMCzieg4gPie5CUXetmpgcT9UhLkQ27GVVq5/8dS
1c3IBfgOLhEE3Mj5C8JBA7EWQ0J/2XFTcdmsGNXCwzkfEcVNB1Z5fOtUYikoGj4sFHKQBZ1J6nux
VvC4WK2s5F67pFSqcGRX3lhc+zXzTl0aKePT7ZSJIDr0cZrxoMvq96pKyljtIeOb+Nvs9IzQJ5ZJ
VsWCtXw8U0wS2/Lv5ls8MXb8uNhPWh4E+/xkSxHRCuo5GgigwBE1FamtBDwD97XmL4rCz0h5lbXl
B5DcAuNsBMjQVyL4drsBGWrZlAJOBf+V0JhZ0RfEFSG2lgupeB0kkfhOCfkVfJpQs+JS27gz4ww5
hBvSc+KWoibtjdoZsnH9fVWWFuwPaYGeqvyj+lkIHn9TrWViR1b8ycMoMH05URQIYWFG6doY2qrl
57MpW6cRx97I7qXXZBO2sLFlWv2KHJf7HHEP4SzSju/AjouWafcdF47Az3x1AzEZtQ6A2nm8zrxv
WR59zxdtH3HK/2fAJ/DV3wYW4/vux7xM9f/lI5kb4JPti4USR0V5KueCGpxymDEmVn31TU3wjWBL
75vqJqQBNKdlAB/8/gdURmYdTID7hiXjGaEKhF6gjBZHlOLqktmJgzE0JjOS/NkmNzFWtRvmJm3o
ct9xfqHal6kWjuOG+FqqF6kfe1jZP8Gaxgl+P7IKL3UafgHLSGHDSbmBAc28+drEIfnd6uliAJ7E
IEjS/pVMU0GgjSki7vihpr8EUeGYMOBPOgqVqr8yDMZ9GZYeflLcDN6IuRjK6hM2wdKs6Mq4G9mY
BEqOT1eREqu7e2L9QNJENASkHN5MVvzwLpsBv82bQaEXvYR7F7T/yOVmUbZmjElhA7z1fywgsLWe
S8qL6jcuEPIQpCYTHACZ34Jv9A1t+BxZLpDnxi0hc9IcWmztfJGPqppBqRBXz0UQE32kXGhxNFCo
tTwQAbNTG4WGw4nxSFBs9XsOBHUK/KoKRZncco1/TJDUDpymaenCcYb8df/OUQzH9KtwuhVihROx
5DyjeIST2xGEqANqFwrP0QcC/RlzuXTgt27/2XRh9SExM+uIE8GBK3UNRtH7sWSFUYdxa5KHH61W
hG8bbqPlkZS3omt07sq4+plbWc03Z1QWT4/Ry1zqqiw+9ZGn3wBWQgYntMHUnQeU//U9jVAMX4RS
uD9vNp+O8BPRkoRJVK2HsUPKmFkWOW3vQKs4EXf9mNXxdJShNASceJ68gsOkeK3cQrda5hnoF9vh
jQuc+REFFIblx5xPAzGXFPhH3+Pi+yokEqiCpromYnyEjVgdDWTeLmIDT7rXJXoniQRgDoj3idzo
unbgLqp1Dt5Xuup2f8d7UzzfaKkjo41zF5UpOdqbqHgcSXzfpj4miaw+HmJA50ERWLicCUv0BHyS
QrfJvqrcupcw7XuvkT8AaSADmbdU96EFP5DfetQ6qn8pwNMLPrGOL7yZWuyQWHaPP1TlwuPj+u5L
Lv2mycLysthV2dAK9y5FMkjQdzrY85r6XF54VirTWnS2LexADSUkRmZI1skqyvuwxPI9Bdk8nwqf
XgYcL1ytOWB5fc4WOEQFbeFYgtF8ZfU9tJrT6fKacKiRx5dTj/ouH8xVf0LMqwVQv7tR+8IBGKbc
YJP70OfM9k0zvUpiXB7rvJGRkZAC2OpimU9JAEW0tMYgIfzWQpAL8WP2Q0/w1akjcwDd9qyEqH4A
AvjmcckHtNQ6AKnm2DpdQBYbPqh1jvC912MqulMz+Q0KHHf1is+QDFuL8cOZl41iK3g1H8bzmDUX
uUAQGmti8BYNt+DitoYzoYCnEuqQFh1L6vn9/tKp9PB5MspdVFwWi6NBmgsaQA6xAat9/lBOPe0N
MYtbv6B6EnBIw5KNVV1Pr0ELlTFUicTxejvM8vhZL1aC9L/ZK+zyQdjyUmjeV6HT2NToyfHisW8V
26aMtePd3vE6kv3U19w5Ab9ttrs44UwtAk5x+ajpwIKfGG1sy9vyyv3jKHdn77NYhppsyyvnSTgH
N1NW8RMmuCQrrRN1SnVrMzj98oxSVTVLX1cq6UtiY3XVjGINpdsmUHrILB+bVsUOW/E184Ldz5VW
EWi8fRkT4hzudJeoYG3O/5PEpmqH7HrCVzK0UrCxrWXWExWjXk/zP2spOJiqRy/dSuB+A87Xpo1Z
BL7iRocGv3kEASJW9uLb2zQIOUzhQHFBKOnTrYRTKVI/1LqqNi/8dtxXY/d/MU4R7iOYlQaj/LfR
jiBQtLK+fGPmOM1Vs+cM/WyjwpvwbMAZ9qYpdYzyyX+LX2PK6G9hn3Muw0sSV6i3m1/nOEe/RKBT
94YfRhtKPMG+BWi/tJp4OtvaMFcvSgaIGVAuztvMzMVCUDhu5tBJ73Y9L5Y2sBszP7bkHuuzOmv+
ahjAuPhwT+IK96CniHDVM0z64Z+Y9Gi7IRSLpMC/lPj8VKKQTwVYrggeMUKfRWSSuZ2qouu/wt8F
px1DS2axBXKrqsQVGOaRm24robE7uhRb0LGkcEP9gh7DDe2DybhPCNwgKeE/+OrRW7so2j7ZR5m3
5AED730K7oCNeKDi4Htq18gfWiPyAGwuoWD5ZRwFMvLfSPLZRBCXXnTaDopv6FkK/lUAKtbdAL5J
dHYNS2QMRwaOxJ8f4cj/uRUdj5F8fMGIgLJGfqXJxEJcETGeCTkN8JpYHl9OWxGx2ls3N05KXBVg
WaACxOgZ6el2/DQw9uO1krKeDqKBiy8s3l0SYZiDEK+cdvV7B/Q5bGBe4ptETl5MJvJqnEtKcTXT
YkN+dwdz0bxKEaKlcK79Mo1ZiaIYCOi5FQaAmMff9Q60e2itxafUsPAjoKL6PnIZFuNG4AeMC1UE
Mhk9SI0WF/ybW7JARSnVB+zwzBWxvx/PhmvlkcoJUX59J/1R+248L/zY8Tl/yQVuEgZvSeXxRuIA
6cZyCCcEpxxYpxvvrb9h2eJEu8QrEg9fDkcPyp1jjHPocO8YoRhK46tmMuOD7BLLI/k+/KGpGy6X
PzbXcbmrOREmNOtD9K4hONWrT95zsf6B/Q1QeAiwTKkHZXOLBZX6R4+qjWDty0dfY5Dbz03Sr9jw
+LdDdKXgo0F8NLVAz4J7NRL0pkPmCIw7YnZYqwfBnMnr4zx1eqPlhfRjIzzho00OY3mWL4GJ2act
789Z5g7/qRher3ZToPBz+qsCyuVMqe60LWKoxacbYClrd1qB5SBCHTI8vB1426Erz1/wLWauufOA
5uV04LL47BTiWgEWjenFbCiTN9e8jRNT73Eoy+cvV1/Q8q/aOyB2tDmZsEpCccdnEGAF4lJbPS0h
h9jQmoQhxtIX1lUkbJ18S+ExnNhvB+AG/JPVjF+/5nM/KAtJ38AddzR9gAKC5hBxVN+ZSjErYwT/
eEhEHZ146kbMbruLGUPaYaL/kxH9Wu6Gn8hvbDTufSr1slfddGfB/YCMO3H6kSQXgo/l0gwTm0S8
JOQGAKkUiHvxZeUf9zahZKkjEUGylvUmfFLan2WFJdGB+NKqO7J1/U+KoORNmlf5xt3mjU1YlBp0
0T/bEoB5eOaywdOLnGGnI5vM11RQKxkp69P7iffygPXJkD/MNT79RZaiNrtA8cYONpij89pTS9Mb
sxPxTwoVgHF7R5yv6ecWLr3Gp7pBohG2RkbmoxkjG//WyPTahP6xyXX3JS0xHt9HqA7vhyrfyki4
3V71VlmV6TW00kqIj9CllOYL0ARTD2EWsxuIAXXcZPWKJw+qyFb7Vya6C1fUMKyGwCfeeDvHSoD4
UGIp+n+4D9Y7gsjgR+bj966N8LZGA8Gw+xoxuRH+ZbsWXFW750kWKQ+yzDI49tVgJSiApl1mzbnC
wezPek61KzCTksKprSHGhNrCncc+8mDWmL3x6t90Cnko8pi7Qs7ivDz2fz+T4Za2iRydc+9xql3I
yz4s76nf+yviqp2B+Cyf0ioHmfDqPCeZNyqXLfxNXcCkljOb4jXQd0zGsb36FgSINVbftzopPm+V
sKMd5gkripxqniXKzc05KIkBctcvT5Bkcz3vor1DvNXSNoI+hm72HWddRC1RykzntJgQ4NlJ5DWI
PaJcmSSf7zoT0w/hcpi8Ca4nFvdFtZEaXPdVkAaPHJQ1mp+NNIW9oZ0+FVCqJ3+FQJGzgWcFxRwO
k5Z8GMKEbM+CgUaXEcAQ+HHnJ7z0++J/RSFJyKkRBvQZ0JGRVvJmlpz/QmuZbqfeYKYkk2/WOhgI
V0AU66hi6FnjgFnIPnd2px/xL6OLbLuQ3eO1Z0y8ehi/vkmqe4G6NNypL51VQ/yIsLPvsKEDrwAu
2dNsU/grDK9urZOXZKwBuCh6DvhHPfO4P4QVNCGA+Dmgp15PRIS3Ax7PblVoVDbjIdRbyAIo6Yfu
HJQ9UbR3eDPMS1G1f6L/GgqaItinEHnllYT18z3pw9hsSFnxVCDlK159liWQw5a3Q7APXERmSZrx
ntP8PTfd4QZ53kBz17ahonyB7zjYMix+CZCZRs194cXw3OdaaNoFAC4AtAnxzFJwfKCTFAwZvGVq
3XuZVLHFNDKYRHy5BP5QIhWpLpOEQ24qGo0tt6V7Mw/IQlifofNNrKyZpyfqLVQ6HDdFfdL2EPM6
6Z0xhBm/gr7pS1q8V7ss1BvmxAAw74JMToXKjvVsHP+L0u6iadoKYgj/gQiu+n08MPvJvDoHJX8z
siEVDsDuo5kL7PzXpsZDOOepJqk1Uc80hG7iCzJa3CaEQrz7OfZTYUOHhNoPHCNzmb3EXVI1VJUu
ezGg6iXQDqsOV/OOXXFJQ8ZWVkV/VyOClCoq3Hp5qfPviztTD6O8wUVnpyM2KXJ+XPO2CVeJ6STH
OX8t6jxVql0L1+femmNUOiEvpnxt5WbFSVDEFfA1WnXGfXNnpDWdtcc7KMeE4U+b7jOexk3ZiNHE
YV5vO13pB86ey0kWP5pGaCMqibx8AdgEhnqj9+RB81H054TfMPvfjaeM2eDOEIc2tI9291Cym1kx
NV4J95ueDD0dsNzaauGP0+gSIdw8Qh75YC61etxKrAk+2JvAV1JdkLTljb9bMArpsiwqlQWiVpaR
3L5WIlPdUVd3H8T2c1AEOBh8apbNXdmp1xDnz0jhREheBRvZYdN7T3VwscuHBgh4j980yabsZ3J7
z7On8zh4MC6DhGPPUGAJAGYHYmWsnmMXOtHssBotIyAgrcZ9MRhdUtLtx5wgn+Awl+jg7SpkmhFu
LOJIDJi2Rd/WOfyHXzdexK7HrBuvjWkxCUO3Tnr+YReMIs8JXbQ4XBfg424mp2Waz3zpNJMPBbqS
o3LSPXpe0Sfe5W8px9n946IDMeEed4Xu2hXXAQLqkmJDt1NzWwppIUyM7XTgEWkUKB8bnHXcONtH
I8nYd0df8xo26nKromNUz/nN6MDJw1bnhUHNm5P7EQ/PyFiTmNATSZCne2VVsW53CvF5bzX/CWq3
TUMPJgXq7lcBAciAGrU42LBaertAOUiqm/dBf8r0BWsk5HPepOKFRSThdp6JVlSf3OB7hpetC0dO
oqzMk2hMCI9Z4gdzlpbGuRacN7bwaYzdMIBtYveqm04XI6LxN3W9zWhIP/2qHMvWIKLhgZQHv9lh
qSOkdZ7815rZbQbOWYz+5CTHCQl5EDJhHHX+Gt9uYCavqnwtEE6N7LGWm77z/1v3FaDd/5ducTcT
V4By5PsjKRAdApgnJEJmcMHkKgwYSX75hzQtSGjDU8ed7Rs0AFI/isdulHD7tUmsmXWV3jzAeJ1+
jYTapPkSMgNTrZqobqe1zgsaZnZF8jUGoGUWSCGjeS3A5s8W3OrivFlK1j9k3+9zB3lmkKEgwSjL
Q4Cyi5YwXroo8fPyZT1uVlvGK4VdlzMZw5/1ScB7eESd5vhBIhvT7cSSVi9KcuivKRyXPTCjzAC1
xfnZP/bG47eGs5nXxxcsaeUXA0LDicQCycaD+YbixT4NqeIwajd98+8iks2q1ClTxLZVDwC5zDld
pQPzp/gSMjCV1xxtzB7SQXJ9e2KvdHCuJBV8NjqZ1ln6fmlcLkP3GGXQOS+cd3WYgF6CW/Z93bIp
5FEO/2bOCSpQ8/FEvuy6lVQhH9mNadVQ1TQWEp1B4VmTrp7U2/kvZfpkw/lnOsA7tqe5v6x5fvmX
AcbeyILpaMdsZN2DLhu7l8MHPSZcHKnPUHco5D8BkQAn1zXPq24Ot3cOFk8hvqeKd6ALQ478dd4N
k1brfVZUUJ1moYDHT0FQwRNWjmpk5wRHinapaBQztcv6K6/ebIyFeQCC8LrGocUkfUXOtKaDWQ2B
G2QKnbunvCkcOfSMFDl+cYgHASfn4yyKuYPVsuM2y7u1l/dA6NJE8lFnOmLs81hPiPj9KQIFkfsZ
JYrRaLLJRGX7asyjRJzXxsu31amKnVXD9330zndAqkXF0WBSBNDCvmb9RmIQbgp9V2HO7QuTyX3T
f86qpOzygRllLX3xULEnHF6AA5KB6elDw1JkviBicL+vpgjDHta+KQ8s+cGFJ0TfSC4EoGg8ekMM
dsJn9XFCQnMFNNyoXRp2G9HQSCkvz31fPKMB4T6Qygk/G7zhEtlxFSoPazQ5PWHGNA3Bij0oVwYt
Q/jhbPWpqb+ihLJqGNkFYEL1VYSmwWGOV8LmrU8grVjup2jcWkJZ6YdfYTEBXvxUiCISxVoWoVyP
5AZi+KNRoI3L/1cuuxhVFVukQr3TgVLS5gouPY1pUGKwA4QK8E0KE3dFzrhwR5xZefWuqFm/Ck/8
jSGi79gqrBV3z2uSAYpcAaTmj73MEZtopsvG4VMS5uK9ucce+vybD9qWb3gEBYow8Fukz0Sb6DAt
9WBbpt/WepxBcfe4543FDe7qMBpPAjM6eKxEyPRM5LQ/j8k1RdDHWbY1zUWqd1SUDMhKHfdejQTI
d2cuYUqfeb1Rgc/S14ErPxSDYO/uukW1vRx+Z2L+5WZQz1TZLn3Eo/QxLnulY7RnDt9LAMfdbj5z
lbk/DN+LhHA65KQrxvEQPjjEWvl595J9mUcSIRfkRGCnl9GJAJMwiReqYKd+FBRVAANplafZnOC5
TxEoZUVSxgWkzKU3XwF0vfmN4S+qHSYkmOiqEDJXsDa88XMhroPNZjPpnwhAoLTue+aTIQ9Ho1oZ
n1rAQBIKgT2VEH1k9tQ04DFB5VUbfhPombFqRnlbamBN54p2KeB69xsuZUKL0UxOUgwxuvmEhr7i
M4hdh1JFek187IuNUrZi83Om+PYjHdjjwfoizhiq5giloBzWY+hi1pjt3vahf+s1C6YewIfRvDhu
+az2CxRofgVjiOdf8IJbz0WPGhmd/593JOort2xa7fgZqzddd6AuhnjHIzjkOuWfrlMaZinwCWMN
gGEGfLPtILtlxELOQ/Apk2dWJMG0D0fAo9z8yXePa4QTooNxZaEyDXTRpgKVwXuTjLgaOW3RPml0
uM4SrCspnpg+Y1OHrMhmcvK1V1J1MVcvNxP2zMcdtf2/CVIr2gD9120LDcAZ+eudEfGlzop8z05A
1LhEBeRxjuVZnO3OWZS27QoH0cwOaQYh7nkiw7JVpzzW+LBLKHndqfrdXEjkI4pLjI2hdVwu/fej
eSlrHPMtwlRVSw8c8wWt4GvbIGMVGrO5rTfjTo1w7e5Y8dQPiblAsm0Ck76lWH5ct9NJz9hb/us+
t0iZ4FtpqB+9AqqiUc3edIv8uRgD2IBDNP4G+L2juFXSN0uDR8eBgTKL0U8J5psu3l4CyUNOsgRT
O2a6uVI1Iv3CoT0poCvIBJLvx7QFF14X+0Ki8zDwNfes/utjrf9uZs1VV5O+xNjoiSglBmAHYfGG
92up8h2I9SyWTTBOlL2RCE637FSWVdbqBDO5lJe/8DeMP6THm9cnzaIB3B3VvtJykoZhLn4bmY6h
o701Da0PDpAeNbOSOhTabVN/0RsFtxfsD0+AX4scQeugaw2OWgxiVEy/yXyCYidzf3jRfbJrHnBi
ZIve0OaDcD0C1aGRtv5s3aDEXrt4krz0CMUJNs9zuea7oKTrt/An5KAEKfJc6EkcU5r9rgSdQa1q
4w/3L18zQXDueVeR9XhFLZpafvRxjNbjRmt8gL7vssDHdQuhj8UWDxKCrGQQVP4l4QemzCrwAe41
WvyMveXPnGRmCvHFQ1/Zdxyje4EBnrFjQqzJZYIG7LkdizHb9z+oOuAc10/O2vnOwQa0c4P1O7Kp
ylhG8dH470QFj6GMbkmZgtMMdBwHqm/dfOustXUZR71oMSRtMHFxlnoaOhmNI06gU9cTYU5CHaId
07ilNJTwy8Xy455nWJtQMV/jLk/th90EKSGnAbeYPjkI0rZf+/JvaWv+SV+t5OPWCAdgXhlPrUAu
kBElBPjOX88HiaJHpCiVkJvwUV8pbPa+mjGZUCOjmu9ORtmBkR+/OJkQysJ6g49g6rKY6bLzTYMI
sOY9ifwmL+2JXQwuBsd73hGAKysmpBfhUzwsoCcyT9LBJ/wOWLvCfcb/v/HHjj1T2O+fNT3/ZiZi
riKiLQEZLCdp3Asv4hpBinhgcqbxwRCY5PaGUWhw4WiLVNVVhm1M8Ri9s6SRY8CFKtj5PJ8BRZkK
gct+AawWOwquQ6soGmqVBZI3paDsgiL2ZERLEQ5pCK8hbG/XicjIhBwMPYRlKc39gouW5q+7jyUw
cEcHgrAkgfG36AnD4sewu/6gj7MeaoAcAtvyTPf/QIpd56mmZmhrlewbT54mvDoSMM2hH6SIly3S
Hem9Nd//qewFwJXkeBCIAUazcI/oH7RatC+K0eDpLdns4S8aUaSxo3JzdxyHbBTGhHLmrdmvDydw
QIyilgsmsarStPbTrpeHq058+1KI0hucajsJuH2REyFyoLllkfuKq3o3RSXg7V2e4/Q1b2dAcQp7
X/zd1f69k02kQ2PdUa8BPS/VZpRkkxR3EV9321gEIDDd37y52p2OONhRmdU8KQEkvdlZHd88bqEg
PMcYKid4CWbp0gyBTLgEH/MahBfdNiykW0FQOAUwxs0pmubArm9SYD9eVWn+KwSFWoDFslmzqqBo
kTKjHi5Ep1UpkbK5bRFJhAKTaXjviNN6HVh8scIDh6Sq/1EJ9xTwgHqF4su5I9YA7grfXk9KV9Nm
rbXzYxoeZYbUAzpKRBay+JajTbzb1GYKGjJc3d8sCgQWxyMfpG5EmybrGvz/bituA1EjjNkipQPP
iccenNZ0YdoErq0pq0XNSWVG85MYimSTNHbvbGyQ9cPw+RprB9OgQnaqxztE0THoyIapmEUcx/1x
xTQje0Ra6yU/mrZhd7kdhEE82CsypK2WvjN9ut2ZgOaZfJmMlVOvz6m91FO2h+lq0ExK/ZgzreAV
mNbp4v+gfIPZd9J3jBceHg8dWXbRPN9r5skaDga+qppQEe6HZx1eRnrLMOkOSRj7Ix5WZgWIzZNm
R1/P532PTccZetbn6KugxWh50JtlNei81dU0q7Tn/zCcU5Tjqx0q3IA0WO1lDdWSCurZGLnfb2xx
v+r0FIWTIERL6Am47rYUFewZjlIpqRHK2YmWyhlpkqNda3YppTP0k14HK+uwle+YWQECk71OYIEt
qcTdUY/3Wy3K2O/Zi4ZTmg7c9GvjHtksiwixzstRXat1UGBwwhfcvUIPiFk7f7Wre2+44sZ7VZWJ
VMAX62JurCW12NmY4Ac8HwHpQwbYOOu9iHYpUWuBZ1xhCOtm9WFYXDmSMEwqKgh7ai1xQ9pcbkp5
hViATLqxsZAc/2Ua3q9+N1Ix4nASc6M7aOFzan+EcdFntxUOOlK4N7F87n3/WwPq/t77zn+LRvod
psygTg8u2Gsmja1oA2kFcfJ6RbSiqwo/vQTCB2urQRwchl8iHzuwvza5y54DNBD4Xb4aqCQ0tfcl
s4pe/dGPPRQRBZmNXg3o2qxdqrofvmHw8UvPsU65bRxif7dU+3bV+7vw5IBboVFERO0HzpqkI90i
3NMdN2sXvuGC52qOJHIvawlyr+OiODZIVx5TWbwCQFcMo+8sZRWsEicJX1rddDyrNvuFmhInjPi0
yZs2sfF9LSMB/N7c1v2GauPTKWKG7jqiHfhi5yQ5x0dfeG/EUazWYDsYSxK/kWZGVljaA90b+1Dr
f5FAb68g2UQglxhARA9OoRMdEf9T9H8yx69RkbHwHd3td1sXGtMGppHdiSiM5pRZttxeSKfUVAre
xPjSI1FBzXPo1eD6XDcyldgTVOvKKE/s/Q60UbDKNa5MFD66ROp8kGeks+/68wdmdmHHKkPUClR7
vRS2rQaATpooyzy6+xAZBfcak45ogo+MeSZuFuJvE6yp7oGVvLmCWiOI9Y3x8r4psh8bTe6+pTtX
4G1mJ4mpMJnA9jDEFuN7BDev63N203LPxIW7PbHx4er+7gYsSKQzbyOF8Gb2R6KxK4C4tHUbcPXi
psx7Chc4WmjrIrEXXYfah22gZ4zY834vqAcAL41YMbBZs1GpLDFGjJaQ8y2dZy6abcJFjK51bvM4
AZ0kdF2eWjm5BYhz26swoQNICunzojvJ6lQLJ2DVMl0+5BTZFfeDwAol9wtFWJlsLBqfnNPT893N
k37rCpGMOqTw8hLC6fgyy8duhFRBRFEy9sFi9A9Lh5C0KUvI6tQtY7DSW2Cf1HUTLzLX5fReVCu4
PNflvqXps3T4mQL3kr3H3PTrzRHosPWJnJWk3s7HDbQNyHW7JHJp9B/b6VabsLzzAPkE4JP4/6pf
5+twwAlT8UtmFBJ0JSLkQ8AztqIUUmitz7hFpaRHe65wNB1el7cUtI7xIAeeFhX4w3vA0tRcraQV
KyxYUbIo7Q18Y3dysuq2bQH4pYAqXJHbJnsrmkfTJ1/Z/6qCPYlOAcpdHC3OUCV+gUasZuIgOsKS
5zvJmjLzaYRfQ7ACM3zTZe7eFbWH6O4ScRfRQZL/XOZwhX5tOeyt9QFY33AIAiFzAzvViGhVzd9h
Q2ZFgpkzhJv7qgAnwlnNoi+PemsYn+PLCBJ3KnZBCxtvASlAUrFIE18mJpZctkZsQbbNrqALQiaX
jcZ5Ny4pP2KJmjW95ddc14II3FmBzKZYrWynVrdc58l2DL2Vw5OhJ6homNznCFopFRpTTNexS93Y
b0ohFQqBxi7EZ0zJgjDqH9fQ5rLQXClrRwvLUpDG1VWZ/tAo/GCh6kpA18lSyXS4leaBgJRBWiwJ
TrYzI+aoC09Jcda4TXbnJsY9ol70rIgKALnfqhAzG8oXI6VtzzB0YZaMA2o88yFWmbnP6EORPMC4
mNsxfrvz+pn8ZvH5XefevNQWji7aDKvbyh4+Py1+JJLRkAzhOHvdU0nzM24w//CT8RyORdZOdhxG
lOerVzxz0IwALslvV9EN5Nmkv2J+/Vl2TU+w3rbyCWYpL4DPTz/qupAtIV0hz2NpR/nYk+fxcn8r
D4MrW1Kobay22YkB9zICls2ObocoN61vVm5Oa/IRg33lkhXJn33YRBBGNj7an0q0GbTMlI5O82Nb
ZDg6COJYIwVc3T2SV4hIsuAWQOJLnY5CkBigrlZAUO17pHTTdeA3W1CscFHXzuQw/JNmXREVelJT
kSD7XOku/KFXXtUX88mFckyO2sowk4ES5ZXVGJ6QcdVftlcpx/jC6RPmIib4xf+M9ubRWCI6ALHF
Xfbm8hsWWe3mIYbk/rAGawDg2baNN4gGXou6q1BolnBk0R5dDkmmxUjc1zTBIe9oQGJSbcuYo+r+
LOR23w8Wm5Kcl4yeurT/jixsk0dsf+6XKpY/6YdwPlBnY8x1zR5w5z/TD13PjK9DIKaJ/2tpxNpL
vJv9OBtqyOP3j+vTJsndBxpGAieR+m42yrBF21+Pi6H4VzzzEUSLBYnSjpbhN+27vNPdALfjVAMq
dzJ/5JSbKVv/0baB4JIXm0c/YgAGayT0FnNCsmfPkKwvHMU+a1X06rK7IPEadK1UUjGvOYw5IYtn
uqaQn+z11IP4SKrGu/kLsWlUvwUICS3E27gstJddOCJjcge/XAdbt8lcwrAl6hw/ucp6tOTYzrz9
deCe2lsuD29gfzWicWfqqhygvwCDM5fpqm4w8WtXkyHSIT8poDbm61Uk70YSkf1dcWMwdK0VsKMD
O7ADdobTLqLD3qmBZAIM+gdk05wpIxmC73ZxlCBQlJVQySK5G4rje/+sQ2HkcCsP0VDhzms+Lmh/
4z5YezsbSihcfEukey/XhLHn0tsQnAUEyc+/EFb0qmBgJu3HRyYkrLLQXLuM35IwW5uURAhC3XWO
j1yoZjmfFbuK1RJWB8K1+15utJaedmiDnovQJcMsOdEey4oyRn3V+bUmHg+FFdnqiOCFzH+uQcd3
jknE6a1VjCQdpwB5Uf+6ylyZhb0uv3ZTeDxtsouePHjO2umh2hfeLJdX7EeeISr3AC98rSapoJ9Z
JNEeLIby2p42Adj9zDNcnOAuMyGQm5FthFbN9nE1M1Cz9Ayv9Vd+I9bbBcGxIGuC+yvjavgTZvFW
/fVy951EVZ6mtKuENcVRuJirg6GweSuKxA5SpVFgbzA6SbnNBlx2nCso5yu3odqsQP9dr2oXmm7r
1sqbNE3Uni5JY1eWX7/zQEYWIyTFDrXvUyzZqne1jS+djQewVV3W14aRpgSRi7/yeKnAj6BDmm0N
qmGX9JxLwaYp0CfAvquy0nBqOukGjvM99xTlDn5fafztbnYVWoc/crmDzzdKAbo37sPVXc9nU3Vg
BsUa4TN9KOep2wiaDDLQ5hEjINFE31YcgqKl91NKCcsffbwRl2S81Ycgdpyg9IC0lzIMXidfoQ06
WQ5PQPM2K2HT5g1WGJtn+5Ui8OiT91GD1dCKrpc7zb7jJ1lNt8eVkXZX8JicCl+z89628bLfrE6U
WDRxPm3DAzIzA1SWcen9QSoXhRwmz/qWFKTFMJo4ATloD5FF8u+SaG3nipv9EeeyhCDCuQux9uPU
EluaH9jBA9BsEAgBwg7Ym7lFgLHEZyDqtANuCpSLTtRw1dWKpMZCycsRRzxZSjUkWqMq+7XjdVk3
ryl+gMsWEv5U4YTXcPQFOARq3y4mE+Pxfq0ootJkiE2AofktOKNvay9zpuLpUiBn6h2I+KP+FtiA
r4VPXSODlnYre9JNle239nSwLoFBk7PKRtKNx+t/CzM1YPuuojSCz7Q4Pg/PYletclpjflNyXBnj
jWL9Lr9CZ2kBWds/HUwd3TjUH9G3Ze2GXnLDWzuKbhafGR3ouWqjDFvsd7+oh1+QDn3a8L+axbqj
FR/g831qbgTEOwBo00AXI35VU9p8DzUVONIIGWThXqfnatWziN/0JXA27lmAAxUiaExsFwVVQWGk
3raizpnBvqp7HUZOM9UwlaP/smclKe/BpZlSZ97YRM5EGH5jf3yALyMPM1ZyCe4lLtgN0y9ndUBs
izGYoWDn0sXP9MgxYql+vOqovRYh/aYio6GOl6cp2yLeE/7qpVsGRj3sToFghXn7l73sy++95m1R
rytKWn0iUMh81lq3dr2or8zM2zTuXlGgbYCv21Gx9K+qG27EaK9h1/VJ1teDbBGDyRGBzK8ZY8uJ
EEV6W12IvQhhYyhlwTh9DXxIifZGU4WMCSkWDhQlFHy5Eyz9aaA3+yc+UdzZjE/3yZYpMlW2EjDZ
g14Of9T5DO1VdH7p/tyhBMUcd9k2KvMtWzFx0oKBhLImyO5+c67eK/rEv7p/Fbpr+NYF4929vrs5
hsyKPlNZbrPORremKSBFDsvHL5XSUfGDTTGwtDH6lDM8V3IgT6DoTggxrn3Lxs+PgkOWa8QKkkZQ
KFZNyR5vf5ZL5CArkIvdN9TdURqBMQWLPownrX6LjcE+7TffGvMCfoJAaPV6sSTRIAiFi95Ebbn0
ElDuKKeHU/XueE1ZjE4HItpX+m1DHuvH+PzxOIT5C80i6i4ILGJ3Z6Uf5u9d0OfhEq8MTpAc5Vud
v8yzNcK9M9jrw+qEh19YGHCFL8LSrQA6pAY3sGPY5XjW6T9KsfZ3vW6Cft8pxA366Oygg8F01a+e
Ez+Ri8wo9x40BC053dFDXTWEC70lqhYV4OFCWlj+2Or4+9JledeDPA1iCMU54MnVm1h8zU0I4KyG
xzLvxz1X0GiyaFdf0h2weUL0yL9WwZFD4Gij8iSXs/dYsiQJ3GRpvsDKQinf3oHhSqFNXIq1vpi8
doqLscZnpS6pFaXRXOQA0dtviSdl7rPrgDyC87EA34dfvyWvQ9L+09Zi6p2hIqGMIS5X1hZS4Ngd
cj14b/ZdNmyllrcjENZHlPZEg5oqno7nnJSw2N+L0FCPZlxPb2Q2cAK+HUg5axyR8p260JCA8h4e
MbkpMMz3+kTIPhIaZTOt42JQfiFF0vsBOeWcsT8YqZ7443aHws4Xwu3KcqGtfYlw9GZ+YN+U7kGS
OiQhAx5nfMrrpR8gepOo+kfyQtiQkDFeZHuOAbzq1iAbLHAs7Z7Xf/qSSfqlAlX955jXGAaE7i8S
TdQ2LhWyVo4zF8lC0EwI5gae6CKzMr9F08xwHz6iI7IcJHOk6nWZbrgYtba5bhSW/vhyhhXM/TGT
kAVtU2+VhT2juzJolJrbSsQ5iqKZB8d61tRowxu4HRigkrIFKlxBsk0dbxO6jGlx7sjF/f/VAVbk
rw6TJc1ydNq8/8k3aDIAvuJ+wo2fXEO+xZKhR7FekioanSX5vmvnea2aAnkStibvgPPF2wkxoBuS
SBS06u2Vu8xw1Ts0a7skWa/lQql9FFvOZDfIaNDfH1h3NvTw8fbp/K96+N5g3q4ynG9a46GcsNUa
/eCQ1DYVLGgDDVISZ8XvyXfLjS1vRDMljRi36d0kfJIsjVp8mOdGmCfCNbwuJ73RzamHBbupiuhV
dk7teWHPp7Kt6N3ANxv3ktGhs+5dNhZrmnAD6j8k3noJEs8h2Lv99JQoco2VRheJ+E5Fp9BSZ43y
lyH82wF/r4qRdm27Poi1yEE7EWKtBg/0HTfrDxIuJMowuIkKqWPkHyEacSPw+QPzklYN9+z0T6qI
p0fmlqmrbwb1xAt4zAqHdtV0BlwTsJzNbvkZUrkwBkdLNXv1UT9p2gt58do3g/6+NMumfPQhYq9R
/G3bYT2kTxoddc5PHIZo7PwYy4QoH4xZqNoTpZ8ygnISxftf86gV98Rmz//mVeg2dNb6HBkYCmXT
JTep3mXQviqpQdFmiiY6gLsuc56CTFcMzWredSCZI+6PPOnNL4x64S4s4iiPmoVYMmjSRysUep7s
Sb/iV0knFpLA2yehDeHnAqXMiqPi5r2Ux23/H61gE5o3VAU9x2LL1m1NjDkjnG7DrFuXHy3h+jOx
UlSlYz0EVZ/vwvlUKOGZvfRLtYoUAqDNX3ACah3VnfUiFrhVJTOgn0Bet2ZjT0xsipv1XFoMW2cU
eKN+pVvWWdP5ZgVFJtP+fGrXYduKHXaIlqelK6zf/0uKyC7uy1KQjaF3aOiTeNY/xYYkiiOKkEWD
BUda68xAkEfAfDpNbh77zfwiTlw+lUjsqtwxmZSswrRnFxTZd7EbbIjBKJuVkkFNxHl7VZ2cIteR
dIe7YuuHaGUVgSw+RnHpwDV12BsOIvvCiYN1BAkQq+FUxXdhjqYhs5gPavUGZUvXIfyLDcMgt19R
LH3mnaafLOlIoid5+z+KFKqxddhk+XoTvIk8puwEhDTkoyj/da/UbNQgsAoQ3XflhY01qWK4amYN
LKxPT4O4GX8DqV5YY494WfvWUMSXknYJDDbJjswkh/lYPD5d8NX0bih5e/x4Fg6t0w0OypvHbGEB
jP5gRzMd2s6gf1O8ng+ZAtC5p/3vFbMo6q4G0s0XMw0kRkz6Y6yEFV7LdGLPhfr5c2cd6SeAKPiZ
oYZShQbbFyqe62z3mT8gbsW9l3lujDL8cXGiVIbQafWlb9NFW9l0TmpgFzimltFhx4pbwUzDcUA9
vslyMJbBXBKOc34AZwyPxo2Wng2PIjk74/hU/59zh/kDBqVik1mPHJDDfkhpGdgHiHHn2HUMP/6B
eL0B+fO7Vr40I/AX3UDO/ckt2bUKAWpEQ8vaQ0YYA38FdjYPMnHY8nAJD9Outzf75qMecrp7TJ1z
p79tHjSARd6lmmQ/Zb25Isw3aXodlVrIVeezsWpdU6OCjzrsLvWxFXjmnFm81EaeAI8/lp/uIoG0
IjlxJI+CW/nPw4JzMa4Aj+JWmH0jpQuPWZhLxgOvsgfuEele8N7EZutSKCjlKrOAklyeM16U+Vji
aGGGmBM7lR6ifL4RzQ4FWTEwJsC9u4ErZXJWNY9VX8AbeJjQW1DcltkiH1XEO2EjDlH0J86OU58d
AXp4IDBOw1v+BwG6ewZ6Y/+6bSsjCehX5Tn5kN1+J8sK+3snwgwEs/8FUFQR1rPllAo5xywDAU9y
O+HslymCPE0RHw8a3e2e3eP/sPOzDsMiLk06F8T+cwmMiP82kb79/iI4dOvZX4LVeXIEhSx+aEI6
8XIuwoPcejIy2rnhfkXdUfi4yhdM5fb2tZDlo7aqGZulPAW1QRUKf5wcadhzZXlZA0h6namte66t
uHBmkukerkpKCHGbkJ+zQYPqq7ScVxTasUOtJmiMiyg7MSJ/xaL2eorJoYysxAdlrH4jS+IFdUZU
e4bFGTVobFypyWVGQu3Yol3YdEXj58iVm8yH/Lqui6OolA1/OxJJ02U3a0XSNHjuliK5UcvWkzj0
i9bIG1Utd8U3ZM3+b6QwsuuJrXuY+JU63/uvwragAmYPlbDlTelFzyfCh0LIr/hOj2rl86iAvbNl
JVv/trjwoQLOonFJ0ZtToqFb3RTxu/Snu7wgtrSFGV/81RNlkOgWLxybT4E+TboDBOjWKyp2MVPc
8c98OCNiibvFMjiqNbJt9PNH5qbYLqqNPeWBU8bplueD1H3FCDQLkBRybYQ4e37HuXP4XxsD3h0U
xzyx6Swpayy9wC9A/hOwAv3/2VjuWLknH05cVk25fe4NDsGSy3NvEuE31vt/oYbZKTgHs7UAmacR
/YTFTcLQW+8ND1zXdhg/IIIOOwcyro2toBWylI203enEZnmlmUElwCETA4AW6lVGuRIEfdDIcPxJ
CBSwzzEkjnZckhQXhJIJz5GXTwtbDLQrHxQ4yeEToxmicIlhv7X0iDGGscISGTDtXFliXsJRmtBW
K0Lqt4RInkW3S8GlsSl7hITFJe/dS1V2qiGlyQnB/yrRQyn+DCV9kZDruvZSZP+fNZPBi8S3ierU
5aNGE7TCdFt/rv5UoI+IGzauouNvX+R/Fw0IG4Oxnhuv2ZXADP99tadISSDUi8h+FOf728FqHQdX
y7THe7AdCFZQLDBIcTauTCpZUERJ0c0aPKb0cP8C+PxWXM8E/ogJFQJt32G1NfHH54nCeoXqz8hp
qEkMy1IPnjOr40OURiksKCBjD8vJoiTsJdCVbyrEyuSdwQUtJaGpytEYqdTdxR7idukzy/Y1zTEg
v27fBUBqpR0DN1m42+2UB4mhkq1EQblQHQ/9E0wvYDdrDBTJjzlAWH9jqRC/mfKVhW4T2Ftm/8nT
HTp41mMMsllgIvj5UAje+0J9Zx7t/N6yHLpXpRYMBAcbzFvgiSoF19rVajYDrqHQSod1NEsCFVyM
OW6ZjwXOSzb1U/ymUeAYJZUnWh63tiFrOsj5je3mfANptbNQoIMHVyoILEDG3aqq82EoVTbqDB7z
z5lvN47sWdmTo0ZFzhP8gwhCYOjbnc5tPpIm8/8+CV0OAjMzG1VZj8eQQxsA8Z2nJs05ngTuNa6T
DYceazai+cIKbIX+Z6A9GcNXY8BpuH3ss0QjjOsJSWznBLGCcxc6XD+jZwouHpRu/rtVyghsOADT
+jAkims3VVcodtNrjDx21Y53dQnOwjQ29mneW4n2+nSMGssHlHCBwom/DV1hDqJij4swaRolBWN1
KqkfjpuF2Tr9P+TG5sRSExKdv9XtqM6GyWqLP/Q4cq9xvw+3fTI8YLlIOiMTlKrDdAmA1UAsQbA5
6ni3FzJ5ihvWwfhRnKuNtpFJ1CW5hXXr8CNxIfzw4+mx1ZWQ68XpAaygJXToDfbegOL5xC16pBH4
09OkWHfbuxtQd/QJJNoOfOvKq6p9AU5RdFi/v1jGdttNr6iOtyWVriNXntSQFi1hVZbMjtFdoLWX
L9Umy6VREjKZ/UPlNDihBGRFrse1Doehf65YyX3+1hgrDhuWC0sYyQB2B3uO7YZSzr96OK3W4a70
ddSJFlxETPU7cvRue6B7hbDdAaSLhpmrMqYnKsR9BmeAwq07p6PVO2z/ywFKLfuz2/ql2DsElWAP
wOKRRinN8kAfVDCRD1wv0UEUZEJn4IACWeCj8p0RSraJwSa70I7oDzDDMlfXrRoVAWMQD3Oi9m3Z
qyngBcYf1OpagPeqdUkBUSqoFYVXmb0oXBBSApJ8PtXJwLfWo52YAxsv2ux2rG9TxPRsiKUuCT9D
u37Hji6aPvdPtbDEf1bjvo5fr8SBTE3PxhR6eZj+9LymEgBs7uUUkS+8jvL7tySDz9c74IO/yVum
lg8NfD/sNcvbvuOsNnpEZ3P/XF1YSA1kd2LrdeuqQChuNuY4shPowk5ne++b/ZSrTPattcTeGlNR
1qCETMe3zm1nYhaGHRPhSfM4kUfGyfYC3SHnWw8/Iw4bMQXl2ZV52f0GjJCpapcUZl42ZKdCWWCn
G02OwSRql+1jnf/R47w0go4UarlhOAv7QwtC/DZDxucKntpt8nWZKcTlUictrxzZntdSxd45EhF3
MQn8aD0wJ6CBniOy5TxpS4Hw8e6NRTNv2ngo4722F59jDwXIocVV4y4DIvVax5kktgwGTkfJbXvJ
lO5wMPrXfYWk+NPJjIC+cSOK7/GCuJu4BFOkf7G1nIqHusjW74snJZVHCLp5+eAi/XiLPhh7s9TR
k8i6SpcYlCpg+EgjHtP2c0GsCJhRxneUGHgs1zIWjYDj2RWVQZgFHq/uJBMiZlBgkt48eIBOFXKo
cwOtwWMPHZHEBxVgm5jgjY2xBkCdg7DSKBzniUIDmZLHjOslq36ri8T5pzNwyWr7bEgekEvl1/Mi
ktTE5or646khvGQPtx7uJvoh8ef7rtPDpbMz2vTK6BJzxM/O6PyQq3QXmPmKD0zi0sb3FDobKZZY
bt8Ty/J3jUcSiUoxx7EyXR6A5uvVOhmndg05fSyUpE6GcmYKQLn2MEUKDcJDFyf1D/WtTx5utUnV
aRse3ovJ1dFWiNo/3g2sIFswRK9T37HZHj/8tGki46FeaDDzdcRphfXXhVcTIBK8nnxxFmj0I5uB
oDl4NHdDQv+YmrNBd2lpoefwfxkVLRe26OVz4R9JozBSVY4Vz8aRK1bfYCJPKtxf6EE1V57jP6x9
9CLu5kXUil7ZZb+xb6yjTkjb6vhUf2sZ6nPwUdm6QbyBhA8x2cn9q3m6u2UYeBXAlcVUJBJUoDbz
Xr6NEitIVnYUrXVdBIsq5lJUVA4u/acaB/oLn0icpbXYwMalxFucK+y/t5sDiAoIw4NyKB4SB6j8
JvvD3aSKCC4BaO5+BnO3GQ4Njy3x7lH0vtvyALgpof+dKl1WYalvK/7PoWVjxnXwtGstemESlfbD
i62tyWrL7L9TUuocRnjiY6b8ehQNnf/TmKdrOR4K7AdnIr2MRo33/kP1nmvncgT3zc8P0gknryWt
lusIgRZ1lzPgHqqjCe6aifR6+x1NXBkYnLKlkU5IfGKkC9iSbrwYuBQA9oBm7TagM676BZI2uOaI
aZuk8+a3XtkdZh9g7NaN3SeyHRmJ+3lQfMHBdPupJQwK5G4JWBuqJQ1RhckR+zF4Cz52meTqgrRz
4xQ90KFO+eL7c0LvEpUbDJ88Vg5LqfYVRHiFDvrtm1r2OwykFyKO2IXJGKM6dqhwXqP4xfI5E8jn
91l+zn4jX5h0yqlzmWvBbN0PZCFqa2Trnz5diGb48u+gWrtowjsmE8w0DUp3YTutLSKCZ89Q61du
UJlzpgnwD1takHcnGa8yv92FP1iwbwoiyC4fCWRJ3Hxl/7+8BdlI0G1vBClz0e4f4XuQcduEV4iE
2Hk5KoMBTERQYCzC8aixpK+JrnLaoHRTTd9zTdRhBPvDsM463/kw5fptZUBaiNkyUp7mFuIGLChJ
R2u11umsYpbQdFH0ovdqb2n6RkTkoDf9sH3E08d34pE7pi+sqMfHqRkNAIy9wr83htjzti0Qtqn3
SuH6VNR7nL/JdAYXU/aYU1B5m+voGcxgTtzkIsK6LYSsxodpTOSLmNaddhXlOojtxdsUTbTbKWfs
3iISbAvIJ9l5B9MvQC0Wahdujo3nSnLmPvApGHRlGu75Pvt8L4unpWcHboZvC7Wn/QOpzGJtdgSX
77fIPuGK7X/n2zjbYJZwZ728vye11R5Zy4BE8OP59sh0ucYGWLNADKM4lWtKnQyQIe2lCK2B0tnU
y6LtIifHJyDneprolv9J1pTldZBazzT4hu8TJl9FouktN2gbl6bsNGZcMfQdSHoxq9gvqa/pWaww
OwcWYaW5Tb/+z6MRDqQ71VPWKsN9BSg6fvVVCPx5G4bKhX0jS/sEIdUQ0cgwWPzNjtSbZEqv4jE1
5eiNL+sLpJm5Zui8NaXMpIuU/b8z5ECz+DzhhrMrfvm/JNgY9Fyd39zUl+LcMKgn95myB1FYrIyn
kJgy9bw9OvOt436dFjTvRlc2uBeMJYdI8tPRfQ57mNP3ZnDztm/tTYcKpXuOWiD3H2ZkgVebb6q7
ZyESlKttbdygLvjXPiiY5MRVVU+U+9vy5ZtXzVnS8ojWA8iwtoDWny8LhS/TMN/EYA/y6NVCp3Gg
7Jj1ybhPIiEdFMjyWmwwcKUjO4M9ga/2wu1pfVsg2XxrUfTuAkEUmq4IUdT7Muy4Uvy9SfactHx8
kmydWjUZVS5LijTaTeI7PPiwDbAcHIn4CkSUwOAo1fVoIkCQWwqhg0zRmWaGCTZ4FzifVYICFOOd
5G1rZq+2Y2MgJag7Ke6BlSWD14n7mZWcfBRYqSPMU8ILf7xdAzOQp3Vx/mrUY4pHbjEf5JMx0KCe
nv+mZl+99h397QPnI+yl2sA3YupXRiKVNopyRtyW2GILGfOQaq2hWLLihlgVlpmAWuHOkzXvVEob
qbBu6NvsnSxj9U2ux8QaSKPWbPu7Qgv7Ges4p7FRy7IGL0gPYlIDo7+eqa1zfo3sMQFaL1cDCbbo
BhDm+vTmzKT/XU0UMBGfeFoxtlo9r/f6J/WskfJd+6Nre3Bo0xZx9DNL+jEe1olwZrWx6eA2iieg
C8OsAxalMNEf6SwCenhJnc3nNUk3p8+OcGW0k+JwgE10BQVCJKWxgTR99Yg7eB5UhV+cTg7UlLrf
Xe3FS13fR6XPoHUdrF92yJzS+7YfczvRClFhqCupBQ79EMlFGA92PIgd5Z90P6/wAqm295BwhEDX
w5kw4e4SYKzVyM11/1pATR6vWSZCpr05/ljZc6/v76H8Fcgktbnpv2/5BjMRx//Isw5Z5Tc1fECY
GGVq+jEXNgTagO9ocbzH/z6/CODM+Xr+QsWVMe0E0vfrMrwz/AMoMM5ExcM8H3p5f5u1Z7ViB5Mj
L+DCBs20ZgNz38+jujzHlyKpEmklbTXXryAHn109sItP3ff7ngRjmKxjFtQHmVrWNh0A5XjSOp39
NtV0sMKJL3xjpgLsFrSmn1yIKdHSb+nmxqUBOI4D7s6tR97VGODzKYj+xou2CnerzeuSXBxBiYwW
D6GV7qIXEKO3R3ygllELRZcNHIOGOAhkCGxDFGGXaeSKqe3isUhuqCJqBZ1Aj/UjZRr8hiIYrEmB
i6bgNH1QUu07tmETdM6aMmdUR4vThNqGr89lo5ZGMRLCc/ucImeq0WWFppc7Qjlu2dEXiwps2W5b
K8RLSMka6jCcWpIu2TctwVl/H0b4zpY4q4QQjECp4lLYDPMX8fuGyRP6bLjurJoleejvbNC5aEG5
WKYj+zOmBZEVDWEhE+ZO2KPBsJLFRpQARy1KMESM3gBUPtRCkhBvE7dkjG4MwkVp2QefXv2UU1I6
ZMfsZbUAQ6M4Usk3BwiaKpVCZyPrHFa9Pu0gOYlN5dBjnW7KOn+Kmztuq0PYQ+hdfouayuw5dXhF
pIQyxpIPrB2/wm5yORGka8FJM/F++Zj60dTLJbpZ2JqrC2sI9owZ7rhm6nNTlrvmqcwa7svNtm6a
ehgh4M0Y4sklesHMeEYOLpyHteUk5JV1gBG4/9BFiF6/KCUmw3Yf5BRuIMpdah6+6c/1zj+sAxQK
3nQ/hHIExcGFQzeN2bVNR13ukGvrUjIK/W4yhu96sxRZoyrd1UyCyrAIlmNTKpBEEpoN0HrjXaGo
1syvNdsXDisfAJb9P6Ur49YJbN8GICugyW1HmKTzKff8LtCCYiU0LIEYP4Qk7FocdJnGVG9V4Xcx
VpM9/ba4rHckdRvAdqf1IbVwgsxOPXMN9N7d2L5nnKZnu1hft61q4Wsgy0oyaRseVERem1+1m5EZ
7BttX6YHahnmj/CnWYmpSiUKiAkANOaCQJGtFqgVYxs31LqtPOcucRqChcm/HpO+0H9hU9cqU5nY
iBlh5arpBqc9GsjXsDmCzsXZo9Y7tDaODkba9VrByUdXvk+WTwSuzGu0gK+bvQ8KK57wM4lO7KS4
+M8n33SBfByrUyNAugg8tuN7g8aZUAUF7oD+FjS/WsY70sLnPSfZkxCPPQOhccNO28OBD83rzzMc
B/J3jt5CZmctFHxJAvz531jaoM/Z8xuC8ulpTdVTwJcLc+MwnZV2SKdCyKDoEpi2LteYo6kX1gXo
znmDIfofpujsnxHFjamdfPK7iIsfNfRVYdwC42R4OrPKMdm1th2uirqin0qcJTIvRsOaTfGyRaUl
mzm4oqrtXrDC7biNEd27kolenRlw7eON0EcCjjL6orINo+f4xnCEK8Oc21ILg+gdcPpcgE/LlUKE
12+ZeRtLsmyHrR9r9PQMQ7l0HgZufcj3luVRSsvmf5Lt386tD55V0n+zGLSwNPA5WVlPi31Pk1Wd
zOGvZtZ/dCv4lMTqVEaQ70b4D2bP2L1zRqVLRKvf+6+UjiLZcXupXM9NXnizJxmTLoS1HGq5ZeeX
wUgvkUhyLd/XaW0dE4PUl1Ca321DqQN7DAH4E4jfSmmMsp6G5aVqPmRYoOABjtviDjGXQJT0+0kQ
QArbljOngkNjtBQDfvg9W4KfaVmSgY9q+8tk2gujbRWRW2QBXB4Ja/ityGJz5VuoMvSEWM/DpglI
W1vQ9l2EZbIkS0mJWrdHYQlLw5f/Ws/dVJSd2pA5EGdQlXKOs9gjPSCddAwnf1PqOE1g8HZPbGZC
IFn3oOhqXVsLnZNMdvI4iUxN5cDubtJDyOcpVLBSuLmgdR3EIjdZEn+0Bzb1YCmAQqVFATkifSaM
lUiaOXqd6ACSICjpISu+50pnkqoScsXQQ0YFndxpyoEzgHXNw/VqI3LNgoe2F0/B53GIJT/wHz4I
RHNC7oLGY1pHKNGZQcvS77/NVYYo+yRFRMclrdKjbIAcb+e5LIIn9FpMzNt2pPa+FgJAgfI9YxtL
Y5otcY0rAT8CSFF5FzqGfSm0of+ZHo6a2nlgs68VSSGSrxmRtiw4lpDIGptiStEEJn0pWHT0Pz6+
Edq2Q7vjDJGIWiRf/xOegPqmZZxSv2/BMpjeo08li6kZwkKW+G6wvuLwkDeQxlh1eciDIWDMVDx8
uvUJvZvf/0ovWXRsBY+Be/lC98EgvFb67TSj3LFYjRosDE8jeQKVCxALNBDJYnB7c3BIfKx0gp+g
7r3GRGF2IatdjRz2x/AEOxPBeORTJMNPeEogxL3Nn1MFj6H4Hn6wq9kpnClnShf3Kv3klfGL5OjY
HGSBBjIvNawvVrHFWDHgKXQMt003P7b5kxFMorZiYaZzsHv154c5iMwfG9llsRyuN+q6aIysdVup
grs/yJ9JZRAulfSFA2dZcKnFDG9hqyF01MFCSF12QVxTnFutYLBpgNJ7d9lQaleKd6Mkv1UE9++r
SHM/290rnb4AhjnDM/LG0nQynftrJqNXfBxkgk0pviWgS2ip5wIDANu8Wcq2rGniUjsI5uZqk01M
v+TYD4gBR0+W5UUa1wTYqrA6eo/BciRegTSSMy/ntH9JfsFa3PDi7G6jC8DX4UxF4iZtGnoiVTnl
uky3KGXpAx7pF024wlTQ95Wh8snqDhaAhYgWh0610+WJw5e8Z9k+wDd40/9SfGFtKx4Pkf6HUuds
zcI8/8oamLJKJ98ObMX4g4oYVTguGd0yyMibtZwqIUAMpGb7/vhUoN8W1BO59e2ALVeZP0kl0SsN
yPcBL7gvagMH6KoWSlxfG4KzmS9wrhtzDVEaZSfqEg8/rj/UVFFoNsb1Z7A4keCY01V1Fgdki4BD
XxoXqehcq5LN2823aRMzW9L1v2vqUZ2G0PvT3PhjLPvQo7z5dE/d4K+wBEHIqsvnLQ6ShOO3R9Nt
rmaiCBBJUi3+p5hDJIw7yPvsnBx7V/mk0sTBtckjGTGxLzztQytJkzFNKkvKmNKzko+gaqOuSCem
1iXDHHqUAu/6ts0jWRZxsCN0/eDR2I2yG5/FsPQLFmbAwSW6nTTXwzxbodFTSLm+azdR5IFkb2tp
Q61ypxdZTw6A+O3pOWTlxKw4zOo94+tzbYD/tuxgjr/V4H/KA+JF/rmq/1v76fdgvhFQ8lQDyCky
Ms+UQn1gehw5gdDVeXl0oc14mINJ1ygHD15IY8SVk/yme69PD4UbbuF6QvPa0Y9PVEjoyFPHBlsQ
VnyIuPUZzfMh5vC27M4q5RwXahd1mvY4ErBpmAz4bTxz3E9QK8ce+0aHXwh6DUK7pf1ArZL+084A
L98ABYrt2iWiRQERiLXVOOQHRnDvA1NdS0xmaBuFjH0ANiRKH3Hvd30OArn/Q/e7jxhrljCZaozK
IsTj4ku0vFNRsctGJv6kcZzRIcaaXlpAQyVEwxtB6tIQzYuyWMykGqzHAC70JJHp3KRMnW0CDSXy
4bnfeuY/I2YvnLOHfsVdvSvVIqQircKxMyW9Rkiyiys3maCp85khpG8iPoZiCRxg2R16TBwahULS
zFs2LdHGiKqrsmt3p8gffgD/AfUcn0EVRU2XmvQ+r2VQ84m2Iww8WNqLRm3s4acUZT5e4/VSvhKr
CfKsqLtx2BopmHjiHUqvWJUgbANt2l6z1L3FxnEMSp8b+JHRgixu5vV1UEEsEMrjB+DlP/JMFZc1
PGrbgJZGK4+QD3Ow+IrYRo5gOgUGEyjgbq1uzhrYSSeOSff4GObzfowz8alViG2KS5mmew9iUZvW
Ja7zob7jdLXZfwpMt9WBS80/jFxN1QtK9TSoOyOBF5sWyQWWC/zvUwRpVJRCemP9FSG6oo1BkB2r
0g0kkpdLlAW8o9hJ/++3lHZMy/HKBCRnfb0+zANiTAYUggzfalxUoWac5hToH8GrODXOck3P8CQd
a+FbLylPA34uUsMGjBqEwbALNjtSNVXY00Y3dAlNzA19iOPg2jGYWa5igsYiwIsgKgW8eri8gnsk
TyHIOX7JNAJczo/mmhDJVD7TwO+EE/nFyFOlnwYhOj0NJ8BUkbF+BHX4kSrV3AaPNRykE6Hm5JLH
tdAWZBcj4IGJkKddgZuLndAfXYFcH++7MeYZRnsRZdtJ6uoah5B5M7q+gPG2Nt1bwVQxQTp5JCrT
IFS6TF3hKhfVYi98IHdrus+bEsQSZZOkBNx2z3UwwYo8x8/N87WColBNsqMdQxwHlj1kE3UvY+Xf
RCe/r2Mn3nCB27Jhqm1Z7Yuo+iQTf7IbjhkARyLJj3uD8Q7+GsBxVe2uvYlSs+jjDOkFa8t36kPy
bHfU+mNs0VOc8iFpg2vEQa34830ppbTSeNtkuyzFtG5zMMeLYtAQz/omU3IVYkmwR8tzPyPe57VE
r95AqbzT5B9k6DTb/z5nmI/t3BrGG8etzOXgm5E7cfCKV+K4Q0haqNk32TS3p36U3XCOwrMP/kJF
+gRCo4ygoDkhjCaBpGIaodu47eCu+DFQGfhH+yxuz32KqFibngwAO5wsbZC9CxTJ+HVN1eFX1KMW
28GFyo5JQtATTZx7LCW8YZCGeLtZGXyqd6JyOrxKEhdKoZ5+v8jyLcMiJ5p+LvjFJTlKdqzk9A4Q
2LUwmCmLXhWHWldWDGSjV3b9YcqcXq7izcSly+XFUnkrXlNZMEOeIyY504uUeCdy8+zv5WI1aCus
aXZXuBKW3P6MIbmDswF+zdwXUyhQLVThKnviyEMH/fctAO3MYGwh14MZ9oYfxOVoyBqessZLbNve
QScmkewC4wZBuDGriHKpsf8pun/1QVQ9cJeI9+zmmbXCxH0fRsW8vntGEtYdGrUVZajV6DvoaXJ9
H/ovmYnq9SULN4BgGsT5wQciESiTEKdbi+kOyT/sfUZN8sx3/M0uqkZ/IMoCnA2VAbZtuep4jJiL
ueIEdmh3vAFp8eEmWuowwPHKInDWttjjCzW3QGwD3klDFP2NMMlW1rgoRf5OuKPmpjqytdTkUb2P
2v3UEYN/3NQCRca+9uGPK/3juGxssIQeDLwR1cz/1edYMSIYIytQY6ADlDa9DGo3cl7beNrwMmKl
Qvclv6AY6kUeKUXQ8ugBeyuJQEgrJKY74PiGTNDiqNiPjkRQzG7SXcQDyAP/uyIVfDfDVjk1/BcF
7faqCAGrY7Ipia8DpBheovw+Vx3bHheodW4OtMRitEiI6k/VZBB5e+ZIH8q+5ZA1KJqMd7hYIMGN
MEntqLq0eYuExNZ9nvjuCia0fhE/1nYNVUrxnObk4cJfu7QDLIdKyiGoOT4R+uy8KLey0SuWPhpQ
Wtxt7VS05gIkxl6vClAtLEE607M6IldwHqgSYpgez8ZMrMg3x2y8gefzgKsZEMwxlXJNB2aKxbUL
vmBhzVwpRLXUuFICYs0WQXoxdCL6eG8IJnrVKbj+I0QJmwcHxq8cqpnGewBbIK160aFPlfrn0CXT
beHnrZePMbBHtWhnRg+dZxbmbO0FD6Yao9cX/YCagyGHLp7AHlk2gVU7To9/CXrJY+CyBZnVpLSQ
c7vnrfRgsBINZHUj1+BTfNCrv2Rjc06GNkS85p7QAkZdOxXBzY2T+HOaJnPEAA6mT15PswdyRDJ+
GRKKof3pNvIItG6Z8pC1/CmXQHVBGIdhWPjbbV+DufUJmkrt7i8NRPTqs0z0h1cFroMR5T7VGH+0
vbd45/u+n1CpzlsN01Oh8nlvS15qLZnO9MJDMMqC4U639+b4PsVu5o9xfiPiZKWDQJ/dK0xJ6QhB
q54Dg4LnEK0aMJRA9aKhIxhi5WAOV6PKsj60GXHzszFc3L/id26JaXH4b7+uzOR4oN/6DJG+U2f5
cj10KoeK7/OehtHygFOAvUfF+HdXECccJ9OunQi2HnpPVw6i3M/x0BQ2BgNu3EsMMVdCGlB+/cNV
jsjqXbpAh3e4WQ0e5AVFAM5vMP30N/8QwNQWFaBLNxk5u8JELKmQy7gDDjxVbDkmjUp8dOgQzqW8
AmihLClp9BvU36JiXezPX16vnxUpB7y6oJpfkDmdmy6Mltq4vSV4n/0rI7Enfox9l2SKwiJ/1unE
wDEPR/SCK1D9Bte/MadcVdJSD7Zac9HfDnYJGCRVteU9kof6FcDjAiWmUqvrlzPTb87bEKlv40EJ
uFr9Kv1/5YcJxKDO4slb1Af6aHjY4uHy1tBuCAqiQwfhWw4KjsxbUtNawQTNzc4gI3I00Hn2+/dk
syS+e9Z2RbNsQyulvL3mhy04XGg+kXX9oOG3Qg8E95fKokJcRfc4rPWd8fxJi3OAsLLtxleMTkws
M00wAbExOoT+RTNnY5cFVm4jyvQPt9mqpZQF6HM2/e171MNqmUpmIEGH9FA9mpVr6uC/gpF90Jcr
FNkdVpxPSD6waeZFlFtbpLtfDoHzLJVSy+pczACoLUWAzBXNG2VdpOk+LSy16jh4NOpqNCw7xTFz
O4Nt5EduZZVA5unwwVOuQIdQjX/D0sHuBxnnXYsEdgEWyaSb43i2Ljq/YSULe8X/XMzscrDEmC/t
iCI731GD1siR6WvBRZLEiHruu7ESK5+l+5bDSF7oesQv4d2vNsChD4qA7nfT30GG1MHZT7t7ZlHV
vDG1vTyzgjcMMqVtTrmixkejxPuEt+6Oaftbb4YzqQuDj90Olnl5d1mh8blN6LUxD4gh/IdhjZLK
DMO1nRgr7dFMl82LiFdqpFw97S3pDZG3D2lHSH/hVoyVihF+zkTXiyIRzW+6sLg2VwmFBodKHKnZ
+9r0Hugs2ksxiRcWyhHgsOEJpzp+X7erbNTFvi0FmyPQ7HSl26V5lybrVLMlnCeMrP9jJ0QmyJe+
w5ekDjgg6dfamezafFN6FQAgQB938oRNnzFrewfaVpooL+PgU8yTYpqemRRSmipl9r4YfUN5caHf
VWuZDV2IY+NwfmJWR4dEznvXWYvGCIv1uaAKmFngn3l+sX/2aoU7HdtkLSTSGvabmGtN5EeHaRmL
Cb8B8kdhFKdQgAI+qP66GVch3NL8FGLswUA4E63V73EknZH92UD88kFZfPQYH10c6H+v0gFhTcoP
T9hHG1oxZ7LPhX3FglWY/LmHJYqK7HNYqjLF/QZ/9bZh5NoW9aJqOF9cpRmEwo/acT4SpyFMfdbF
GFSWBxWRV97+y9xYDPYpVXpJLeEYeQ6Cz3zYLGtdbl4Rpd2khmQSN1iRUgTI2qt9A75K+Z+6NP73
qCO2P4ux27SKi1GytBGgLu+dHmBHmFg+gMfem31ycMXQTxRALNChrSs+Ne2Qi2MVG7W0yVTa5a/W
P+h5DVwbSkNgb7rUKT9WR+J8J2cHYz2GROICQXEmHVVpKTZNzGBFb7TQOoVVoy9Dlw6zFmVPAX4B
naO0wHY7s9UCweeQM5crTrICjZQI2nzXkjU+LrWrqZ7t7w3eAjXJU8pebj7eSybGflVgM/FdAsUz
Cy6ZIhhtnAGpxaxOxkB+VQ8BnSOajffuS5kLjNkI7OXMPCZ312K1vJWu9XbqP4YYEIMsNg+HZGMA
4ksyaqVtTo1SakHy2ooEMdCHg7q3b9qYlvSuipD3zHWT785ry8Y6A1GPyqzlYID35umh/P66NGkP
VO0ENfUo0WeHxBR+dc3vTnQxQgZaC41ZZy3h/m+jAy96Dj0ECW0QRp+6JwVy6thEVMT1fhqUlGaL
ohOgFSTu+GunU75ZbNN2B6mUqdKPCpod/HovaVq5b5G8C33XSP4DJ8u03gmvPZQuDGl8XUuL05iS
WkXukODMk+nNWNdVPTAn8gUQHlsUNg5WQM4IPo88denkMMS5VXGS6uhCTQlfHJcy0Kaew/hDvEeq
0iBavRMSA4lCbO+gE0NG5l7wCgMxH5x2kXAdRT8GiStYIfppAXE0J7HhT3lpQLeAGdqNUkEYe/QT
knNJSLGtvIEGeTt3hx5TxGMHi7pcc4lMsTF94eGigthxd+xJjVa75BSQvmWSWnM1QtoImGClUcby
sEz3R+k6awzr443aawBdlTt/4L8yFQYn77vDaDbaf56jm6R4Yw8+9Ei7XUFijsy9Omzrl2ZDcU+0
I0n30mtDdqGoROxGr2Ln7DHEFNztwOzDPNeBvGZmHC6pYHNfmO29wuoOWPjltoNCqkQC0eZR6N3c
nmUv4stDb68TJ/mDSuEMPvUVLxz9OArgasZQYjGntZV4ydOA0z0D5CjXlDsRl3K0zzaaoE3n/jKn
aR3wcDNk4yx5d363zZsqSsT/tv2hUZG2lqvAInqunz3mM6lOgMy45Jq41d/G9OC+DKW0OJxKopO/
RUdPsal9cqhpzYzpW4LsBZU1LoDRHacdDFMUZD1y8/2LpgWTXobRbR5135KFaDqbShTTliSe708U
ijCnfgTbRBaVp7SkyyO9iVDXjtkEWPBv7t0WzDp+fPD3aujCghsaBAVnsSzCAJ4XXPMS4QqoQA7d
cimcAspqXRFX6PYgdLVJAbrjll9zR7QEI9RnVMMA/e9Jtvari2RMpwJGqi7wALFLedTmVZzcKAoR
FSmCyLRY/nAfLk/Kd7weE3GguMXEF0A/WjI3argpAcLeUYk7AXGkY+USTGlM3cEPKTSzP5ilkPrD
EeoLVyVTAbcJpgaOT2c+SKr4ct2kCfl89Z5gWK3E51S3bk7WnLFBnXFb5M8l6+sLcEMravKSok3K
cr32RJK6zSl7fz5xjypQc3+M3RdDvzjYlfI1UDZH+AjXc0yaOyavdW/6so3DZHlUj5jmAFuQ74SS
84FU/E7iiiwTDzlMB/p+Sxyt34u8Rcz+jz5iEHSyG3/iEhQf2TDCjePMo9wVfDO7TBJDVdYxbcq2
2K7EE03VMPfKR4dV27rfB0M5nc7i3yF0EUfNp2KrdxJoO6dH5uxcF8kSSJwXe31M1aEZ/gCItjni
5wuvFxi0LuQeEpdM0KdEt8XiO2PnwkalptWc1HZYPqD5jeyugpQvM8n2ip4kR/8QTbzBcM9mhEGK
WeVlRib8+95+FujXqLIvJYKRdsA1T/oOFdehIuC+hZZhuMr5tRjPhHgX0RpuwTktYyNbNWRAF26k
MN9vEeueq4F3ktS30E/A0aNow94t9WABo8ERp3em8wkAY/zp60uWOvxaMWJOkuhTBVpkUgi6KIYi
45DLhKrnwVePg/PajpTo7zovG9jx1eRC+kYPTK6Hdhu3gr7QRq3MFRi+ZvKF0b48LKLzphO5x4t5
l2sSEYe0rxkXpbFHS7i/xqw5RhLOTnKP8q+aEZonrrMX8eHfIrEhXZ2n17tI5duZr6RcjTQT6qcu
XY6Gc1YPd/ak3rEYaEG7QNXlgopv+QqtYUZ3hbgeOzP/r0m55S7D5wnh1txzBeZ0e+LbEKLzTSG2
w9v6QqB6ovMzTb5ojX6PcOpXQOiUfJsh/T9nu10ynxFu5rkLeUzfmlem+qDGTtgqTGnO4K6am6wg
okk9hlkrDBG8zN3NswDFa72WMObmscxeTA3CcJhU7xsixUDy7qC8/OE25Unv+x5DMm5xPYmLupvK
BOH3TORo1+5I02yaTQiRv9R40tJnPLjNbWvOBLD0HTxHA1rTyHk/Z6mZfNI7YqrMUajy+dek4ZEM
SrSVsmWrxo1By8pBqpVjZofHMuLVEtg5ZCGX6s4/SDOGgrYllamRyeEdQ3D61a9neNrfmir8lJ5L
Osu7YIvKHSY+/WS8pxYckmwMobhyc2wS4dKV9FfLpIAPcDdatYLxT/A1KrppZx8z/uV2h+uH1gjX
0r4GkPzT4nxd4Gr6LMN1R5RAGyof+QblevOsENE7xLLcXTH92da/BvyOlKjEOFIjNC76siHXVz3v
AURfcoVLw2qegkswQGIERo35jOdQHggwevuCC2c4jBeQR81yRGwEFjiMEgVDhl3zQuVXAQO7u0Lo
fRBH6dQBvhYUo7e6YKsCdghV537BR3nq5NDQsCfxZplkwyWUTRqJwBtpyQFJuDMpSKPvIbUH4mzW
9L0T8ctWTaSMRYyC6Z8bjGP2m3QnxLZMAkoyPCJkkIDg5TsYp73gFMNRy34FvFFodEIEeJ/GId9U
aOYe3svXwmcvgLZjNawhsVLluV0e9mG8l5nqpws7n6NEcfKScce1gR2lbG8G99Hj2pb6cNJNMeb8
Ad9prGyOEiaVzDEo83Ln71xl6tpl75xj78zYiMGXOifaG/8YNnWE4rrPbQfOGEws7D+sZTHcP2/o
Bd993Leo4mgY0fnWgtg7pDFxGNfmYyHgZR/o6Ng+17/yAlFFc7lROM18zOwcggrxWi/I/Fp4mJ/D
JdqZtuFYi6HznphcX4p2/VM0wS3JczeJKok5FkQttCvgBOv57k+PnXnLzuRtjwo/kHNCiTaR7q8C
b3NNJgSDFCIyClTy8Vk93dMx27NeGViYCv8JQZEWssjxlpkzhLL0xj/cyKriTpZZEUvm9nrv/t3N
rkV/hGXbP/kv8rpU+Brgx3A1jKBj1IezuVYGDBgwLFwGXYxjNUCPxhL3xCh6HhwHcTY3umnLIaH4
ZsPdjltTi11NI7IuA2z27nHW00eJZ/CBo/y+hBnG1GZM1nhuag6VCKqaugdyKJaS4Qt5zLxzM0PH
0KOqdHutLEKLomoTTNzmL5M4gIRvbPd4BjyKQfav2dRIbPNtW2MzGcfDFZWR0ZbGHzZnRLmbGWt5
+d9BL18hoFWUEmwZiklinJ+sRX4l6r8yg/4v6oG7zsIwoj1hQRsCqyPFezIss++zuT3ZDgtGAtXj
qkCltPMB0sw7Z6psb/dodekNFtyXuZIaJ45Srh2rH78RZHdUnNG/9chpA/498FYiBEu4NZjsKfln
hLg3I8BlUXjqaeZW4jjBIwTU8WWeqjgDsR7UZgFNRReJDzxtQVYRbBI/OkQEi3g+x/ZAouLdLp83
2NtvVwBB0kZAV9vxZZDKqNj30w6m6UhGma68AJQAvhKDDmRfPaScfwXfi946VVaka06VY3VFLF+F
e0fA114LZVBTBP1qxQtADp8wFLpNBpfNIsa5gJnQ5VCswRYr44FDJSfkr4Afc3u1O3IDHZ5K7qEu
vm2opleajxcGGqxw24y8JntmRPP2jzmZIpZQX05YtrBxRC2bcU4gUcX2QqmT7/ZdQ+cLMKhBQmIo
bzPSP2tng8wagINY5/4Fwz9ivM9Pect5qHh0evBrh3Sj9dWgTXQvyb5Nf/ConLRFPPCQtitggacF
mKiPxqshij0OQFS/IeplM4nQB0eNNkXArnIjNeXA5VAPrayrEYpeXmKjwIC4IzsqV1BXvjrCegUF
YnIr3AlDZrf7z6ALD+yaDUsvf+ONLjqqGW8IrnxRRm8LNmRTsuGK8pxkjr4hBclSGyadmSRSJyVW
fuBmAxC/trdTSLWmk2gd27nDeoifDomqTeep4Cfln160MqIrYj8pwqcwuXXEYTh/Nefrpb3UUdHb
xR752D9CdYQMfT7y73lZ13Zs15y5LqD0ruH6ivrJaj41exKXl95WirhOkdiTldJ3bIV/pupFLu5Z
c09rKjhs9LkiDs9iC5lb6MGE2JHXjVOYbxFEqDBbBSX/tM5PDKcJqB6osxJoi3OhijMnFZKE1nJM
Qj7iIqVDsHTw9Y3QxqZVI89K8aRWOqTmzoOwpuWvzsO+OYkJ/nqLBEF6pI27No7PxNNgpITK4w/3
hiTI6Mc4L1qm4cxz9Xdsr7CAKXCXYLlcMxwAADD/bXH5gGYGbdNdaPFBVitFcoCpwPRgGlEeKoiv
5ZmEMNoB7gaU7VeKsU9kAhFGC+LVHqE7DsPtuCfLh2KkXXqyuEt/v/8A2VGINF0Lmr3AebyOPlu9
1C0Gbv3i/9HrwmLJ77rrxZQFw5KwJ8g3XtdCQmq4U95a6g/6Q8uZosx34in/qXxsNPoLLPJViUZK
89GGvrgkUFbWJUX8pZCKmBeYB744eFN7+YzMHrANVMIzTF1xfC5fwBY0W57sHS2YiN5xNtnBxokG
AlMlU8NnyOEvCyUDVT5241NoD0dF9Z/9t7/FPwn2ugdhYYDmElrO55YeQZkViWIlKfjXUGi1U3di
mf+7lni+oBqC+KFMkpuX1q2ipzTPHV8wgdfFc9O3VPuUduEhcG99G/XkChrurM2pi74hIUjiskIP
qVeVJx3TE9hS1GNXae0Vhr9pPasNu6az2McxPIsQo9uiauJcAWPnhweTQCXs7dvTY3odG6WEr4VE
vq2zm2yEhNDMB7CjOFxkQFC8nPpA62fDexoYq9hDmabpFvTfMPG1CR3HkNQyo9YsgCJR9QW4/t6i
/oSR/FYx8hHEs5iAZySEgYsad2JkpUqshf8bB+HDJWQYl7zGRSVZHulAmX+cLK6bMBqm4+8pFTWM
/tiEw0CbX3kl/jTkKfrgMiVN64N3mO8isYcubWVzqaKW58tEC8FiV29jzj9VTwb4TiezfvdnH9Xf
rJkGSRKOW4TUqFGwsToa8u95YrMG6NKj1xAHFjupwolu37tZXagDZ1ykLPQ2CjL+wUbtmxmtXGGK
fpvZZ/Bp28YEVdE5Vz5Wjb5q7QOUzRfk8dEKE4OgYks8c6yeR7p1ceuWjrH75Qhr8JpFC6u6GwTc
oHkqoT2ssWP/JAZUNx8KQWYSl44HgcFSKhz4zNy160CcM4kd8WmEbN9wQQClka6/NVH/lE1am5L3
6SWPWf+d21c/7XYTHxAi7SqVvqQr2jr33MGXC9nuL4NxRLdM5WZIgqyh7ruOwmpuC8TD8TEcrema
IKADBCigxwvoxDWpVzWq/n+Y7T+tJiiSnKd2iEzh/AtQ1Nfz1yleB2qKYaM/rsJafWoJj/t68hLQ
lWslPef72Z2xkg0dn29BXcHaHOGZaIFP9s1gU8AJ0M4Co1XcIaCZjPwmqxECl/dvU9RSP5TROJ0A
UJLrIeZpK5ITuL4ah4PWuvz9gYaygzp7mrl5Vpi55qWwzY/CYevx+1EdTL2XPNlOcpo8Ypkz389v
dMmda76ppYrUM1HO4i/wtsPqOl6I3UBNGf9Qm4Ny2/QYG1A9NxvAUW1dJ49OHRWsEQ75Ej/IRMmx
II8mGqiZcA4TbjtuhJJ6gbux8B+FfUSKHyoPFgMKTxL9icCPX49fsWD5oQUH0FgDicX/LAKhZhsz
sz6YLPrkOmH14AsraS1LCOfVap72FY+XxFfkypPuCIYqKEIFDLagRPzHpdEs1rrpAsDjaHFE6xun
Wc9Rv8wVLDU/D6qtcybi2KJad1oZZ6nlEp1jXiOlxMsakxJshDl6HrIT24pbVfV4DfLMHz66lB5n
CY+PwpDTZ+N3rq9HiVJYNsP1TRHwjErEU0Y4skzDo5MPY/rEYTq5SQIA2zFS0EZX2B2KA7mD+KOy
kzxJ8sl17zmZrYES4h5bsVw73UX6qTVACSCd1IFJD68gtYkHzvdx7CIEJKq8dJnm75LKurPRboJi
FRWKXvdBZv55QPSfaOq0obw+Mdlb3b40lpohYeC1MOpN5E0m4j1Kc5RjImXtD2UY/sdQBBRoxqhV
2zt/GIC5ys1ZhA8TIDBfbQGjbMnrQAWU3mX6JgqLr1Kxj0J/qqVR7yM1chawSrnhtZ7japypmBGB
ugIis7cQubprHKwh2ZsQ+sn/UwhecRrpwK7FtBaoJYcnmhDZyO/lpoGB1FZkC9/onoG14nMrhjgD
pRR3VtJuoh9OcW3m+7Y8CgVtzQO+iR1w6RUvG6mv0y5c+HNlhiWiw5vykQr9kqtuXc0nuUuWnhXu
uWVlQcz3R52B0a8DDuo6MeMxoE5iMZW7niNZAgdu92bGZe2AMUC6jlF60rL5wE6/T4qo/GTtPzS2
S+aBiPsf3F3reCHf+xae2lYGekWREevOjH879f1Hc+ohhSqWuplpd9TQQhyGi+EorUICWtJAeJ6s
Z/a11YRlVCYI/7Prtoz7ULMcMT/MVSKUGCQbaEs3VH1aGQ8bBp5qaKC0UvUb6c+8JoklzBQ373qT
uquNynTSsZn6oXMiNJEQQn7K7S6ZzZ9acFbySGA5UzgM47KI13aUf/1aSN9blMQEgw3PK/JcJmDh
WurbTh83Jx/w5045ybL6myGNYcS6gAmnwWYbs2+AjOkd3mR+q2nWTBFJ6uGTtuTYaLg3LAajv934
2khrWBjVQsbfSSg+LsmCKt4xRZzmrMTwJ9UpGYrDEYwfAH6ax1mYVvKS4yIrFgmE3sukr7+ytE0L
khc7FiZF/xjqApZMRwhYnU1OADmXDOStxCdvoWcS/N/ksfIjhq1auzOuTBXfqDByw7IFP276r4RD
iha8uKPX54glK919GsR2JnFWwIEKV8NH0/56j89+yFBiJjDs2ICjSl+kZgC+AOUaNh+ZCSrNFeYz
xPjMxWzwbjodJFsaQbEK56zYu/0hBK9UtAggw9TBDwiZx0yFwjjxGeRFbzxG7tvksQqjQRmImgq0
CqyIAcT8y5WEPCl2lQxAxv91u90zhBW7yOHJqc/mxn0q4PvNVElUS6v2dAqfcyv4OIwEVPlkTau2
GaX1RpELD7Bx/sU3hN66X0VHT569AL1+7Uddq4eS39G+O1jpHbY8WwWNu/AXGdLK5HGvNxMGUvLw
untMHajghpCb8nc/goalyeVptnBlB/jB1d75ELyae+SEGsBoRCN/dfgn6Zbz8GSqnkEmTG1mdzl0
y7LE+I4YucsMIhFA1SHLDSjmDcar0hpbuZOTXVxd372bHrV95QpjKvps7kv41Tp33EnJ8F3djWJz
Clor3OarcOmjbgS0Y267vlPKrIEFJi1AGwWZQ/hsubMwfD/pevXhGdrgcxY8Ph9Fje+RXv3cC29A
+KugMXlSZPJ6ooTG60GNnsqw7E7E859n3FTEwjuh7DVFJWp/UkjSEPHcb0FsjpOYQ21iouvoSItM
n3rczOzeooX5p+NtI6rzUkMWIABMrIZtRNMu4c7EFmEUye8eRdYJ8q5MGD67/Min2ANGxrWjNJCN
oEg1p0qPp6Vw4dcErTwXr/rh+W/i+VK7fpWSMj9KdZhnF+ET9EP8vo7tvIu29R+vRNVx8ECcfv+A
JHUUy9UUrjc4+C4bzXsLsJSrrUEU31/qKXyCfJI9bR5BrbBBMPapoA1GXmOiajBfuatAPOCD94Vz
zrMXBjYlaFtwRXvjQTb2jEiLSy58Yub+lBhbTylfBCOAVdwO5Kfyao6qasVJ+/W/7sy7Nl7ifmI4
qzeEeupodsI43OgM6qe7D4IsdZwbphh8adD3MkFfFpKdJqzYKIES1h+MR4hLNwz4QAnaS7cv8X8k
7oK5DxvG88oqVXyxztRsuSqtxLtqIjAzzS08Xv2C29WnN9cHDUTpFWczP+GbkXLSJ1vHI30vrLfy
0duYkRqHwZtnGxpxiqSC4QE/iWystWdqqgagZzofwRzOW6DEK165pxaAIr5VnNmL/TjAun4BiEIY
d37OtZQ2aAJRmSYDTlf+spgjQl9OELVrWL/mG8y+BogZNNhpQGMbTmCwYqL5KNBNdGILr1TGeT5O
b0JFMeyY8RQYCtGQ7HycTpQrMoeMSpdxOmnTSCzWzGxJR8V37edfI7CLy5kXkOEmhtEvF2iI9LGa
UPzpRw/Zi3r2FvltDzThkQhtObXAX5/+Fl3lnILd1mSCRqZhcJqfO+P00MtFdaVWQ629gKVy1b3D
QMbSxyWSoOz41Bln+XKONDWQpziVGmYnEo2el+IzLgcreEvWU1mL4AjFm1cy899JlwjZbyUmbsJY
101nzF/69z3jI6MIEWknqR2P+dxi4+tB9HQHSRplFm/9jl0HRTJpX0GC5mQE0iq2FrbEmTZKQK6B
qkxT1k47jNfh/TCQzixYxKKEaIEsTKo8qkm7F7yV/+KQpdoGxxG7u5cjNfQwWwE6M22b06PU+I2Z
UAV/2GdvIwlb6/SfBPxtFSdKh10qBS+oM0RmCXZWZZnVLuDv6w7WbM29GhcevtXYVQHUCmyX6tz+
KYrvCxFwlWQjXPFbr7SVAQnCvlrfR326TaaCSEOdhdrH9zXnAaEpZJ92mUHMKUDAH0EaLhfjgUJa
6FOeVQ70GMtT4g6bYZ+8xgTZ00zAEarK6yzHFzXGx1p6Eyth58nMgwKQX10RmWvlHWR6YdaZShdK
Vf8wwyqwVseb43a+V/hjO1k/Wcf8MtD3USL0uoBhS/Wuge8gBjwzQOJ/73aXd2miuwePqCs2gMme
M+erSA9J92hBXmMV/deHLE7fcXNKd6vVSIcO6gsIDwz4W7j6cwxPOwvbhuvIhYhPnD55LrXih6Ax
RmwOkl95Tb8Q3hIgB2/b8oNMaeisF8YCy3GG7hkTCBKlbNPyBqlj4XQVdqjaH9Pzb9hj9N6Gv6xp
4zo+JpxZUe3pUp+/RTOC2MuwQRf2G9M/FXXeVMAF01RsbV+dqO3qyRklXGQthzq7V7uVaKOYubJn
dbaTxcX8ldvO4qJRg+w1jUuSaD0MWtXvTTJDvaPPcIoAucxBTFtFkHvwjQu4UKLNTwYczxc1ztcp
ur8oWmx8lC/Gg16JAV9H0WBc34xgw2jn9kgNius7jIa6gBGBidy7YgKiyvpjaCYatgQPRSojdNG8
HYtWWONHU4f4/FW8HxMpxS0sj5Y22mhZjK6QurQGYjCQOTah3l8GMDuQ/iibe2+BndLKsIbkgck2
+0IIf5dkT0ERz63GVrrp8H7xG8RLTVbm0MgQBQ9dPac4iILMAv1Ub84rQnVz3U3SD8y1LEBZr3il
L9LFDrV5XPMCDZvmPqstSr0CjXIyuzt0EQ+tf4GHXADKTnEMz2NL64GRN+Yl8aezohAd728khWJt
UB/pblmIPHC6gPNor/+mDI4zA4KzqedWO6RhtcNUC3nLA1UYsoucCKzmqiP+WsJNHv9guIjJEYYG
/tHJdSSzVCt9eBT7joZ4+supDrVdvdcRoGbeDIPsUHzdPlkihEtG3BCebzzMTKeKZRimvBDSbPjy
8JOMZyhnfBoySJwtcBevOyhvRI/vh7dNWc6TyD0eoL63olkC/in2vNKyqKynP+Jb5lAM/fJ70O/R
rs4WSsomQn2yaANTJZ+HU0FTrC+tSYl5YtiaB2IASYTUYRhDtFyHFUC3wdBsMMyQ+rvuCFqu33Rr
Xf+7G0TIQdiNw1t/Sm5qfK7L37vwnJZabo/1EpVBeM0T0Z5YJ5ZuC/+XfVIBlNTHJ/RQGyWHtkl3
yOtIFKny/Embps7dbnVaMe4DLOgYMpeBTROz47SW9RUiwjmAP4ilFSda9BaJJHtoVrrfuSWM08q7
Bh5Plc9OsPkV2sYe9K4O4009mT5DzeRNAkQ51YRGtDDbWeKKV1UqheLEdkBLDG+ROQq6tufXnq30
pfpTeQxkcuc50tKDf8O7QuZQMzSXJq0XcCyWXU8BhsQch40nQtH/x3kByV2Y11tY5NGVQ2/31V1T
Xz6Ffhy1WI7KGF44OT+9kY+xkHO4VaBczn1D1VHMww5IHwO563RS334/pPmVArW8wrcXs7073TDo
Scq0JdPPnG3OzIUM/InlYETdEA3VkBY9w2uIUXFXkuDOZsRFdZa9r1wE7l+U0OSatlbV7gddn9qV
ZPtjiTw2+6WXw0mjai/6/Uns7P0+nX1S+7W6Wc6lu7JdMvSUwjtDB8guPzPJO2kQEd0RTBa44E3d
BFK/BLEM2MJBqraa+KONNC2IzPskWM/8sLTocgn6X/GrttdP16sC6Zxo3jj098XSaulaeCsVDOrx
421R/l2OO0bE20xCnUp09ppni0CBaMEq52wHbiTh0VwT2z9o99629BtSQwLeyesxoxs7OQ/oYgnP
U7E/h3tdS923XsTic0EU6fShI7sHjWYTvP/UJ697V2WKrQnihtYzm3QQbrQNlUXcLwhxnO3fil5y
g5ZH+Kvu0b2XKsXKSD2DSRMgIu5NFl7icbW0WyLzVqjVTn3gYXARxUlKM8rzwsRehRwf6QrR8GxM
eICBrsMe5FH/7IHJOMtbYPxNN1Z1PWELHySn5wliddQhaOpPhEiBiI19a5aARqeps5E1yF4HbmK2
GrcJHJr3kpxX4GgCQHQNl66yV6DLjttmSvB8Ace4/ggRypl+Y6wbGKSLyqvRnzvpMAt3ETvb8B2T
DrbdQcjnGn0s5GqJsq2zCgYb+ihhF3xXHuZx807R1+ACoicTMHz0zUZ22GzkagA7kYhiN8pNwApb
C6QxSQlnCrLQbSuHVI0Le6jFdmzM0nwgkPLtK6Pr4yCpyE4gIlvdtWxMho5aA2aUX+e1fsZHen76
6o+FIwPXqcy8KyOawtdAvwrU062lC6ty6t7vG5Id5WTp9JRGweOXQ+VcopfsJxhtSdEC7ZPCBHHC
el/MwQkCoPYTL0gXp2KBCBUYuldHMmRF7bRQnp/unIi66sz0H+YO7IaF0DleVwnyJAo8Q1IZ5lUb
d/9Sa0m5FrgWpECzzaKhQ5sA/zX8WXBF95khZZrYarxKfuE0fdzmzF79ncuJ4KeNa6lQ853aYVHi
4LSOhqrTlecBc0BuAfuy31FOPjhz5Nk3WynP1GC/l62fCYX57w3SD5iuS3khEEIsV7bbGEOovmFm
D86ZhXecZP80XwUJySfHOEvmL9JMioCK06OGe9SUxzj44cXClB2Mfr28FVCktnA8UJGhVvAAKPiN
Fli7NIJY15lwlSDv4LBh5dVFqD+K/t12hc6pFYyaey9nV1h3ARr9wqvYCqvNWYuea1RZT0E8PzJh
xaTZyXZw3D/11NMOXAJo1c+ZSzEJTyhq1jWhAAHN9FYtAUvHGHST8a45wKN3u66/r7p2ri3W6zh/
P9LmFlQPfWAwCSGZQlu0Qb7aTW3hHbuZ+tYLE2zwgy5hjY4s5pGmSHFx51b22IpPmbfA1mVBuIrk
O5qdbP+nOUbwdTQknncoFKmyjGHwQVXrbgTSTqDWePuy+4It7zehtRFk2z4+r5u80sU8JuJbJ8kK
Y3R/dIrhTjGNv6GOtwuqkdCXoshBQ0aGsgH0aPNM32AoKNaW4AfNBaSQbLkM8toa4rq1Nt1CgFi3
Woj9qDoo61f9MkCtj30LOYKE7/t3SUSNnDqoX3L4veu2UzSz559zxt0QG4JEzoVMcxTBLYgL/D/a
BSHTY5Qa+FJF0JxvIoEyCsROVR2if/ZuXUvLyrsvc0Cvuzd18A+7jGm/hg3xSMAezX36ghzqBJgD
kBBhksW76kqrvozSCeUvtQ4/ANYiAYUtvO88McgW5MeTtYn4IyUr+K5o2ViEpybEcnRuxQ9EVM3Q
m2L/pUilVcCBlcLZ9iur6akRLCZjwoH+DxN70WYzEkYfyh6wMvStVUIRmsESG4MogVDVkOoKKipB
6vEXail4ot2byBtlw9vQ6DH1BvR5ZyTikw0V5+r7RXJxWzizTxcbEcUuwPc6VzX1xlKv3c1ffRSs
J0PVGQD+PBEa4hGJSc4mdFmJSjRbUSNv7jXsX0iwOCTSQ4NKOz3RSBG6mBB8n3IUClsrdYcz25SL
DtMrUaeGniijdnj7e9o43sp57Xy4kyA7zQZ6taRwlpMfsVEpiEvLBmEcxISR3kP5cg2o2NtgER2l
5GGPfG2gstQAI2H6hVZBtTKQ/P09GwSkqcygjzQySBV9VgsbMWrnxJJhxD16jkJkfwRA+LeV/UIa
iCzBWOVW6h500SCEBT3YxLxp/IvgwcsfDG9x/TqG12QnFpvRXfemh5/7xx+xYvM8xg79lK/uzejq
bPZRixmdrY7yKp0Nsg3ix0hDbV99BF6Hc2QBqRiiOTsEvcJAv0WOUd1lg/eT/9rkbkREnkUPupd6
HLBuBhIW7v/+R7lPXyCVLdkkraCBgJeZrAdo1MJi8pM+WUD3NIh+s3d1whNJIU/ErV0mvZ1Ey7PE
iZ1rCkxPH2xiwyWHyOls9Qm87KklZndcIyvbtlyRrk5Cu9BN8vvuP72MLi05rGUCzXvbEv0UZodA
2gwe55xSSTZlsE6q2ybhUiQ/OTayQ6OEQVvNwvdudSM/X8TUtmyV1sWgarhrQ9pRsaFEezORhK8h
CZAbMKi+8P95BtbwQPzvTJDWQ3d6Vgj5xlJi1N7iWudO8jskcqzMVwGbyBZJev+MsP17+4f6XMcz
gq2k/ap1/X7JjAUy63mm9045LRT75f870vOOWcxjlrxO7FyybrCncekDr9JqPiAd6/zWoM5vQIGP
4GnjAubpOoENn+zf75OkwCKz8rvtT7FTLlKrZeedfzSIKV6u5LebTXqF+BbmUQuuNSiSeG6e3DVT
bX8RbILLw/kjIXGNDtvkxrkxlT/yVDsITCECyskqCR1VlUhU+UqIAkHoxhKLTjZIqHjNZmF53baT
KVIxwOzyQbcftZ+bdXcNiPZ7UV1OkS2in8dVc8aHgkL6ewWt6jgMlGmZ5JX/hKjCoGhO0KSfM4uh
O2Z4mDoslL2CuWx299JtevVSfI0TSekIl+mmFYM1P/nHe681Ui38EDb05fjODvRNJAdif+VYL6OT
xFs/AQ2doz1Azj8zna/vldoGtS7CjizkXxtYXAdPS1IPS/3aOhat+T/3nR4WdG6XLIw1ZixtlA3M
axa3oPU2x3SYxcs+Xcgzx6GSD3GMvAsZmA+kkgKR5L6WQFGoYfLGhSGE4EmeRlxkpQqJNc32yZqU
9arpfiw/9nEMRjzl4BYG+tQn+D+AB1iPZ/jIo30Aq1b6tqzhnsznRRNhJgLxNjwuMX8tH2LSjGRi
dEzIyyN028UeAywEdYTtmneDpARAMzkJADzZWgX6ZpH1qAHq3DpP6yIpc51E4GyO/7hzAt+2i0ZW
ZOgS/DS4LhC29oKpD0378J4M6FD4+KgdMH+GgPbA8+82kxvrO4TmWk7ppMyIFpJwIu4dE8KKavJS
BlZpG7fb48F9YEPbVphd7/fPCKHbAzQc252LSOj4sHj3BQHLqHYO1zs60021JHU+SC7PmrCXQeja
tcDB4+xe4RKP11lpzKUbVGb6hNccAA+5HnnHP5Wl2nv8bQ4I2mzlzPoPIhUrFG80W3u9M1H42qdT
YX3i3lhzHE/NHAHzkJNr1jQdJkwsfmokxtnY3n4f6fIjmKvghWQ9a19kePc2R8+mAu17hAxxNELd
0v2mul1H7pAMzuPSk0pQsrAPiEtjbX8gZX4IVsEl3uU5JJurasYR2OA0Mi6rDV5XW1aHisu1M40M
vqVpzHXDUW7ejXd+Wgh9mc7jFIDlLRv1csCROqDfE9tvtQiQyPfUq4TfGF6nkKcZuSOoedZNY0D5
HMKPYnhEkiOP5kryx/H3geoNCKs7DNQt7nahOt2wQM59U7jLz3mUT+GAORhliysHtIZKQdvJYTfD
bqwFRzf1X1/dUfZ0Nk+SFR8AtnidpqeVgB5QsbKGCx28D/AKPI48RFazHh7PocVlGKVHmqF7XhKb
J/DSis0bI1V73KpCS4ntzBquXWxGpLiSRKh+IVpjJrIBszMVysX9lgkZbt0vhqvPM3yN3rnVLG3e
H/8yHj70kWPyfVWVeQ2OpxfP19RpeMF92JY0NJo8cXmzJamR8yXZaVrmTmoBEHFn/SO8/mZc0vLh
b4mz7FaUZkTGv5UyqJSWUs4WfgeqWAE9tV1DpyBkvciBJ5TxvyOBK9itL7o+KXlWUQuIW1G9HjI2
eJ2mR0i5z47FwbaJWg1flCpBcdWDCVZv0RpciNz6lQPt2f7obh/HLM5MmLj457o6ij4JHc+mYMa4
lHBzUR7KVSWPdZ7FDCryJ0pLU8qQ0LfvAGm9dmFS3IeuVBdn/++7BMiz5ZstHc1PNrDSYvlt3dlx
jcYPpkzP5eGpWGK6xB5t9qFiuckFMm7Q5IpOwR2BX9U4sabRtHEA6ibckQf3ySVVpvPHk1x0SC/1
9Pg/AyN+ruTdrYnKpCJFDadZMxk1iT9CZQS3jsufWQyD1DRmhBGHhcxy+uDoq3n0aG57yeXKIV/O
XolHsEBDK8eMnDGDC52qIeyH8qcoFy5or2+9PRY55+6aL/qBK8mdCXV/KzWOFNsR9zIKJrm51FHz
zuzf1sspv4I1KUcRgo8YLQIXw9HcwXpBMDbEl6Kt+CTzusVxv0ht8mpk4B98QqQTqQ3IxyWMZ+kN
D1wf/OW4euDXELzJQAU+97RFT34pKqqHqGnb39xJ9FBfQf4WtSmJy5mwQxgtSxkMUTNMhtFm0w1W
c5jdJ6I5aHLi/J5rEY7DvFeyt53pWP8SPGaCH1AbdcR+S94aNgdLYo60fp/TMipG5FM9hxe9Udpl
Drq33/caWHU1ZcNrxOJzhZNUH0IpGy5cN0nEk0TlvLrz+t7+mq7aFUXMzwQy4gQip/x/vcNICNb3
ka8gfbEDeCEkFoukpxYj9Zd8hvrNZHi2tDViSzrt6+BkXum6Z9/iGsGPyn4wIavgxuITb6SDoGio
YzCR/DBKVvbDx01EqZ6soFD6bBde/qNbjAiHG8HrYfx7m1ep2xE4FEFaOSuWixyyLZp3SpbhSNfY
di27d7tM1Azx/Dy+oshIa4zsH/KVMuZkS3gy9ri/NKDap06JlqhjzyJAE54coMRnmvtngtVa0ce9
mk3LAL99bPsLdmX7msaWQ2nBI6GUG1X/dfTwPsb9vtunoSQDlSGg+tHKDvQo6oFOr/xEu/gwGtiU
0SQihJHl4MtzAfCyt5aoHgWJKfVc8v7XiZSKOQ3Ab1mWELgnUQBZvBbuDZBnl2yf1bnB1wN9P4BG
Hs9lKiRVyBnocixIRresDbKS+QMjglmIpXoh30joKqNQ4wJ0d1sqL9JYqJWVWkVdjfiaXvXGweud
X41keXRI53ESvZdVAiUz8LuUZ1FtaS9F1nRebjyo0NIBdj7J0QYceg6cKOKAa3b1qymQm07jPqh0
SJLq16a6AvlrAcw4m9/OVKSpnfwJfcDJF7UUu3JZjfpoLjqvS4052ENpRVD3rDaMlYUDQzVQEa8N
/Scb293u/qpdcfNKk5hCub7XI+44sZ6tS6HULS6b79AzVR7dfJLL24paSp8viCMURpeQI2SOCsTW
bUdy/AF9y0wL7XwlicFREOltmWH0FdfsTEvGhSvfAzIKnM2aiidmaVZWyiAbPkgUadCg9W+7bhsy
VWjrnCCTHIdUd/zQ8ZmwnGS0xljLpIqCVOiSWLCFmGuJ7VovQCYluA+gZHpf3TDDotufzeLjw1Vn
GHFBez5/9W5ttiKjDI9clOgiavYzvcBb9OfCvePf8DmPOalPJ6DVnH1yVx3BHTiljPjkD/4iVYHb
EwWuIlZtwDaNeST2luK5ih3zXFCH5bJUMLdW1y5FTU8ds1/RS2bkJny52R2/vNy9uw1rxSFgJdxi
Ps5ONJgRCqwvGv9ywmfJ0Hk7Ub4kJuiLVhRCNWG23SffJZSql0uqiUyFLviccOsFCzOnvcb/OWtV
IJUEk0JmtaPiHMQMUuDlqtCnvL+Wl7s9+OU82BM/yOHetSuUBeqCuCNRhuWWME1XmWxEHE3dd9iU
6RzpmWxvTKI93DvVQGtAeojd0gAFbJl8qqkAJ9C/SQzGyP8DpClHTZrojAOlrxnmzX/dGhf24vh1
A3Yu1zvjNGK5NhVR2kzzeRFBxUIcroJ4fWXGIGue3DwO7ggwTR6/Gn17Swpn/KybeC15RDjEx1WF
VNu2G9akYSwTIBVFOXQr7MI9baZpwoa1RNetTogheoTZJHtiBWF5EccHUF0ExXSe7WoiZpDoG9iq
LuywXMdX05n7n4MPDogt1Gcc9ntRG84LlwSlLWRTLCZZEDym1mFoshRo3PUkL77gj3c63Wz/JirH
8PVZPlzFBlo+4U3iHsb8MAz81uAF5V4+33Sx5tOV0t+WfSNyEqmmxz/jIgQJjLungUYupYAfABTh
g8WXgjsSuSL6VfnXOqM8MQ4FzCw8/MWT4qvqN8lu7C3FNNf7bS7jQmDr74V6Lg5ysNl1kMu/eDeT
ZLukB5CBiMX6AADfAlMYnbFpyzq6dg6o1p9KgEevbvoi+S4pvKi5WTXhTUB6nroa3gTRsSfcgj/L
ziB2yTv8nELy3tP5iPdoD6f+SPvZFMKEGERR2AafYt0sWLLZqf9wDL0IfImDxijjCOyd4VJ0QET9
Qw9GaSDqQJz4ByYzRAc1+8zhm/jKcCgl908sRhYHCqkUEvWmCwRVUEBH65UEEFdOJiqVTTOJCzn6
WGFVWKK6HN2/VLp8IFD+hlGE4E94maNizmSuPn3EKslpxOMMz0pPI75z5OaGWyS0OAqMUUJ0eRNJ
BUJjYXUpzFASuH207z5Icc85WIP5Mjt19R819aBieA+9rwJV1q8HV3rJU/XH4394UFCSvNeaO5/d
6iK2NWWfTNlmFOiOP+aTber2zBUiuSSFmlk5fu2Q2Pe07Gg6tpxRlwBgmvPgSBTZPA25CiAla+wa
H+CDBQ6TdjakZROmN9WLJOHHbahmjMGkcNAzcNNTD+o+wEdY+kotfmDYpMffBVAWALoabL+B2bvs
1bkevs8Lg3WC141K20sdphOcwZRoqYfs8ihtGyjbk+SveHfFG1uj1yJaK3Ta0ORrlbUaeVop5Fuy
qFJrDPdm+xV+nm22QwK89/SwT/f6Eaw2D9i6i7O33Nd07TJQQEs7jzpwn6rdjpGROIUy5EjDAscp
KbXOfFqWzDnJIzWqO9W+BzKUCkm+5jWJDiZbwGVJI5VUNadurdc4GsomO1c79NThWgUlj/A89Aoq
f2EYX5jwrd7JHN/jt/q6sgc+Sv4QmyiX1ujVMZHJrMkf/q6WBgcLhzVbK5QAZ8r/El/3f03PNNmw
bVb7ws8vRzFtFH+gXcJmei3sMEvrlgqywZnlrZgZ82vX+5/ibFiuaguPkfVGkJA6KyKkmjDywNC4
1JfrB0QTVC6DWrCFYdERF5MOq+2P88HCZnJvpzJmEvNosXMnV2hEYHl6WBWt27osiXK0fsw4M2tb
0v5JcJPR1TZieUXZKuMe6MYluXG0oM+BPF9E6HOAlCE39blZAMeRzQfwbLUlDZykfr8lBefcqdGF
Avm+lBsJLfGfjKHuCzlYnznt1cl7TlKwLwYioHQqNLmkoAa6VCYyXAWlqRTFssTvdJWhGS4EeoyJ
gqsEtaFNEP9Z/MJmpmeaBB+Ny3Osg+ILFbcNXNdDOYk7e+PFWGDwTwOq9PUqEXUM5pITE/Kar2Nm
UF25k4O5wPtRaSP1lq44fVaRy3RnnY0qKs1FqR40ekgU5QM/5hxSLNZDABGm9ErCN5Edwcap91xa
3m6CoQVqWVAKXnNonsyFnR42CynuTh1iX3MwWZjU6qFTfTfIXLNL4GNul8TRJaGfJJsR9HXiZdnA
kbb2SnOIt/d/LX2X1kgjiTGpF8CWz0fQe5il59G/2mH1Scxu3T5xkbX6U9NmqeGZKZLuEaayDdds
MTUDYENsx0pm4f39ID6BpzVaePyrNx3cRn8fGHAiD9STm7cXYnGMq4xhXQ6d5qJnWFsxPxFHTjnL
D0eb20f8ShNV8sb4XAQvLVd3E83PusDcxTbt1O4ZGTV+5S+j8OsAMGzIkvPFibLZQhC+LjqqvmIA
iOKBRO5s+sQiEk3NqbWI55bSEvJuNeOZk7GJqiX6Dpn6MzB0Sih/PdnqrAURWJsTztX8Dy/aW9i1
rc+4POPhGs32JUTZJ1fmuVxNdlGHsU5Q4gRHiCKwqa/MJ99F+Xne1aoX9PsclU58BPMmt+VfDHvf
mnTPY/MKUc5MckxzLl/sK/Ow1/hZQJBQujfTpmw1iAMGGzwV0xEyNBsWqvRguKEw29q7zVhVPOS0
RLdqCLdfZ37VAvp4OI2w6a2L9KYbvapdAm9deuPrY7Vohw3pTa8XzOBKFPCIzpj7jBSkBR3GvVzu
fZQDFRqQh6E6IyE6eZrpYSG3Nyv+y6/11D1UsLSmJ3gHJ/40bwHDJuO+dtiUZ7YpUm92rn5F/h+u
xaro5I/33r8JNoWuqVjuDC4N5v6THbRpeBvGDQWGYA/XEr5RN7b4YYQeGtHRArPi3g2Gy5e0lU0y
IBo6Ys4QqzbVvV2Py+nPNOdG0+9eyqVBQ0by+ApeCRH/Pi5QvUXu04R3ufAz8D1NJDEKDIGD3Zqe
h4Xw/khV28hzal4C+ABGq14T5fn4YgOMGFcTZ1cRuIb/BhNOdq0GxBL1fk4p17k6LnokZfu/7CI4
0y9qj/undMyGCidaR1fkmsknZkvpF5yihN1l4Q6H42JwnBWHDS9wDifhZ3cksftXmZgH8yO3iTPn
O82W65wvLJ7X2uSauf6hMO08RlBIRSCQrItwQNgNWoavU5zR44vWjs4nrp/11EzhIg2WSAlAhICa
jEk7LNJcv5PjLidHcc69/t32hSXq5t7cjBkhMuU5yGtr0WQa1bjoKgqbheae3HtlDilW/nIvNlo/
SXVJDNTArRYV5kfXI6WikGbl/lGNGHu6FsoptqHfYO9Qlu/LjUpGvs/VIqkMJ22UT6Lk3n/yFVOo
4GXVyG1dsgIdr1Xd/l3UUTgIVxUUJRktRwx5wka4fVpL0QMgQH4i/7S9Z/aXh7UZmnJJ2DZroNxb
9FJDOOZ80BguBfjKYPVpZxDh31W1QuIVzISIoQ/wTRTUP4pwgWB5lKDNtr9WP/Tgsbt3A5fVItrd
M2XnqpxUKaa5dTJTCzX7gW5OnHTQwDgsVlmJ+kvCglP2xBk6tTubsiTpHGrbj//M+xISV0A9tiaC
VxcmLN6GyWSS3yLkdtoZq8bwnjiDo3Z26dwZZCc1Q1WrQViEoQltvtlPrxALOW4UbGJYxZLsl7lx
7MGvMAkb4AfRwplNRvpL0czrD9heWH10bLf5C0ld5yG3qL6zV31rTuPDEC/FYjZByrB6MYjwzcXC
l9XElcCnQzajg+z4m1BxntgTH0wCxPLJDlZZfvWbP6NAFBzXeQTbQzBZo4DRzMo34V5CpJKZTFI6
97aXE7+HsgQpjxyVxwx20xZYLeD7o226j1oFsw6TPd9Y1ofLQ/PpH1w1UgseT3ZpLKCObd1xbfwE
cX4CiOydKxg8etoRLwixtfSOKZZzRjHHu0XXpKyADQHXS3FMpzg5QKpC5OFrUurG3gOFcZlMf4/J
a119QEJig+XEWGcLH2/RWnzy0wu3+MapH9Xc+s/aqvt1xrpDhrIZkE6/EM7QPkNeJjGVtM0ZSxK+
z5CeX5w23jimAJgHzRVz4ZyHU2/Ys8MXT/CazVfnAT6LvI1ZuPWIgKyXOWiorrs7JA92khivWNwo
Ed0ezDzscPIsUZolmhLFDep4IZu0Lua2Kov0XgGU0lQXajlBocxrmu8XnOZO7DkazFTJxt34nt0C
0kxZB2yAloQIw0mXVTfGp5lYzkjKUv/ygg+HlCoT7VQUgcnfAQ6cnhqZW1dSIjw+hArVaFkfNAFq
lh9xvuueYMeURDx6Xr/EPhkDRRvjdGY1hz2vwzPrSYHrAiJuoRtO38d79zxQBUVIXGbIlNdX95E9
tCiplygOlTY7nkqfizec53XvjAv4DARKhtDi18QXu14yNKawqDpL9c0S7Vr5fvRJeIUxHUNj3dDA
zLwttGi+b06v1aVJ0b5zjZ0Yrz5RrOohunG4O9RryeBP663dRRo/V5S909twUe7LgA+arxJd2x8k
2xgo/2wpNQ0Nb805CWO3ySKROQDvj3sFwjDkCa3jr+Y6E5FCVrLsqIIplO9h7CLgtmER5GkgVrYe
ov5MU7n08tlCgeuCkzE1/2AFTTdypuyE7e6kDWhw6OFzwAVvfwCoCfYZ5u6WWna1+nYeo+AO8dV9
mtqxdpcnMH1f529rNlBAoyKOif/7r96Xia7thoDC0PceFcrZEngcIuYhd/Guk7hOb0uhEr5gwryT
MIW+mnZA0alq02V6+i29yVYNkbNORX8jErIu3Bcge8ETU52itcns7Wf/9HMtbF594QZzgCkJtFr4
wjGQ5L1ZoKl2UfYEWE9RFK02hlx/EHo0BfgkvcY2jUeTtjCrqcceGCN+zRKw0xb237EU9eD70v6F
b8VlBaGX9O6ZC+vNqDDRznOaz9MthxvIhOPmwOj4QRTV8qMpqDBl+N+MOe0UjOymswHyrc5LRsYL
Z0QLYU/LqJK8FWAy2lyxFfmZnp+7dfNyoqvkdg1Z40o2VlsVjOLcknMERMf3LCA9DpmutBsJqFYP
LqhA2kEAKBy0QG1QMJ9O2gjzP+06HwoOh0I+8r6uAWRieUVlZ9xtR+Vpu2Za1tUVjyFP1ELeMmMX
V1k8nOm2+83qHnxs+vwJoYl+hw175ALtjhRjikynI3RB1Ny6t5xPiu6FJ1nniZrIDxEIYxZuHxi4
wN5XyGqcsaN95erNMQeDX0qZfqOmkAxTWfLGacRu0XsvBXzfqREHqRdMdaxVB4/00S+EHHIYlOlT
dGNNMx8TNEMEoywp7A1K7zAyRxIrorH+IPGa9RWD8eaGgLC6KyU1AkyeYEeXRGqYSoUg8uE2b9BP
14N3SG0XxiQFfArQnlSCjdqDUWlAHkOQslgLQ+w+mXo5kQ0J3IcSvMjjwYI3H48/xrKob4/5UHnl
MGb6KOYZ0GE7WmYmfPB1Zg2Z0752CV8/oqgqfrYpahCo1F476qkxVytOozSyMuX/OdFXCuvmT+SU
Q4sbc+wtVBopJcosqVXFfj6G4AH/kR70DVJjNfa5Y66Cb9Vo6aOZX5gxn+PgFdPIpARJZR+U55mw
U5FZmkCTZhg9v0NlaaQsnSBcUc3zMjib4abaJxZQsgDhEVIVOaunsDUx8XeaMGrOjZ82JNgkMO4F
50Fd+ELTojd+aAaV/6hiH3teT6+vl67HrO94adPWiGPNECLxIqDfcMdprat8WBDxDmJ4uYqfm1Lx
4Setb1XnhnS/5AE7ovcXT/Bo9OLLyYo5/2TvuengFEMvShBHwSAUkmbJaR4tU4F3fdAM22UaCWuN
af58xdOmSQ68IKWcpjGlq8J6lz5BRcWwO3RnA7cp51V7F/td6lXwFUhhfKKM7QSCdSqlgJaLiXUJ
jJfuMrELEVivYsGS5ivNONeTiS2dPOsgOILXYOPopQmXI0TsrnS8OGMPsRhTtDje3ZH6QkcJ3ugo
rhOgdqY/lEa2HD8p+QQ6DHDWH2yj9+z2yj5CKfnLN9OGRdsdknPnGexVwI67xQVcuYC+x17mUcbh
bX5rRDoKdgczyzEjv2PTAzlAIgin87tEtnGozalfzAjrh648jK5XwivNBtvbuNuDYy/qiOF/RFrA
YDwzu6DP1Rx5H0B8FzcNl4CkIv85MqQfVoxV1DVOv/OWSgdyXRmI8nP9Ca1Cdb5mIlZUxQqf/6qL
9FB/FurpESXjfq6twSM+FKXbBekSKrK3Msl8Eoos9WPNM2lIPBEnt2ZJraPEuycMjjquXmJiI72t
11ObCWnZ9EH2fDdW/f089QVdOLvRwmS002I6VG5d0r1qSqAHt72ad/kAGdiWy8OXhQ5F9vtXZd6F
ltxfImDiLBRV9aD3R4CPakIoGaLM9Fnvuupnahvl4oe09nipyfL5BnKcLOhgFjrm8GoavPhXlwUY
t1E1pXddO6+N9Zc4M03xuLG+xzcNaBR0IZt1wdcYSiUgtUveWsBMFnKxKy3zbi1aEMMZn9lZFiEM
E35AngRT3cfAvIk3snNWZ3y6VfNqMjrUf129WUszffrXRKh64SihBaxWj0I7coY52RVevDdmlLr7
Vj/8U9DaYVqP09LnHCDEUInGvT6SsYW2zQe7QA19LNvQSSNGml+hDgU75kwQk+wz6rIy2Fgx5LgY
CEt3fwIFsXW8pI781qXo8AUfun8L38kRF+a72dfeLuYQjr39WmlalcxngqxKjaImESzWhfOKgPco
IURytL67l1h9cnoylksAZGWdlwQXbbuvqp2tW1K2o3ZPSNGztCLCfdkWtIsSzPkiNFVdeu8tjS6I
aQzHlnkUlnjcX/t+iqYN6h40Bpt2XCKk5iartDq88tQPDDu3wer1kMm9KGljX4NPUJQ2FMPx4pM7
MPyUaROr6XixmoRb4jPJr3ZopcwPnvTWpdpQ0Dfq6xuwueIz65IC/3iWkMBQg2Co5MUm8vZbWICg
mSW5zFDezM0nU+88uepPPd3H/nrg70CacMG1E6NG8z/3rK7x00nFOweN1XtnMemvN/wBfdfO8R5I
m6LLo41l6xLZ010K7FcczFYJ7eNbdEVBPMlTyDGKq7j5h70qLYwIuAu/unaAEki8jmao5YYZYN2v
54IFKix30DU6JvH7bfBUnr7byvbqdZD2TfBjPast/upV83MRqn1s43gxwFyKc6A//NzLK06B3Z2j
69Zsdj8xHSASYq5T3VWoVoEhLfx43hZponGKmhHqOFEGPZLUVVRG8mV6YjsrIwaDOL4G6vwaS4F/
goS/qEjUA/n9Lo3CuSaEhw4yvMl+2Axesg8mUlbys6ZN1nv7K0NbUK+7bWlBjQXqWFnDieCSMbXR
JWPhIG/hABhtDMujxylaPbOYbEmytlhGF1tBoTWIUFI5JDBko/b1ezJ3uKh3gNv20iAubPme2yYH
6Uy6f5jhVGumnRThWe8RQThE7BoU0WKlqNzjeVMFyT7tf34uLFtezXDMxxQyMPfDDdaXi+k7Znq8
VTD+2kD8oARkA+WbjOl05MRiTFt6zeDP25IRdCVyhC0nP4EGo+hcVMOxwxZo/hKmBHiyPDlsl7eZ
br8+z6OjpB/llnoVJQ8Ur7uMr3DC2sewu9GxpQZ+Q6uBYJWLzX3K7JjHgzmlOQBUQSpfBULw0qih
sRqVt8oAsEOxXUvYIttX7A9rOmStNHDMac0YhMU7Q/Fc04w/IDhyigu7co6nIwIHaEPRi6SHuXB0
4JrVzGHfSBGgRB15cjxMIAWiqveE4N8JJIeriWXQihcol/++pjCxSjZMeNV2RgfuI+p8q2srW42n
qwUv+4DgJz3ZllSvEiW6BtgQJEod4MfaMc3j44qcW9J5jf4F+EGt6gIAGx16C0EWeQ+lAHkx2dXu
cv0eQ9gOKnGZf7b8NZCG6ukgJUrD9gzXvY1C4cLBwGmXDJpNdAObEeMBWjis64jo8eBvqdnQv6M1
oPXEfLjawDDYJHqwxKFYg3bW5Ph92ljjX4PFVLt/DQeDF0Wy/XWHFZJhJ6hfAPQivPL1YHSrYLIB
DjrOBDdAYdHQOqnRV13ni7XdxAcerNXHySyVCJZ1ZEvaCEyfltEULIr5oO2cV08XB4loo9G0/nmf
oph8eaDka/wgSrY0fYHY9Hjh/EjCqEA5K7WQ+Q9XyojriGXt+u5Vil2XekGEEi2eAGSuVLQK0MtB
sAj9C4ZBMFOfrMP3aIraTJLt+rhXSegvFood+khRrb78shFx0i/IOj+2rqERyGfjjrSOcCLy12+M
K1JFmeof6ykiY7hbfx7yzZD3AlEu9fk/pO0QwKIr/olCghKz9bljlaAqu9ZvwQTYtRMtqUdok6qw
UvzagHKCK4O9BIuQQdHSK+e6lBW1JeXM8wE7Mw3qvTH7e5msNd7nl6e6pcT77IPaEaZCNNN+fiGZ
38MukvvMlglHA8fzwiPCEgh2lJNGimQQHoouO5bpLiaUMSlIy0FzLz/h37WNwcVoxiGAPHjWf+lP
WVrBe/9eW8lCY7Iczb9LyMj3KnfBh87K1yLFDQsq0FnvZd/CZKWdh5/2PpIX95Vn8SVjSPKnT2/Z
M9RxwYdOCr5nZmGAaIoDVZZUlo+E/CecilRIsgQMan4Rg7gkhqlC5zoTewqGyLUziGP7aJugyQmY
QuXF0YQXw7tZHtJtoNJdTpbhpbV3f2NSyJrA/gpLHhkEaKLqnOIyxsgw2EggSwR+EqUSRpe9nunC
sUU65QbAHMo1p1MIL+P+9h6gLBBy9bPORUvvYK2bKwRFnMkxDl5eveuEM+1HjvoSnD0FZmlE4ofa
3P5jivB697kqXCKTPhX9+NdkJTvUjt2XB6ZNMmizlo8ujSbyCea4tIL9jB1b9UUvZXDlau4ZZhQ7
RuznCl/rKSZNaub2CaJOau7WFZ8gECb+PandOSVg1HsuU2fC/hRmDEl21ASA1SEalCS/ZNZyrVjA
Na0C0QrcebPW6GkAiMUEKXwANueXFC3f2BRq1PYmf/w+L48VTyavbRlAJ38UW+b5jlcobWPJt/D/
pztmJn6dGMczXT4tAyK1RcwCgydmmqJKxvGVLncjAwDYhRujwDtjBOTkMFmNctHPVtTrABrE1y3z
5CXBb1xXjvhx1FveZ9o26q5k+55hTBdh+CMuMD3YqjBLTuYm89a0EZionAA9k4T0W95YMf3ZC3cK
EMuWTYJpTlz5hyh2b6hKPPlKr+uSMxyoKXYnPYDZyhYj+uSzhlh+wdo37jckj0k8pO4F13te3kAC
zYBhYD/Epp+DYxMdTzuMHw7fOt32/rhPoCkSf0Z8blnQaMdnwZOOmMh5a5A03t6A/KT3ghN8Mr2W
N98nvF0hpKp9c6haiTrlGHYyzbux4jMQ6eTMc9a6tX2RTnvfq9vWX2nC+JdLli00V1dKaUu7K5Az
HT89u4KSzHJAVR7KkkwLIrc5n9D3nFPBsjxepeng7D2w+CDSCB4W4WLB+WsnZkgaZq+qHjLquuT8
RmIh1vMa2lf1LabDnoIsqxhnIrhjU5Bx0k8afZsFdSHnlNlIHVrrl7IN50dwRLxvMQcTCx5nR4i2
84CYSmXiy2HgoXPGPjtnwz8SOOV6qWhqsgXtMfjn7WZ7APbbK3yoU1dC9Cs/wvXz786QUH4d1tpt
UrR0Zo+Q3hJQ/HJeUz/2gz+1wdrF5CXoURgFU87Sd4omuHRbC5Ap756vMsr6hSITOZtxgEIEdN8K
IlqYAaUUoXsyI6YkUtrDoGSuBde5b0csQbm0EHA6Y/Rzrini7UiRFfUlPWEG9ARqP8YcSN7ui13v
CRwCXr7+hzs1psE+aRPvoqGKqTXUiz8GstrlAdezZ63d78NbIy5J6OcexRi6m4S1aTM/23eYNdc4
PVW/3mD0exOcVCwRO1+3djAGdvtSWwH/cc9rGR1S7nLjMfVpU6wmVdc6SwmRdXZ+mHE/z34SCHaD
E8iX+pfGMJDqb8x6P2UfPsVIRFzBHrLgIh27lRJu0cBjT8mAonCWE/5puGvOlslZwFqe30sOQxTQ
HDMpJy+icnX/VcV1CmA4KwFBOQq7P+xbIsMlfifMCqi5OlmMaSA6RDrsNzw7B86ZNZBNMTCVwrkF
JPvkrhmHbA8i5XwiBPni/SSuvyH2i1DsUyweAJ6sF8hz/Yq0rCSw0vOiv6fNQyxMKePePIWPpJ0j
hXx0aEJZWzNoTMCaPLHZgm+K+JW+yo/99vkWfNZtT0vk37baaVCifFI7lnffRBha5ub5Oa13B72P
kDrcwmvJizztZaAuu40cI8VE2/yHE+KhI7cn5MgXTJZdt8o+Z/YjZrZdJTr2+ZA5DmCzY3T4cLbG
qdweHOsLDn+VXjDsmTAZwA/WsTaje6mVVcLPQZxtahiCo1BGewHXI2dc+yHfhxZjMpsx1HLl9AL+
hWcdQ/fdofKaHBRn2BrmiTZpW1VErnY20s+4z57b7mmGPs9q+oUzIXUwMjqgMfWPVr4gtH17Dvrc
CPE7Ov68couUOzGDhR51yHHqFLaUao9IpeA9sPjV7XwuhqnI+0y1L5/6Gwifds8Fkt0cvh4IVWLj
xx/UXODnvmRi9KoUaEYkxPXspuhVAoPWJhP/vAJHSjqfqUTZbdtlnDpsvmFhwUEGdcfV+Ir44ZI4
7pTqUVVihDYbi2hW14mVlRgfNoOTa78iQlySTQLEbae4EKxNKVDGpxxwyscj0fP1Ix8chF2pcW2s
+UHCdm5gHiU0gWjySGp/i4w6p5OTh9CE9/hkLSVeQz7g27IaIN0gTDiwUu4v5ksgg4mSP3uwiCDW
l6jXkctOfkzflRiPaBNqdQ7rP0G3wux4hQcvPK0BMe48o9EWEAt0NEVA9ZUHC+4TUAxU0+1Gpzwv
Z3xPxwaC2VoLiiUoNnus/ZXb3l5wxaoH/LiHS4bfscZkX/Gvb5ag8mvCe9Lo//uuJetUAMmPfWd4
TTV1EVmHlqQt2NJLO1MT1eV4VzKXhbrha77G9PJNFRtp7puDeJitaRTsDG2u/uuNRnhM5aBWfMNX
g5FueRrd75UfcBsxBWArTPi0+zZ9wNgN11ebvse3GxvRigBcRnd6rnWtIPGHh87cNBYmwSCvSCb9
7mTFGT7F3cZk8Socodxm6iZPuGU96g+yHLw+czK+xadH+rP3SlQSyGZlDMCqjxn57XlOFJdyS1g9
PIfmb58HgdPSJBSRvJRMIw2YTf6qoRcwfBjO0o8QMKWB0V9Exo29UaR2SKJpb529DbVFyXtmTPST
Tjv5+79YYb87NSQu73mcji9/EKlWCYbpV6IsiM3py4RD/Vk7cD/X8FKLxXPIhhZDx/HJSEoS6ZX1
7bZIpCkKxm6QMWy62ToF3pEyYZrx1PXW5WLvIum/NX4mDwhdzfXQ7bdkdwEBlYFyXUwP28RAKwT6
d7GgIH8zayVPjp2WxCdRqlVvE6C9nSlU/v4uC79dIliTwhlH7uOfu3rV1Rph4EGfcC6EMdP01DAr
qXUimYZK7Ct5IHvG+jdiKB9BwyV6YegY2wSgzB6S0n8E2eWs8goeDMBPWSFw03h01pU54+/Qs52e
3VbjYFrgzOrKVU0RN7X8ik7BblFFbkBGUubBpdploXycm4RD/5P28oIVLi99TeJZT3+UFivQITot
63LBvd6a22c3L47ochBNGAjIc3gKhTPcvrc5/LBbNWcyj/qq/mY6nVvq9ofkSuC0sljEki8/7Fvf
NDkwPxcNoVyqij1qbMI+RpifbBD6q1tDxspQUeeYvJXc5G5sIlo0wJJZ/4UFkKmibyt2KIsKpIaU
6YIKceTIAmkfomFW24padYGat2a2WHQ9h46WlbIn9Q3bVryHvbX0AnUE1WfPZV3Qcn85TgXhwMS8
VmwDPC79u3SjRh1VB54Vpx3EMuniWZTLjpydLUtqPJgPSzcaNNj9EbMsrHR5h4wPh4yEkQOtyOq0
J0cMheW90lW8OccEsGkL4+BFQF/riEH+gylK6Q+zKbL3iTNbfL8GYlo+y8bhcesKE8A0VrFFGmmw
FJ3FVasvMwkap/o2RKGmgL/lJd3egsQDCsNgBhz64zULJyyBwyCWoHxvfB7Vj4rd1L3W+kYccQyk
I9SDjU5IIgfKrCC2W0pnF/ca2cgqXX5uamIflVptOx4tk0rs84zGScOxmD2RAx49KxanCHmhEJy8
8sitfHr5XAhbzg+Ll3h/0Ltri9Bfa/nGcuYnbqBkclkuckMJOq0fPtBBGbeAl/bAgan4jQl8Uc+U
oNYVvYmbNMHLAyxsIhzUIxucMumPN5lsbk1IWe/LrLGeVDzg+/uuZoSPznw25UJiKu4mSLcGiuhm
5aN4ts/ibC577LywhR7yC7bUaM6MibNzVvwFOdeM5Pt11dJ03RtvCTHaoxGgRNIv0vG3o2QK3rWw
ciSxNTFBkdKJyUEjj8nFGdjfU/oPmQblHNOET7gAfZwT0caYdFXFj1sblQi+8T0O5VzwS+hF1nA5
+oOqKLBxtAxIn8dbdTr4TUcrS9ehbPBFQAs3u7rYRLmnTwUq4X9i4khSHuG7d+VHhCx+VvS+c5Sa
OF8XxgaOKFZk3wgiuUFjZ7uBcDxDgTq7ZOdJu7LOp8zvUWqAgJ5Y795LabwSc1YIxu1tLpWO0kQl
N5cOp61hUu96cpSICTDUCJeSazfeQsog3wp+Your208TmR2htcV9QIMw+Ir6XoHd8HQOhQ9fRzRd
uKt4w3TaATbyWmDBXzlytRsNtVfx2+CeIpbNuCLC1WjWXPDjtVBTOtrSiO91V27Nm39GVaOHRxVo
ZdioWppjfxQp3NDBpFtYirNhkxZ60ytPlOWHWfnviCCg7U0Jm3I0DyEG3oAEKBcqyYdJ2ILZZDD7
3gdc8U52kq9JyootuC5/dwWBFlLUIdkl6MwC6riQNbL+ghgEhgdsHc6v4oLNPl95rpoPkXjWjx9m
sS3qnFhQp9TvPPHRQf1plnyM3hQppsVJFqG3UL/uHTROXuCQqoN6PhL8MMCGFS5CHdK+QTvl+574
uaQGFcVT6i2gl2loRmCQ9oJONA2m5o2mukGc9kxSiapDIb881JtSlUA8gae6lbTUlt+npnefuOcY
oUwgg6Y4I5cnn5p9ctN0qsJMqBpYFl09JZPCDECFBm47P1cqoxbt0kTw5hYrcjX4LpNu9l9jUXqg
cKlYq7gUW4qqdy3lcJOjqw9GUCasn1Gb8j1kx74eGOt9v5IZVJoxVDo4WabYDWX06gaDoGyCzoxn
SPj6MXv45ZjEm8SLnNK+E4p5fuorwyKexyfUW4CVgNFpxu/ms5iMLF0CapCxyjXWIqkL3HvRTK7X
yyhI4tWWaK/AgoFn3dGCyn3Zx3jm2GHVYCiZpcm/mwgRuNgFAHYeojqlxtrZs9R+PCUDki1eOJwx
e/p00PSbVv9uIgZAeYQUEldNQsSMK3jqxAmHe3Bqu9tGcZaTQuPMOsOJzHEB6NCfnGkgrAOxJoqn
4ugBWG3fmu9tLDzW0eyF/y2VAilYm0SRhsUfFq5kTBEDdGLlKiwZJJQD2bLPRADVZwG6q8B2TEZ7
Tjc7ez1/UDdFQgZg/V9H+JBg0tWj8yjrc1RRYMiGGlr8nQoTU2ucd2D8dTcquuv7aD1E/TeA1BdV
j3Be7K4EWrd67iK7zAMwyl0z7NBqSSQPCm5QXpk1AiQN8O9KgEM7+5+1JV6UxXAg9HEYHI+wySt6
Bf5wvwxWWtSSIk9F0skpewpaKp3MVhCHOCeeIl2ymgHDUPsiQd4xxzRqe0zQROSh7wbk/fmZfLCi
EIb1KfV64tUOZRgSzp4KTZ2qigC8D9OUu9KJ21UD0aVGs1I6o7rig7iCuh8+cL/oVlfnOFnNxTKa
FQ1gGjerbJ6hKgE/DwxS0ND8m+BdczYiVhr/D6u+jjkEYo7QVpezK10/UnbRGbQH/n/7yMzx5icE
bS8WT/meBHWeNX4zs6w+VOTgCQdIgKqexXxeeY7c8i+4zfJoWiEd+jmicWCouCBbKyYY95W91uD8
6MqpkmpBmfhhM7scTEl0n6SKt3mAEUAyK/e9XNEsGiG2GwrecVdwqppQH9JvThQn9aYr9+S9LiVw
EMiY3vIsT9PchGd6ClxO84M28WwwR9DwTMen/1eWVD+fEHO7/WQmPeRGqF0Zf9c2hHslnREXOheL
iuVF/EfWmpjKPmOGoxo7E+KzdOrxxQXNRdy8x27ja0Y64lIyefmDEuHa8mrDM1YzHAj6VPZMbepP
8Zn57ZdINJfm1pAZKEVg8UR2bo1XBYclO0bOR/1MqMNBvPEJqE4AtOGod2/JurZdI9R15k0V/ioL
qFMQCkP8YHrbs7RdHCHPy2uLjLFK1U+NyBIrxMqrLPRGW5qEQP7P/iNbFtRAixo74znYyDPigTp1
D0cr1zJp/OIWUmDRKpSvYRHliKCd0+I0s9lZBxDTEL54plZg0bgXvGXU3FTRzyWrnIY9kVkXHlqa
PnhoOIgm7WrR0Pilhgz0nPCFu/rJ8qU3tPu6/oUGOrZN6ZXBcLUZKmwAOKLd4XC1m6h0Iab2zCO/
RDthodLlBRP8XxQhFt+WzQ1i45J8xgnsejwzQ7+5I0RZcQrHKE/fpdjiNpEoAEmZgoVjV2FZleiK
0PorMOv0sEWhb273pKPLfu4in0NwMzrJRBzlM/DyIemILe2E/f+hiPY/QecqP97c5+X3yuoPYPS7
BGIPMzNH66Y2QP0TfOmEh87nnu3tzwVQeWvsX2rbsXKhSAZ6mAgk1SouPwQ5zGGxr9a/aGBmjsBS
vDU1NwFzdfcHlUb6JwEbTjMU8FBRmGy17TwBsGb/0+Eeg2PlnsPmoaCDoK8r8jwQtoCSav/AkDEI
b0sABd89M600qfs2IDo7rgY6bAaWHfYYt1qv705hCmkB/EFJW3LCOyL6U6RMN+Viqh0/qdQ0s/Hb
k3ClQ5J2n3YxNJvCGi00akvGj9iTft9xs0O8GcSfoECnEvvORbjjI6uc/gtfTV0AIKp4gi/tLfGq
0KBu1Oyv4yZ4/kpCuNqpVAmJlihMOZWLDBZsH6StAz58b9Nd+DfKojqyPLr+giHCDcUfBP/8iVyM
91hkkU1fGqfghZiV3PRSSA8Qg0BnuRLDMhS58GLP5iOMlC4c56TcfxHBIJ+hFP4k2BKzr1WrCRv8
CWgIkYDDoRLmJIOptPX71b5ZwW8zMPyfnTNGtwefWx/p5pEmBaNWQDcRY2njHqOm97rVzPb4MWn3
ezwRKq/UqDChGj4sLt/1nR+aMZuLdjZb66QO2u7xPgClA1BrJzMU3YdcVOhfkRzXsp1wyK17g8DD
xOuxYW8OBakEaWsL++NYd1MOUxZhx7jC9mFooLfUPGkrMezD6K3rfZoz0ROC3VUP59jkcKOkt6yU
YBLvb81VFWRdKWwJODy4kbKvJtPhsZvZIx+Ndr6PKaC4v6HwWnXIq/Ji7KVhy3sRrYOHU+7JGdkZ
1ES88qECV5MqZL8dPokUW45h6VloHEbnEnAnpdqCI12ND23XUQAwNsB3TGL+ay8Ij23/OAOoAZ4O
Ku+7uCcGHoP8oxorD8urZ/pLbrdxh+QWi31E17mmAhv99EPpf7oDA/RggkW/QRSn4ixpBti9mwyC
9g7ygDmBgSC/HkAaA0GsqOEu1OoIgP0e5l7EIecZO2gjoG5sRaZrnehOnirmlH9XMhnyjghpOZX7
dsyEQXmJuJjFVboajjGIgikwGi2JwPawlnJpHWUjTELO/HC7YtkCUOlp84c+tHGccH5fRAEt0joD
moprLw3RuAgxLqb9/dWVJ7BYvk3rIvZBtd36Wes+n4JzOiuZYYO8mSfH3oChrBuj+IBUfIUyCphI
xHkk6I/xlfdw8ff5OzAtVl3z13xq8LXOqW/l3lEL/r3yeJqrJiHsyjl0H0wHA0FklPS3mNXlSwbc
zU6149j4q/mCPTkZZLt22AeKlLXPm4hG1Adzp+sXmgDZ316q/RQ04WX9XUYHaSv/EUPhd7UDAA2E
JxMH6C67xS/7UNfkf4c23JIzCvxoPYQtHFEyBILaRYJvn0sZDeJN5yIsOXxx8xuOaMBQGIOcZimN
s7AOxkYrWGzSKJmyGNhznXUPhKNyOn8vq26s8lvhlJernCj0Bi1Bq15gQSO8edmSEPTm5QyIRD4h
mD9T3QKMXdrIf8GXSivX+c1vzDZ+CKn7HVV0MEDBPbwnYwG2h/BeGQ1J/jCz9qA+CdUjx7PUVmkP
q7sd3zlwuppjUaTzZZD8cSsxRiH0+4L86bupi1/jgsrMnZLTPpg93dsIeDIo0CzpTiPFvm8I82zS
xXDJrpLjbfyWkHz5Ykwi9+WRukxJc2lnzMLQhFPFl1RGCjzhzF36lg1uAbqK0IN/ZDzLV+Qfoc53
MYenX6OA3N5jE64/13OH66TChz1y7R9yRgKSKnvuBci6W6bKNk83Zwf1G6fg3dR3ETsSn/50o//i
sS24CZ+aghWwIcDNGiESkILdUZD++WojPc3We+Ld81dtJ5QLvR6Eur9RpAJ45ZrdEbpSogZF0VSF
B6EeckpGMr3UiytwpN7IqzDtGRtt/0CkrKLndcl9HTxAom18Kq1HKSi6bmitZhLWC6Bqhpb68LAG
a/uiT9zjPiv4okqoxZJcN82G4LvscivhrswRsMAvdWYTSB/3spozxrs8yKnr6FchULWdi7t5KEIW
hyuhuwXXEEfarb2l+dg4ulT+3LELFLCA5UL0+zcFeGsLehkMMVv9mBbdQg6Sgp+tyxoMRZNDrFcf
Cc3xjRzTbETjTd2dWfQ/52db2cQ6qTm9r5XtCxI9oQ3T3DAhu3gLbr0ruTFBCKGIAH6EaUYNWhgh
DFZMy126eIYL0rPpBe7tYY3fXEvGnvAg7zeFGNywEm68an8KHY1tkwXp4WU2MqJFku7rMlqi/A0D
nNRx2tuElDSn+DdhlkVT9NYhyyoHM12nTG/hOZrvsZvIsOD+60lL9qFWuUJkCxWNXR3si4ayTr5w
/bhNVJNk82mIAn5IFfrsPvshFZS0iIKmTmzQA5LcWBzNOTBeZHsnYH74bMTvMJonOpgxq6NXbrXj
xh3IjZg/O0Tj+iY0cfvGYAf2N7JgU6e6xIbLmh/pb492pzc3xNuBa+M+Ze/054uyP7tNVDAaWJKh
4vqqJ0Yi/sbfi9NcBjhKI/FzDpk7MM4xas+ZxPV2gzoqM/13cZGs6A/pIKy1WrFdo1b1G4ZblNA9
vhp8vuHfTddsu6l3fX0EodNRwAd7EiEzmMlavI7Ivo22R2H/b8jcBsanPgu0DSL9oboHLPOZo/13
wRMCNYE7QcF4NkzC4Z+npVFXf2PLXSpBKASQ16766qJJzYMUItFCu3UzqMNNBLyk8d3puPFQXP9f
doIGPjUSYCJLPIAzMmmgcmyWnYRYmzOaw9T2ckojNuV4H+cw9abC7L+0d8JOUAelVw+ETZ5k3z/0
N/h5Yl8FuRiJ5uQ7I7/KR2tlS8ycBu9nF/Kthoukz6pA8LYi6uqnsuHnEc+R3MDVxcjhyTiHT5Zp
tQKmPfs/XNiLKTxMv8yRAedgeWvUrI7cpdkvxO4IoJNB45hRaCxfl6v8Y4Trm3SR6FwEkzbNxhRe
aThITtTsjdq9+zvSFKPzMrAKYHImNsFMXbdRKED3VGaGTMMFTMEWbcoUscds/FVoXw36yLCGVQFl
+k7h6q8RmmHh/Qlmjhfan3ElWYTDQHS0aPCN0SoAo7VwphD01aMaEXKIFPJ1FKLZmADKt/zOkta4
mO1/daT6fwjrb1CWkozmQYVWQyD4jmMmRtqfdKur0iD4WZ6JLzprlHWL4Omyoutxs8rr0/zOWRxk
MZXTxvJc9HlPbGdrGOMXRx0zWAE8txfY6znzFVz/cUilf4YzOEbp9KH0rncFCXuvIiddOBsnDDBm
2iNsztDKxZPPEU8Q0PD7hQqJt463xiC0+DqKqndtEUllI5wCTNX276EWAhT3tszvCH1frvSlNiTb
tNuqrG4Y2GXMYXjaRHFEnc2+GRKHZdnoPyiN5uGwj/Gs5vpAceekTHPgPrHHYdg7M3FxQLgztTOZ
NvAQrRZnMVpO3Z6Fk7PcacEoCSOLwuRCm3rfbp1WQ3JeS2iYjbVFLvGy8BAVZWDeUT4FpHOH+aqx
zbcfRoDZSsZkSsrZNkpjeR/lPUk4Pep/RfEh7AjbdlU7b8N1xB/1qQpcY7uJluNC5aHJLtV0AaDu
mg12leBlTFjTmS6P7A5d9/pAWB+9g7bN1/mBZIAE8pDu6HA5DGL9p80IM3AOAJuGKRvJQIBmNVox
xXPAtAeqM8bFNJEr7bEoAgaonFBwBUSGeZyUfwtNHSRc2xmQzelgQEfNq4S3xFUukbEhZuD6DPN3
RnLopH+cU+0sc2xmQUzAjarVsWB2qTIvuBG8zJWcU/xEyg/8EboLOa4ZVTcfEGKFaoqI6kn26v0q
fq9zWgemrKBBa3cMPs8k42LSsDjIgTs/q482AKxW/PQFeoXvHk+93NiyM8k7a4XHkDefoywHG+EK
7SBOvOTyqnxARjd1f5LTnkN76wvvkLrZpELnLY+LcbszGUYVZoeCdIU2eOsJBTnvfHuXPpoMa9pB
UYijiL3eoN1ik7AHO6nEeM4fvoa1Ylm267JVWh8S3qVHJfSMKLCXtlYxX5jjqOoxV1MmT/huZeoO
jOmiCbJT/S/l5gGumJIyD2QYAIPsRGkjynrZ62vVvsqLjFV1ShBArxsJVm6HglJ1+kudUrN0aPqV
dfVPUjnzZABhT2vO+HpemFPC7Y48oGdw8MrDH/sjsb0yUDTm1V7FXzQmi69cPPuLIT4Dd3CoKaZz
UZ5sioT5tXeKpbeYOVEWrePAOQoWXRFiyjFw28nSzLzfIOnO1BsZKblp7lTrMiezwnkC5LEVRbfv
/y1M/0eW0vVyxMkfM1RJsnCjbfDEUG6xKi0f+NmdJ6/rfMP0eYDDoHYR8d9zspPiijUPHGPvpZO4
65UwBv5CQwgt55i968Ug1Zf/vf6gGgQdhRSK9YMtTRulRV/AsrQJHZ6Lo89WE3KABU/Abc0wQQ7w
WxHen+vb9KDYv1Uz0/dla/kuieg4Fke2MpQ+gc2q8cwFFD4Sd+l0Ho4FtX8t0f8p4WM3cLUdUwuB
NvcLY/m3Ozy5LQFgCTab5g5n+l7I63MrEV3lN8dGZBeYVufQlKelq7h9fPVbK8hrQw+Vydehf3Er
aCtM/R2f9k9l34f9d/Mqp9MCZKxNfO1iLt4BjUOejkk8MxXD0Yo8hJs+jwg0VGRuj4+D2UUrJ9UE
kNvY48sdQJrYLF9KmcRe+B7HAcX9TRo2xc/oRAy29rwPXdtcEi6k7GclK3Fmb1r/e/eVbPVEyKkb
aJXeDLp2IDOgppNVxi5Ei3mpzSQg7B6ESeUsvA3IBYkK2JI31X+pJmZrW2IVjywlBSDa1JnrRqJf
66EHpNCiSVqIs573E1/0/hq63lY8q/9dKcrdzf3P4N4v2o0Qq/AmCrdknZ3KhDAfNSEhLGfVC3lx
rAmEdYN2/fk1lo5wOZEABM/gr8zgVg9sy1PxX1FXOB8FdUBCjOnUmzA9TeAb3jKjb2tiUtz3GMOU
EyPphPqT0jyWXoEMVM/Tdv+utcAPzVlk+nNX7kmcBVVlkDxiIP2Xo9fslPCEX9H9bVebyZT0zMIp
ZdVaMB/xrE0sOrxjww5QUp0cc1FZja2TklZmuUOcKTCV6PBVsJ8OqKxdWH3IhxL8aqHjQmKJ3j2r
3KfjnWyc95yGGoCUr4qLNlEKMjG+3GuBrI007RG1ml1/o6pMhkfrFZC2HrMXB+xWcHKmwNDQtT1T
3AwsbjYEjKahFfwi9hBCn6CnU2TbGiS0pYxCXTSLUymPMfnL6E96MkyVjHFDJ9vmEh7jG5LzeoG3
nCTc1HwYyVjXU0GTY8v+M2G4GqpNH09F419kfRy92B9LsPWjoGk2Kp8eapT/QW9MXqarqXhBv44G
xUWp/wlgAZ7VOfC/FibzlxWNuhTz4EeprI7WfTaA2LgiwNU2PpY++Yzzg9Dp0JfK4wvjJCsSMWFd
B8YkhEibiYaE9EPkTMNTHuBiblE8JFHapitwsegfXXA9rMx78NUfRld7iFdMvCh4J5LSiqY2/nd1
xfytbxqZ+bj2GVKQ5H9t2h1mpXkRkoH3j4r9U15cYegqq9MFtCXe7jqvYuJfC4x8Is+SVDgQLU3u
ugwIrSSHHNg0Q02C33Mf4h5OSf/zjGAkfLXu7iDshh+lQB4Te8YR9zSJrnx8rwvnrsYGjzqCVid6
+gZgkUuGpS/lSno/NqK8F6IK/dCJTf9pYCArZV3UQAxOEiev1sXKh4EuO3g9LVUEOzfBLJun8Qjm
y08P57ByJsueH+pFAXGyxRk82REuiqkCQeNM3xWhWPat+TJ6N/Zn0AebGP4kzXeH94iA3FiUyh4k
1SP3le1eIlodoSHvQ0NPw8KGkqk0iFQSxZH6nsD9COMY85oI+7SFIjA707NoXEgxzDS6W4vZJr2L
DNM7Gsokffk/nZc3WHW6Z2TxxXqL1g6mChbTTH8e5b9t2PkXtqflwmS6//SVjGmuFuYftUtKW9cI
UahoJ+Xhy+T03ktZGck1LxSVQMrNl9Lbqt5nNJOWO7FMG3m+iNhwFmm2KExhlCEUqN/eG1DZTsxv
rE5feg9B5TlAACFayswmI3syG3vs64ZpEqeLbCXn2NFmlpPjshg6Do43bxTbM5m7RfvA+Ap88EUA
2UbznqlFvL0fcmfiCwkRM45nyQeZgeEMZmnYtjsKZpwWd8+QePV95QCSqyhMYW2peMyTTECzCzqn
U4Vi9R1uaSF4BAdJbA7InQFZ2wn/ypiaISdx/U9YhM3nGZC9AlTqkj0niP4l1fsp16xBzDcWR/YL
0d+R7h0NhqvL55E4AkcRj13Ml9SsT9x46AzsVfwnU1RnxQCsDBME30j2q/EXVgJ7LU0YYd0AM7E+
CRLIwpGaTJYz0Bn/vqVuYYvSD9DXm62c5ze3+e1yziGq1mcztP96TPKeBdAoHj98/Y1v/vhspemT
Relw2xIJmVxi7+0ZBqeIt9t0M20frNcnkqugdHPnwYFQ3dMrKtfsIvQtSeDzxDLAnzdKEH6nZi/X
ET8uD5IfE9+Q0u2Fxfgx3K5Wiz/CKgA4qaOfzTi8DgzsAXayrTNUizFdsOjPIE/WKJ74ED56ZgPr
3I+83A76uBDt+Kff+ZlMggP32hCFFAh3tbXi8cSGOk7NnAzmYCQMkpwDSrTQ1o30uZqZtebw5mTJ
i84XJ945RZ8l/DRH+OcBpGJZbQe5maZYfcSeY+SoMEAxxcF+2q4WK+1jOS0G4+d/i+Cid848FVld
aKRvJLJbrcfEEOngcvVdujhcN6wiOzvYpLkh4r4iSOXR1HyPR59aYJ/448zIXyUg3mogIoCCMnhk
Fjw+FJhwaGTXARDHuGPAD9psjMb0iIc0iarLmp/NJuCVpFEZg3VVpe4D0HqpxdsUjrjYngm65irv
+bAbyV/gJOqO1lI701vMOShSLkIZIOtXe8QxFt6TTJrvjOlhebE+l4HtqpO4mA5TWt/WseMGr/Fx
kSUabYGNoE4i94dIpjx6jGxB1+PrcOT/qpyS09ZNNuOIGuYK6aN6HM+rSx+VPaXbDU9dw5zFyCgO
RoBgOmJStCVfyNrDxRV+NtVuhGObemNtoJ+uGftGa2LVNa/dTNLr+k4RicT58ZzuDRErcyHBXtRy
Pw9G+yq0zJSuakqmTie4CBUX5JAXmBC3IjH+CQ9owcLWdI9wkZHyErv2u4CzZByP7KOnU7yLYFvj
yVAqgU2p5dlIxdskTPU7JG6UxTrD/sv0Pz0zqi9pRCsOwt2sgxv22bT8/mdvJTizel1m7+rPcXaX
OqaVmwxns2RexRhGaVleQvTZBsnzuR49uTcwn4Z3Gt0hD9ib/mpCAW7XWPFQPsJhYIrubk3lQDrM
HDEPzlH/EoFXH67c0EvujvsYP6UrSHN0qSqhfSmwVQDLNYU8oE5HHISqmNLU4gEzFSU19GU2JwNq
nBnjxBQ+aNX8awMVfCtSEojHhqOTDmuBDxAxaRwiuB+8WxyjuCG7IG0FOlS+RJ9lTbQl//XdlIOs
Q9ESqFb6h96cdK56uWznAhKdszRpg0aFEMQU+EPYTABw9+v4o5CtneEuJxHKTyj/7UFrnK45qWAa
Phr7TgHIfWcoQDaCIVwI5Xod+xpSioBzhDGQpp3Rdi1LtJwedusNvBBpFtZWx5BIUqQ3E1tnaWpj
aUnNSEEvzS5TrLCSUlYXPoQvcEY8rzpz6OJBdBIh+C1nvd2s1G4OlXFWIVCDHIz1ol2zcRK7QUbf
yNoLdy63cQW7buWQdX3tPyK3PiFvDwK6tFG5ZPaKodDagfP+m+7VUrVrAf3aLx2PfwteqPYP4/Ja
TtpPXSyAnh5Xk7Lnge67stXWYYEjqbEnNKAvYPiwfkLtTkIRifIdWKmQPL8uq7eaWdlks1drCXCv
+GNXmb5Lv5hlYFyjDUm9vBf6cbCwANggPpS/GsAVmVQ2Lvo7NA6LAlc0NONDNjpO2y23qaso59xl
lDgZb+gjGEUj9f4o+CTpgOqbWsfZkAQIWYKQN0RjCvn3SYZ4NUYgBj73W//VL3NCXQgYmNMHGurl
GX7/zUYXQdQamVnpuGVKX3Z9d37C4WwaleReSB1jz7R0oQjB7cmjtA+Af/quQ9hJeex5sBbFtV0E
kMhP5dUSkYbgW0KUnmzlSq/VXLCcJcmKHV4ha1FuT+LzBXU8n41daIczxTTxioj5jGfK5H9yxYD+
ocHvgx1QtmmNEosmY7YCq3CoL4RekXeg2QAXcAg9YmLGXXGjBiM/Ml7Ta9avG86tB84p70KTO9rr
cfGJRFo2HlxSQ0PEoyzQM3oiwAqv2yV2bg5WUwvOFxJ60uFele7rBgXEEybvgFCqwmKcmnvlL8eL
t5qnU3n9FnVcm3SoAXU8bg1oWb1cKWrHFvrS6QCU1kJjXKVG1Wkyw+M7UgWAuu1nT/toJ49IjsY0
2MV91Wz3gNX1ExBGdZJetSdv2W2vfjMkmKFB/EcXVitVbsY/BPwXao/M9tGEJs0nmH3OS0H/4sjH
eYHGHo+a1HucWkdL6WJ7nB+ZGSu2Z48XtrkljT2WcuutlO6kWxJmevskz3LTDtrGtcHd+7mNyQoh
8Jz8rMIMgAEh5ZNo5Vvh1BuY9RIeiEXNb9ENKuQn06bopGXd+sMLuHonxMMmWUUGo2n/ldzxh0bl
ex/vZxjCtpQOONbkcXcqZt4VJcrL+cMHQ3GdzMKQ1l2OW4n8a6IC0BOkg36eyTeSgpueZuxSFnD2
131o8H++Oq/EWLyAGFX2EZtRW3zos0W++9UR010SH5BaeJIND0Q320BdIm53NZwW2NJz+xaJtg3F
TQgvyPeC7ZQp/XEfQjQ3n3RxItU0e31pcRz0HAZy6DLFDqvVHRhBtx/JFQd9rrzSJlmH+2/8l1CD
OIPHdNuFw0Q2LDAr1mmbcITsiupz9ZY+bZypOpKniSkkg7IrZNbbYfzuxynMuSplJK0wy5WsXHP6
XB3CvjHf6dTNnVf+70yFkyKtHUZrVLxIGPu9pjaKFVM8nWwGqbgNYpjJqnRw1gqmwlphvkVVeO/W
AG0561wrLqNQCiRiI7G/FhF9riB4T/MM/EEpbR7Pps5nj+Pz0PuRWUZjN0zCv8ACPR6ab08XTI0N
j097w5luks0tY6vOrtp6cVlYG38/wbKWB0ptdTkzwTdXU1Sle2+dtiXKs1un+MTK50AXKz+jhueE
WZIE2BHtKnT4hDWHZOLC8u6GANQJ2lhM7s0UUFLItEfii+jQi7YATfawaSazt1F0x2KfD3jBZzk2
7cdPiWz3C8FoUmaISjSqT4QYPFg60cbriXBjPimnfaHx5eIZYXoeSHWB+uUlxLl5xAVBuFrnvGgN
Gm2bpqL+RjWNAC18lmmHBdObosiFNPMBLpEv8uE9g/XhLw24gF90Rlw4tMFPETVNKGk9HrAcFnc6
b+s7AZ116f8GSsYlp3jHvmi6eq+xiS/6qECCaZqVMNIf8lOqrq1qve0RoB/Ug8nT4K/mOAOeohom
sGoFFqOeDxbDpNHfEeGyBQrHsPLqHeuN5NFw1fuCyjhuV7V706n3hT4zBbu+Q2zK44SSFGnqkH56
Bcck/LwQfDZfP6512kk2gBTyWV7LmjVCFFbop7KgHmNGHIsTj8QQbtJIdi3w+9SbIqgLfbPWg+M5
LZqUSMamE4MSR4ylG319A3wDQQrWmfw4BkxbEP5GlujICpXfTRq2KQnTlktCoaGGL7krbMcB/xjB
rp0777GH6QvxMeDhfaDJ9MQLQ3dddHScJJVjfThK7AblHHCRwDN0KcOix7LSkwYxdbqaxAv+5mNZ
JC17ps/60RcQVAryo9Ll+2CogzWpbp48wF/8qKn/itVhn7a4ipR6EQsSahKOSNtDHBhKaUg8vWwP
YblEnvAg/V0X+sFVSuEDrW5hzeZdxupqI4CuCEyK52y3gXRtDfnP1CztOwwgfQ5TfNYfZ4HapXlF
Qx+/Xm6S2ObxpgmauHpG+z9Sqayv6vrIAZlKkDcx9JswzSB+CjUgftp91mx9hAc27ERsEJaJdzgy
4QUPVC2EdQTeTPXgDeP/6eEY3vfg/F8CARLQKVBGHsqU3x8Bc9Oz7Vk+xR1x6N5yIxWQBUjrXwWk
41uVWYHgU2spfs+vOl1Hex+Qt1qUBsVA3SAywAS6XJ82oHyg+EN850C5hRrCGdzcAfd40eP2sT/0
sPyK1mABE5n+GYWea7+S37720t5EmD/L0mX1WDGyai8URTUpoehcbgH6GxsA+UfSp5zPCohghBcL
rlyFjdKXp3OzAMdo1SOAsOAAiz/i4vM4NOY5qwEe8F+1lsSr7p6iH8dDRrrEILGxJVrRaUBgXKR5
ABjlAYUC3aCuIkIklgoHo1LRngjZxix4RcEv0o2wsW10OkuyheDnor7iTaBxKTJq1IBliC+2WkCp
UKZxhUq5ljblg9wdqScWV61rLgB3Z8zvUsoRNjAki7rdwtZb9JfiMLhJJA4RTrRdhgJ8eHCkDeuf
ZRWUP/qMpAr3ner6pd4OTUeAnnWEYFowi9kyDRfY3L3C9HoQjl+/UiEvj95exDa4EFNDuqM9lgT/
Yd5tC7FIAUwXNmaEKeKmBurmNXtrZ5sSPeWK5F33CSEZ1dhuEizV6Y5FgS/33gjMGnSkHsD4OmK2
Sy8veDtWfahpK09eTvr6T/5xyKd4nt4ZnOe6zDEQnFIICcn/yt0z6tixUfVtsxqzst0Hj/FppN00
GP/Au+zW9XHChmi5Jp23ZhLoq7Ke+K7my4CwssJ6Y3QM7uVcTLi6bkyX45/k+3MzLuDzrgBrtGPh
lmsI1rpcNuX8YCqlFL0FYc+i4Wxo4pueMdSt9uccfGey2HZV8g8tzwzbXx4BuzMnct0g5HIaIf2A
cLbWicg96HutvMCszUn+4VVJiWizbIAMq1a3c0fTmoQzOOCzN/+3QeOCF9G4Ng3jibfN2hvzCzSg
zXszPE8w2dnEHp4S7GgvUL3oLtj3IiJ8Y203lHsU2KF18shK6SfSCt7BF0m47tmyj05UeRoPXjJC
M7Zs4HX/cc1/4pt6e7mZ1olXoGm3NClexI3xV03EZlA29JEQNolMAyGBc9qxQtc9roAazWswupvm
7RXO2BVDNvPIo41MKRvRE1BML7/sZD6eQQpKs7sWr0iaTffVNflgGJvXB8+Y+gFbfQZNsP+z4sjI
TNRl29GNUzbT+vymcuqpKRnMw3WcIJfRh4jDUiuHNHaNiZVlVUUvgAF9DSygMcJLIx9CfYoKDPRt
ZBht/XoRnJ42Ck5oHBtJVyYWkKK5S6a4SCL6gLhEaGiSfTDwt6bDYZTI8z8YnLi9MG0jatcsajVK
DjaRVwk6XMaHkLpGKJVmjbEirDG7vI6VUe5eBbF0VMU9KjGL6Ug7vMO/117tPlY/fAm//tH/x2nx
0CRPL0sy9wk+hq5eF49RLczGOPk6OzHZavFqiLiC6Iw8zJkPWMFSuxWYDMq9ZxrvZv+/CyU3s4V9
8e/jqkUjv8TmjQkO9A9SU774OX5md3BgQk3whmR7nEt7nWOrdX97jbXIQEVV7UsYeDAbPWRADFst
WccEmXCw9SrKGGre2zsR1nmyCPqfaaCGqGt24FCeKKbUxQ48Y6qG1meRJLDZaI9azlN2NPBt70wB
phVF1O74FUipvkqu1XWEgE7cV4aThKgIqumJugKAk8PnY3mgG336VtoeBL95YsBCviJaj3rK5RLz
c5zOgYNiXotE286c3qmaHnAKGUKf7IFc/fHQdcP53IpvVQpPSnSjlPN6lo6y/8EBYPRgYDXn3wIe
YM4QannMTrtaGRKpvArqLJ1enfXVhVZDCQNjbNmm46i+6gMZX4v2nZV2PnptYePhJwzLDATufWzJ
l7yfoLvR+uGIM0wioO6sx+Ojj5BIODVM9Ofe1eFPNCa9ugKAby2OCg86DQhMe5DCsSopA8CH1pbv
KCRwcoGTJ+HleDwFMgb1jdekk2D0O3WUCEg6PDHRDDQ/I6kihoxU6xzpmPWFJCkmmOEXArKQplOt
XuCGnFRNlYbp71x6tH7QXjWHw0mEHihB0Kxl0gjioVq7aLszE4i8T/rkvivJrRnK/L0dlAgXDlAZ
GXs+LRpH8iuwab8jJpN+NxzA072qSlAhKI1CcN8sFu4B33BkactY3Ub+hoeS2fQvae8LgUiAm1SO
JVAMJbcprSHqZ3ywZciOAiQMm6m3Q2zPVulcjjRyykIeu4tWn9r0DBcvLqnHulZts/8Jl26SOQz0
WJzRyv9pL6dJGGldfq7zGOBM3IEsx5OUki5msuxX8/FB1aazhZDcIIsbP/JWSD+PYth77qp0lJza
ibnLBpfdjktd9YLE7edERhOoG8KH/au5Y7MHbBw9I0c2vpM0aZh/h0+B02mm1Hvt94Zhw1ClihRu
zJxH9dpOzV0uYL+t0AKqMzf51qRrdxLkOXZNvPFCa3mYmj3+bh9ViGCqnmTC2A+ctArb5pYjWPnL
sJ+ktTpchReUMl0ad4/ZkhXoejrEv8QKkkdApI0OQs/ofZOOzgpwA6n/BAWhHoxSZXD+PytbwmE5
hcEEjRy+nq0GEleJYs9mxQhkuBcUXfBei1w07VvFpLeFvhya4WKEup25hKcAaP7H5M4hqxALrWFk
roTUb27cpU6Fpm5AajDFLF2fIheuOhSbhY1kQFbmB7ZyOClOcBifbU+tIvIw0DG9LhOp1Ua7gkQM
CXuxj0/KTjjeiRj8JcrUm/7pZzr/Vsq/I2VRvaqgmNgTqwJmqImf+5V51/UW7OEfJHoIJ0lAI2j+
ZpCnCsZbQoI0gqOauVqKfeqqm2Ha0AVrHemmXlffq04iFNokYq946lYwwybWjhRwiU7FVCAz6Rc3
mTNtbPhj9oT9iss94DUJ5SGUrGpsz9eIX/5rEBbnQ9TKT9eHS3xn36QjIUGLcEVyle9TbSWwwr37
00RV2LsYln2i4DxhNgYt/ZESVk1a66lezV31npqyd1+KJerePCaJe1r78PVSOjs7evkiedcxr35X
B7+Qvc2putpd/A3gyVXc9CLCAM34QIyGzEorMygqAsqv23xuNY5ygLiKKzdEbT8swWZoznixPf+t
zyRKBOaaHPTe9Z5zP+xOgGqxCSvOW9V2XzK0b4Byz77UNfWzfryRLzSDeZLZxCT0Wg9zW9BKWIVG
l8dEFO+/1IfWx2xfiuLTCEQnsBEEmEKiaMirt4hyk9seIIW2ZlpkOE11QR11gDesrzI3yLHLs9EL
NpUKhOVxH58ctUm5WG1uWAMex5hsT+UsPvt+26PrxHiSuzl4SPe+Cka3x6lSRO+AnE72WNK5bElE
LhU1W2FpajE2F8MBYhIXTvaqOxCNb/H9vui0hQbUfsOMu5kwILhJy2U38biBQ4dsRd0r0n6pfhO5
Bo7mr/3KeYOVh4xRMUhKvQ4/B7/uhx04QQqAdd1RQCjxUDTrX++k45U+4BcxE6mJMWebkRSeh5D5
ISSnJ51jCwrDMrzvWxXGu6HGgnEaT0KBj+g9CgB4K7Fk1z3g3j6lRu7hrFv+8co0TKloEI8J1ipm
flEboSNSowJghRu83NMC1NZK+qvY2mh/t85uSQE/WiACCRH+dECj6VikMrCPC6aKXK4Br4+zK8QO
NykAg2O+m72GeHMKhDZnPqLGp++7kIdwLquIIc8L29gWdDv3ntcTYkxk+NjKcTQ2LmXigtyCVQYg
LubOoOKtTaapMyinJVV2vBcX/F6qSCJ71IbXYKYoNuIkBdtzrDkuV8Xq9P5na8uTOGL2rJ6m7M7R
huHcBcz3YEHEQAsEQKh5nh4v24p4g6rykuLgXCQCNr6QYKt63PqIlDQeXXaiMc/kHzupiqHCyxmq
aOBzayfnFurbnuB9+Ta6p/ffe5+YRfhQsPM15IWFiNmTgmjDx4uG64DTZhod2J7dF18RWGgixUxB
OCmeyrgV8mVfGHL+vAARnFKTnbk+70Kk4KbkVjMLGGuDJ17BMNFoSjLNMTUcHDzYirS7XzN+weLB
lnqR5rndgXcrjWWPUFjc7K14BdYE4ZA3kwAnRVeP3qpepW5B0WRb3EfFdWQAnkDNMcGZbOclxGgJ
Kx4Wn81bDVSHDciu6dkKrcoJbnfZ5dXVO97DyIz2/vrzoOgW5FLpQ81CN/6KJaQbGCqRoCDDUPyK
P4SR15mb4ZDFSs7e9YAg0+yowyhO5lSuN8cAte1UOcZjyx+E8JGgydI1BFd7mQAu0d4VAlsNoZPo
P2idoiy2DM95OzEkfLpm+e3ztIT+E3vUULZLsbZDqLXvn9RaU4YO5d2Tgx2VvCGeNN5LpaqqgcoT
VMVF2zAdySm8rSzeugv7KK8PazbrAQ3HmUFVESL6IYCyf0hz4WPUjiI87onBxl9htaqJ+IoUgzwn
iZLhvri/sDjA27hF9CO+eJ7e+4xZX2rkAGM0XRPKbJsLWeRSBa4/WGY8V9w7FbZVfas/NetNm3hg
8V6MkIxoh8y4sGo9lO0jSdr5gj4xkf09Gi0spLl0g97vPbwF8Sy3ockWKhKxqkhqFJcHQWAYIQRg
UQQwT9KX0sC6qh3MpthehV62jfoFCHU7xmSCZg6z4Lx3pF5vX5eakfOpCHQu4+hx1cXIGehNFuPB
PjSDlM640I14zU9oly6vjEPadPI32irAuTUj6Tn/I53ej/OEOSSKZxXkh5vBKTH5+g/yZyIMcKTD
K6JHxN6IqPuBT/pvxRL5e9M6HLdcCRMpl8eKro6p4OQvljSupke8OQJl+PHKl0UfUKLHLKQ/Dnx9
u4kvLujvNFDHP0ya5+hT8tNUsTtZR75yGjJEgloRl/jtXqiolt/yNRNDFJEaPioGfcaPeJygFSvq
VZMocCXpliG229yGfjWyqNpKbk9IjV4Mom2aINV8H6E/qHgkLT+5DqMYtgstgtLAdUxQ4IRsK6aU
R1zgi0ukXzl4drs6bpEVvdorWGOpPnZS59SeMywBZ38u3dkjCzhtf1ExKd39MN77srAnhpHqQ/r0
6Gj1p0Ego8pp0tIU+pb3t2WMv+F94JG0xzMvS6i/A86ElUwDanFuww5+Id6yMFY0WHZUNFo9nXnj
D1htJ5iX4qK5nknHWNvm8pU6YkK4oH0Vv7HlS9RTCbzPZqgOHrZL1flpnvbnPrcGxpO823QlqvHy
PM6UoiFPxpAxVxTc3B3RKpPvfFdP3EWF1llfh8tshYDLs5+r73VoiiVvvRq+Y2eNKbf3do/SujEk
ZZGLFXXACrT/y0aYElh3aTT21xGigtyrq3BKCTy8eCb76/m1S0vlCdVxmNnJHtIhr8j4WGZvVCDs
bBaCsaiPYnN7XZ9BmvrlRnPGao5NoiuNb1rl4z7alb8dZi0sy5hIWLkjN9/yGvzG0m2uH0pYL2jg
P/evubeCaI8I7tmpgZJ8psgdP20yH8cHfFsIcgQjoXxy6UBCl+yjpNyN3pAO+Or12tmTsa9SN0iI
Kas1VOMVh1oETbJ/NLV2x1qAwEkVqRpF3ArJriqBIV/q5ToOYzFARsXdVDZBqGqvZLsUXuBy9cMt
xau6ihk06mAA73RPA9o4IpAbAUr0Lfv1KCS/PQW8aOBHuFBvWfEzNmjR3uOAkA0Fdb17xCI0O13H
yIf4F3w56gAcXH3u0gsVD6dRbeHiYdqylK4ySgxlkKJPFHBc+l+hGomcsb1jWouSnQDb1TlfJy6p
FFsVxa49aVUovLrWQuUUx+4G+jDuDqPm7VgwddYxocM7ylUzPsGkyZkDC9XLn4oiPT417xwd6MMP
Z/NEeAum1DldoQ4TItvNggVG2iJw+IO5il6FPi2OunfezMLbpAsKMK8rgrKPFTSzvjnTUW11EJLa
31NPuAL53CQkiZMrnfjQblzZsqG62erohbBWgLWC7Hu4Uea3AYsxEvb9NLTtWGrABBiLJvEfSDXl
hG4BcNdKdCxKGpnWUd157Wanzgh8gqJIhrqLYHTQ1k3nFo9WT7aqNkrBacNx24VlAF+RZ7l8WGNj
TOlQz2JVHnHVDnrpxGfUN59eT6rn8Twt5nnitxrrOxhnY9YTTywLHYInbGVykjKV6CdlXVCjux0+
HV0EU30RtcF2KVHkPHruJJwoEz/WieuuRjwG4gXkFLyLJQOMF5DCOIQHOD3ArzBvhCqXN3chCLx1
HeFepNU96YvTL+/+lEac8QgMoLLw0ZTXG0d0mxcvOPTYZtGfVGflc8cnxESkEvDy/gGYN1bgXVIf
TNhKA8vxTFRJeaUPRDatdVg9rtLzrvYAVdRUuNxu7DZNyuwo5uh6iyF67exfrMcHV2JIhy9he+e5
rN0WNriKUcxLWLsLIJTYx4Y3T2Ynw/9ukRziMRErGG7RJ5FWPkwnXVLd8d5MpJHQK2yL/maG7z4Z
Qy7kiiZ8mJKjzRH2YNnFqPWKlfwWfuJ3bkyZBKyj2aYD/KO05jPLSBKVG/8D8M0oKGnm5C2aYkO4
G1CIHxuRd0WgWoD5xP5Vn9uQu15FbYimEQg1OIsbUsbzezMGkJmvB3y3FehkipGhTKSGdL12CdyZ
ftbLZWXIVuhjEOYTtNwFt4Uk9hGoC7aNxPH1UzWi0hr9NpNQf8gOEF+lPq2ArL/Pnt/5ZoKfVJaJ
1XIEYccFL6HC4gYubPhTvCDopRPvUzApi5QYCM9JQfVGj2jpakU6Izj5U7XPJuEVnD/EfLw0DHmu
/k2aOXjg9WQkmmshKsmtpZaamDbyordHFLVeWenvDXkDsE7z5ZRZA9ErFhEGIRXVnyBqaUA78F7+
M3/O6DekHweFJRP0znxFK25LK2w6IIaur1olwCAFoHnJrBOKHaWjdiJwmnGSYFl7F4KRcROfRuKp
EmTG/UL8kqFl6XiXPveI2LEeSoN4yMLeKuqqOtKf19LLSaqAZlyI/JrJ9OYPK/YR/5qazu5yQGMp
CnoumcIRuiqKqAUZK9FTGcU+jP5EayewPtyLxNRsqbcXRdHx88+fX7AqWsRg8ku2vmlRZ7m+rcf/
Cr4kpJOxoZEV4PwYOVL2V8HE7U6yCvEq+fAzRipJMDIYGJmSsnVbS+tOY5AaQPLrDPT6FTEsqHAY
SwURnRSb5nB2/q5wqllIJ5CfzIkw3YQNfS5+PC32N5JjgqsQ2aPMhHFmHRP2VFCHsLbXVLr0mEUQ
LY/WB3XiMw2zN4lq1gJljCpGf4z5d2As7aNgqgIKgOGCTJj4mA7wLTv6MrOVf9YQOBwpnPISeGVs
i372f5hBQE/USd98B5wzz8s07/WEn6BgLYMRZhnlFYRgxSFYC2jkxjvnG8AH4/K1GqupPJ4LDWQ1
WeanKU0Shrf1ScievnQNPRi/Ih2ribYy8cY9B9JtdQ7s+b91STD8j8ZBUxZibYvTPnLNAb4BtY/6
0kiJN1ro/0x3h5sBOvOPixTkHllLeBZuRLuhQU6fly9Zn7rU7tq0DOg6J2SaQjudGANELE+oDdGS
5DpGIarbeUe7hn2jH4GB1V5mJOR5QLAHLnS/YyQztsScaiRWWQWrpG49ykbeY6CB6mv6xVfud4sh
MADiGoZqVZbt4e2QU5dyBDfrrOVCMvuiJ4vozWYtwbTrFn6RYmsZ1x1FeDbgVI2Uh9fYL33cp4hL
VCIq1Jhm8KpWE961VxIvyxJwtJJHufQAxkA/xhYXKGEpm1GzlnUxwuXGgBYdoaGtHX+j+0lYwqm7
/EVswG9iWVj6mdV1mDFK3C0/S2sz3my0EYZeOxySze66nL1ArzYPedT4CiT/XNhi/g8WQfxT+YuB
s4+/rmdudGLR8F6sEbMwBjblpRKsJmaWZSgCczZUQgaAWbDy9A4kgssbZcFY2wFiOdXpAJMnBQwW
BjheVJWQg1Ty2xSDNYLLxBEXZg7HAhOyks2qFvdQJNhH2uvine65qwNm3KSSoDB695zmsAmt3Aes
wrkdBSh84WBtB6dRCqhAPS0nnkKPlVz1XbiCuBdgMRHtYpheGND/HWsLSBKzB2x6Dv5jo0gCmO/d
+iueEiwAeShKC8obJx21I3VjiOEDb/JZ35OHjvLY7qQJ+ZA1k0t1nw8ymzKd88ZqHzBHGdNsaldW
cCYR9XiO1fTBjiykqikKstKoXXZSBpd4TUxEbJtbq3QLSw5xyvATYBy8ujhCN+zmwJK8Sj/tA4Cq
2siCvrQGqm53u/5jNOL33SdJI2HJykv7mnsEdVztd3idnIFqmg/YLFZznVMN5iDXJbb/3hgend/V
RzuOg5RsT6Bd5SMtAbi6ihw2y6qD1CNnynNn8aDkYZ6OVmrgWZVLUQuzenrvrpzJECy2+WGPaz8H
40xJP+PWx03C7Vk/Jv7HG3PWN8kCYiwjqOSm1pKwRPoOjei9yuP/BrCjeE5gTFbmAsOurcfxzndB
9W657PaDTqS5aobk7iCGcu9nc2EhlpoZbhWIOLmuUKiyDxmYiGActokLDM+bdg9sSVIn2LtUEKVA
72eehAEoOa1uX4eSNSftGCsitrShwhRwysqbw+Qc3VNYW2f3Rb1y0BC12lfKZXspNM407lTRLaO+
4OQRhedBNH/3M4YTWdaeyoTrIQG347NlmLo4BEgzCFa4zAzukPTdXFo71WdFlEBN3z7rzTyChL0G
3uaWjJtXnsybDgWKM4oMyl7G8ehnh09M6UK0qBLaLDUAS8aIMz1+JK26ySuCuiQ0MzV9oeaM4R5i
vLC2qiU4H60gkKARADcan9kdiC4z6Ao5J9H869bYsSMaBRM0s/eocAxVYep/aZ2CHMkhPzPW5TF+
29MVQYsu3Cs7V1m9LG2nztM580sUOv671MEqQZ6gLSnk0OzfdvfgxHS/BmngpDzHL6txsRlt0xCP
Tk61tkDnDp2I7EzemFIBdHlve+1vLOD+UGP/M51zQwWYm0ipzufuZeYXtyAP8EBR+KSBgPa2GBqB
YsHfU2PNb+ksFHfzHQbhqukUbOOWr+WOfOLAG53uDvg4RrBbhZR2ZzkY0CWAsHiJ4XNv/B+d+Gyi
Tec64Zu8QTM5giNXEQU0k+4qEvR95bVJRrd2r04ethlimGvx69HCMLYb2hr7PH77mRb/VwfoIVlM
VEUSyp+pzEv+SHM/avMDQ1j5njTvMS7YDj15+puC5uG2UDSB7UmhafF6VeG9xT9X3eB+NzbUhP6G
8xGMuJ9bCb0Bl3VdX28brBjotNOzOQMJUAVF1dAl8k9OBpP+CnaumhS7CztIG8HjXqpta5SAyx/5
k1+rqWfga/D0K4Xs/Muck4QmWHR8aMfWhn1+8IQHyJoR/fDF5Ybb0zdir8cSx05fRD3eUiYhi5k1
RV2Rq/vA0I03brHOmubCkQ5yw0y88pCIW13tACgMBaycClEO0f8Rcn2PVOVggDwxAwf/QZL8sFgN
4YvSVdXVYJESHKTTY4uWBJ+QpZN1KxcVF2OLVYlHAsfFs5A/Ln1NacC2h5BMhU9cgUPqdy3JQYTP
GNJ87VDY9yLbAhc1vNiideiSa+PY56DPqkSBsR8O4em0zvgJFNpNf8e0ItTnKr9i50Oxec206yxp
9PRQ0J/5i7ZWIxKL1cUbbo9NBGX6xSz+rt0hx6TJilPSqZn7Webxa4wNPu2MVvHShg6lbM4crH0T
cI9GzllL9jgbbJ67+RwQE8oaXP20kZYilk70MCh2U4iky/qSnsvliv4ntOhg+q/xN/zMNCe7xt+G
7sdqnVJHOSZB/HNLn0d9aFvl0FmWBfoZ13lHywVys9wQ4wzqRxt2UuM8Iq2ddeMMv9Bd1n0/1pxr
WYh6IXm1QRWQ2wSsH8KZFjPpf8E+wkopTNWkP645sSr5oKBd+Pk66wQfcmpQPbH+rLMwQhkZiJBR
aJsyhkkmLAhgSgUc3tu1aKSvbcl7XJWplf1nMPZs3DPvsa0LqQkM6y9p4tCqMRPUQWY3HFOfjUBB
ldv7icrAXxW04VGOunOjjTEImbfGhDZ1/MazewrshFBglpyGOKFGRarXg+xybbfrLAar9YQptuDk
TYxU1/7cnwCI42WbLM8eYw8nm2JT9ImKXlmC9aPoIsA2XaeK8So0J4rhAxFsBKokhDmHXGloMxk7
7d0ppSuQS4CBbIbrui5yIijjhXZqPv4tADQAEwaGjwoktaXwub3p1PY94YZ/Mzs9zTYfgsd5+uxP
mB9f5QK+eODDZ1Mr3CFon/wr/7y7bxugt5n/TjUjMhBhyuHwOHeB/SlK32NeWhrU7nOJkVfs2cU2
R3wDD6juX6W95LCie/C1YVU7SmJUQQMwiAOXp7dmApYnft7hYKtJupuAcRhxxsrVcgzYToBbLFsa
exaeXd0JgFoNUcxb8QTse/IqpHBq8fAw6AjACBqKvEgCtzSi2ZBqHXr9gPzBKozCQ7vREUeGZqqx
lH5o9phs5snAXP9cEwIaGDN2ImZ+HJmIqkLyweZmbBGKCc9t2RPX+i3Wz0qOPxVCm5iG5QOtgNly
ghESAlXYFZo8siX/ZsZkVJd0Y+8RhdALVaAQ5Oe+a+Lcxvq3VxYfinm0eUE4khCY8eF9xZjFDpXu
tp9w4YMJTZsRFaFwJmFJ2CVFkD7nQ9wtuHk17aGEiEtmiCLVhtlSTrsNSh1SutwjprN5QS+OXBaf
pDPXamlRS1jTQ86vBVbXbxow0PIN+RO3m4nZKhVE6pnllAcDy/68SpeIaN0UM/C49Gh+WNSVwmar
0J0V+uxBpBOD2RG7XgZeTPgAHOYxn+wP7s/z+CZ40HryJaWX3OtJu6i1k5CCDJmFUK8IGE+0lZlK
FQNUUMMmKoW8EXPrw8hE4yPPMK4z4s1GoVnxXbjNvTITcdcaTRpoF1pSLr5e2INtWh/w4je2jIr1
44UmRQESRNm0WLX7/FJ1AeyiFH6l+vpjB/Ha3sqGqjrysTYg7fqweLVTrV0sFuMXPpo0cWJawyH4
EJRiIVreoEu0nCN+kGsQRj3Y7WR+wuALhcSezUtVq2Kn0a4ARp1nb4+5keKnCMHEB5ig1eiTT6JG
J6AwytgRFGHpHAT+9p/HhTh9Sbx5pAfNAgfQJujvpIeEwGuzXfl1X4ntuHFDTEcrFP4BjW8t78eI
L2NYmM/KhDbCmcXS7e+O+Kp3f6T9FzThaxBIHGeYgrnPmAzPqpovRyn64x4zP59iFnzQG0FROKMZ
Y8UmB8mkercYm+pds44AEJcsAkkO92NnJF8EHBZB5Y84ar/hDor0jiqtAU5CyxvHqe2wR1GKMBq3
uUk5LjrK2NejOyShTW8nfRh4R9CyZe69dlrv6GRypTgHtUXOCMEuGkBh8PfpX/qSTKevasbYscqV
prg9x8m1PP6h37ics6i+5fd8OSgii6OGYYTUTzzrVHUAG6m6Z6uJsogT8X8Sm1FZLZKgMISjXNmO
kO0+EwIJs2E/XdFUgGNsLibxw3kyw6SUphW7shnbjcKKNgWAYcvy/1Om0eMqjCPxDOxYX9TVqhsS
B3Fo5PkhbWv9hdFp4qlvqoyj8z+fDE1PMNZcDdkHdExkxHfxj8rCCwYWGif2mtQ5aOZIXcZQqATQ
3k3hxtJI/1VtFPzUSSO3SiUoOZXn2HfqiUCv5YJAY03kE2gXFGi+Wr0Fhm9c87Z1ItJoBblD1fQU
tx0Ju7Xs7zCMD62vY4GHQEuZDioO+6/SOY80xksruKAaqyfqcOPAajv1rXZHvcJUr34UnmGYFxyE
26bLdOWhZKFatrbJQK4Yo8OpDX+X8ojDMsYnhGUrly70O5hfRa2s0V9UBPupFoMrIeGUJdh1NCv6
6tJ/C2uSSBVt04cW5sdZI0+zh9bH+3egYoCbiAC53bxI4B0F6R+H2cHnooNQ8woDNeQLitxA9D/B
obwU8JhPYHux05Nyxj3OMqXiplHDICaxJNNBBQ4WGLZRdpsFQzOYwA77xt1ecXRapNbE4pqnbdzJ
2fvpqtbOa7HRsci8Il/VkevXRCtAgASrH6f2PQ1vVbvZRjjiLFFdLHn42MDBurZfBBP1HHkYKmK3
FywWSZlhutqkTNnxfLbfZnDDqpttW4V+H0gs8udp0yNkkMQkQ8IEfZhvNTvl5AHsudeiwC3ag6qd
OC+SoXZ8bc2MQyjlZm4cN3x3NoMzjUZ5TvDiKjHXYT+oW/eWWZQQNrCKIXxfKG/dumcRROfKn6/C
UcfCSMfA1addRMjh6pxPeHihPUsBnDqM1Q+07bXZlDZyZP8V6bhZSsGsmPlorP7tb7zPrwhByrhX
J8CF2dztPJYgtOqFhjhB/qokcAbHszD7VBVxYbqEXsD/4sD9AVjzOaxMGUsR9q+b4eyF1c/8rELO
4x+Pv+3Qdzi/WhHUEFgNNG1rz/GqZl5fkNQHCBij/ogoq5cEDJQxhL8te2KKzPOEPxT1uZOJibAy
5lgavK8p45QjvXX+1ENSddCZEPbgwWRfyh9lPZcThkm3KaDzjke9ZoZCcJoU6rqIXyDOxl3EkNBQ
0/LjvvRXNb6dyPL0CGfjj5H3fiNpsGmlIi57wmAYinzUn9n7ce5u58+4FYFKvybcdmp8TvNZF5cK
feY4cnWLpHunEe32ClsboD7ZP+fnZZyRr+CHVa5+FG2DDV39eK05sQ/vB1wKJM9WXxGWXZb2e4eA
ck8B8gppC8dIawoATFtTpW8wuHOp+JQXjDxYfym4Z9BrXeCmzq4gbHwt4xdkfO1LkwbRJYrbXiCD
+D/ImXApp8Tu1fGUnvFmzKx+VvOzb6C6OiQFsW70Hue8ZanZQj1c+shHx9XS9feYyEaldr63xn7k
THRLakuEi9zIXbmQsEUn1XPwsaJpsI7tZdj2tyIHadUJJZNPcd3x3ZoXPAMiLMMh/pqbabUsu4qz
Sh5UrsmMuVSn+SLEOMBR9bbh5JU8JJiprOMBB2XOsf+Cl/1l6/RPHLT9F9YplaTFl1p3NsKRJRsW
SixFKfZmHrL6MPbEpktsuVpcgdUahcn8N2gf6tydS3RQmaUw9GQUkt93ywy9y/Jj64Kjy06g8VNF
WbCdl0zMuUyyBxL5QztlujUcLPT7wd+GwmSF6G26bF7hpzzXj6bb+s6xPqEmC+DjM3KqvM9TP9ei
rXptJL+LAQLjCqlRD2NRicWfHK3wOIrNm32tGRkluC9LBplLBuVsLy9b3v91IodTNC8/uBmXVz/7
EGDNJMzZZPOUGpTvJUkmVdn2I9k8CAl3cBlcs+iUnopPGyzJ6BBDt86FtTJymFZ5kpaobavwrw1P
ZdRzHqpWgF63ACjORNtKyyYlN6zvtX5vG+j2mnc/bJLnmBI54OOKe4gBkJVmv4L1AlsBjJ8w85GH
WpFBKz9eZhLoKe6fkFzGwRgPZrMxXxdaSMwEM51vs+8r9n0DyQMRAVTNJo7jEOEmpJgzLeR+B9jq
snXxsd7Fs786y2r5HJaKsM9FPvYGjq4KE5fa1uEFgOxWIvIWwdoXSNFF6yZAXNgkTSZp1cUJhpdm
9kkLRSW8kBljVzQ8T5/URApqkZ+UehadV5XROO5yOcCrzQ+b4UtZaOmnedbytCHYgWeRHB1nK8tZ
B0JLhU70tyZ3MimfaYjbFNd9f/Pr5bLHH/qI/MgKAo8roCB57X6mw9iF+rKjrAQeXGRrFZchQM84
pbtewlrLTESvWzPeomTWLLDixMSU68vmooTtOzvBdha9UH0GHkvVZIDbi/bvjQxgSuBeoNVZPdO9
HRwK0WbD6TlNOmkUAR5B00KtHK16tbTF0boWu6TqPb6LX7zyNFV+IWri6bpwo0A6kfcOgXzV8QdH
VOui77qwzb08m1tlB65ZJY6RY7LAe6QcwFOKgB236hMDUl7Oi7v1E+OuCAa67JC3b7W4xMp5vXLH
NFqCx94+UCsA9MV1S19mSPQ7hZEFo3YqFqtT7ZO1tC3XP220+d6uWLuAVJ5hIR50twRNw8ZKvE6D
BqowtXzekKph2QwBFh3INgPP7NSSHkZ8VvZgFKRmeKlTyY3nNxeBE3k1MTrjKB0LalfKq9eucov3
vrVwKNVrPic7z3LXzUnYnXBh9p/IFPJvrY/bqlYVJixFAaAoRHO0qlxzIWlJz7fYg91RNYPfHqzy
tKm+ShfDFAezIDK8pQYSUO2KOaBurtJHY17Y/ZdcMg05c/G7YhJirPmFBKx1wcXdiSQn9Mji1r23
8tZSL6aHmHNiGHDK21Vh4+YRbApmePrYUm36Cy51Kf/MYM6qyjTbHUv7wwoB6CVkeJF2/f4uL/JM
zrIPDzQuEMITX958719iZCQqgYCPCvuPqyyfgE3qXEdlJ9VNYH3JRL1xVMnxqC/AbK4MPRymFTXm
EOx222FeS/K1U7SMjiEgwSoqyz2eU5LqpfeucZ79erWvb4AaHmXHMRPFdNbKl9xV8zsP+tKpxzlt
bfpyUnNEG7evx0QA6cr269f1azKggL03k5aJveyVPAbkZ5Tq1JdVGGd/vJ/3YmMQQntl+xRKip3n
X9ToM9+RPJP7Gr7BK7+4gl6azUe4ObjBoYRen/tfD2HhtYkQoJSeSeUY66zqcMDXkL0plkUjYgYG
RhaJ0i0ynT4szfPlErd0UamghohG/AQCubkmN9XAfo6TFDO/Kd08PJrtWQhblVG1CDRTLmM2qU0f
CdSw6ew0XoB8SA5yfAKE3e60irLVsdWUdtulNYFpTY8KBV1WyUVgcmCpj/+OyDevyy2holcGBJoX
EbngI/FeKPKf6kLoa3vPjRpT9P2hezGfj++IWR4mFa4/XdDnfbZDJTQjBF269g6i596UN66insxF
icGrqsI/qxi33O6kZAwjajKhGptlIOJkuQcCh4R4ph9zDZSu1oPa/D9PQDYracX/vuMT+3x516mf
+9aaTpMIir/JKXrFNyxONWdBckYxGXYcJ6Gm3BvvVW3KxW6T+eTRFAxejJzw6cTw+C3TWhqHTpyn
e8SWzOe4Vb6wvYKuiFR4XwELzzkIKZvjJx0NnqHYXJ39IPd+UyrZ23/SoYrPVP29zkS5P/Cp9jNa
hIeixSHFM3He4GpubWcevcFvX/dujU1vCfgLNYJHhKqoKlFjnjo/PHb44E8Wh38OMHzB1gL3kWqj
KFH1fed7NMyK2Vp3niVQ7jRF0PLGVaKjJV7rJqufLXeEh9lIY4MJ/sZGKM/Vbm623Zos7GkTctVR
pkN54N5qJnaVkxu8K0JIPt212KXuxX8ei6gsxzCbfJkDN/JPcIywvdW3rYyknJBPOfV3w2BCd46v
WA8xj3s6s1z2+6i7qws6F7P5iBSh+bN7T2NGMoS8xZdG8TXugRqJzV4a+lq7csg0xzn69zXFpLzR
2OT+IGalHgYZ26EQUa9M6dEUkX4sTsh2twRhw3f85rmRzXKK+9yGARmc4Q3sqGR3mt8ewVk60wT9
YorLIVka6ciIx+NNVI1DjFQyolFdCbId440FUd/fGQyW+UkaE+4yPA1FYB6y2Oq3JIFnHyaFhn+L
/CYLYE09xl+ikF1xLjntsh1Zd9GVPy9upTUaGOfpvM+FLoCwl5r+osS9iYW1E8pCZMffGK5FzmJG
ZE/LRTZlngIME9ErTkOUQq80s0i2a47+g/5L+XXqNUQhWb9nUOUIj442/ioSo+aFzmP4T97++HV3
Y5/Pm2t3MMid6yODTSE4P/vAP0AmVEEgvIY1yfcb6PtE2VYCj3vq97Ws6uvfToP63d3pjKJNUnK7
eNuvAru0Yq/RGuzBfdxkuFBsEbz/JkNP4ndMuHMWyPae79lbKvpb2LUP1IRtmjA/fsmssAJT6UNm
YL4X3GBotab6hJPMFmT+pr1Or9OmZNFhShk1c7YZCiNqupVYjPGPge/fVcuMGq4skBDFgXn8Xgf8
sF7n1jeU3Mp42Yv29PeHiANE/9isC/cLlXOQwRzVl/pjuLFDoxhKO8OunLQ93bPYEfzI3/EVfmvy
7fza/WCwawaoPpq79ueucSjBPBWHkYCTSae+62Z4VHopBE0RsAnw3P+3G2klUpdVcbEE5fcqEHxR
BmzlVBaBmACqoBiD5sugHvBZ9yrk6pgl6Iwx6RB8la6T84vu/KjSl8dx3t1QoqIDTLX5VDA13JeG
vpU9DD6CXZxk3hTaBw9Tf+EDGP+aM0ZQXoof5TMHtQ5l1QvxubptePdWaEkLEfjnV43GmkyiHlkK
Hl6t86eBXcS/ww+66aDdS0FXvrCnhgaO+EQymWyeRj0Lbhbxi2HK7nreBtqaHhS3qMicBYoKB/Pw
/0tyjNcM6oqbux8TI4llaS4K7ORb2hMdBvkMuziAXKdbePIFdwsvYSaQm0AKU/lkbwvlqG74rZjM
iCuqf/S5rSG8NEkDWn0uAp9PY2pgw54ZmDJ6Lg1ptXFZ13DkPwG6SDUQrsQ/1ynExqZccMVE0NCO
5B9kDzM1DjdKmIJn9RoqA4pHT3eq5rRNzhxrN3dRH5kIP2IN30bry+CC0ht0rqkNAMJeDoppdqJX
lW+3ScJdq8LdezR5762jDPyC2RA7Y62f0kvuByHAsZSQd3k/lNgzlfJSr2qABzWjdhwFJphKFQk3
sac/NLPzNAhN8cgQZC6V5cVpvvGbZykdvrby94ibPhP+xEuW1tnQ/BNSSMiNnDsNJ2d7YbNn8cVn
4YblplLM9eIcZo8T12yydHyT/yk8Jtd78yTB96Q/glbG8AVhNpvzNG1k7RR6y+Zi7672Aw7SpODT
sOe+ZjJhWxEYv0JE1GurooBtZi0VR3mVmHq2yhm/2NZ7u2g0WAiCMLOxIf1jF3JdrrgnpbbEJjKl
ngMmrRaARYkROw1eSGrPcZpH4Nozn0JTqTT6dB1D+QafYrCSz5kGhCskmn6FcJWcXQSs8qbPoQnY
NDsARSZ9c78P3lSSfGgd7qJrBaF6cx5KvBdfOpxY+oGA6y9Fa8PZQcS1uMl8mD7jdgr88gsW2yg1
9CcutCSDyq7ZcW/F1oXAARcWppmOLRzxyzMk0CwCvGP7kfFmsQois5yEPDlUtyb+8EJ1JnRqHAn3
wHvomvS1GOmueAAd58PAq4tV4CHswWcL9HhLfDdIuV2a45LjtXN3C/omKFb7CHa4n12h8kaD9lce
WxrDK7XKZ2LDi8Jr5RMjgTWWvUe3GmhLVpbQ9wf7u6O2ifIgl70zgbw6b3pNquU38ssH/uvkmd5Z
zitUbgB4BrWgy6PO40bGPgy4FCWK1QERZ49QcQ8hceoPhOl45RMaX2oamoaO9l+j1Kmsx6nyH1X8
ZsXy7sZYdHAFtzR9Tn7vvNoVbeYliJRBjKpXyGNFyCdHMMMi2NZJ1dpTBRSKoagrRiGcaUbN1vjJ
tAlHBpgEnWoSYEm2s43gMXJwvky1HJhlDt8iTAVmXkOBwxpW6s3Rnvg4m616r1hInh4AvY5gllbO
7r0fm2ge6DgX5Qot3KfL9wzcRcINfxpT2WmhlBXHbl5CQY9IuNSXHX6jBTx6kYGu8GFBvXLnkf+f
SzZKchVtFiqN3ukdztyrBKLsbGLbNuuFhpcKh3fBQ3t8vvHjWtter+E9uZYboPIrGisgjNfJEGHr
i7oaJj16G+Kf8K+n1NHpPGwl8upz7+NsuP4GuRhhnVYzjL66wfmMEjErICwpkOBmgO5S9+0qQOD2
NYv/yrlVuLMDPDsE+cPjMm9+YPexE3aVUn5euiM21ea2jOO3tdmh1StwUQzMLrnSNMDGQHB17JaT
dfHMfvmJOdSSr74mRHkSf/B71BQU0mmIHJANmdgUpCjbQ3wAExRKsYS5cuI9sMYL8ditxbaj3B07
2f6yEPW+wHYO8cf3OKPkWPTf4VEWmBOOLN2QrRSbpZu9QfGLPb785vQiEgIPJPoPdcQPr70KpECX
GrTPh/kJjAYc57TWc0sIGOr0/snkZvBX+b3rP5JWn0fwd4g6En9MgHoxmyfe5XWquuSj+IE9bK/h
1G3cO+ebRA6cykqXssRPz+XAcPVM1qrYofGG7H6AUAjpQ8tiuHXksurNgJuS1+CkuPvu2hIwBivE
jycp/Qj5p+e3MvjpZKu7uXLWu9OBEOwZ+qJ5xPsEikZ9nKomWEmxBU3EGH10fwdUo+YCfF2Je4Z8
goQAPbp3xa3XZuZQJM+w7AUWByNoah4MaIGRQA1IHRllmfvtAaViVctmxue+MIS79hW7agKCsaCb
WICMPunV/N53vDmavAFJhqj7uRiwrAAsN+cM9PR+zsP05dj3aHrf2po3qcRhaOWj7vJLDzvnmaBo
BCgTsddrjnEPeqKkltNEjjF4kPUxO+ZpTyTSsxHNaG+GEnwox7bgrXAQjSzUF3loAY+eO9e7QToG
qMTIBb13iaU4M+f2ghDw7E+LvtYswEtZ5sUFMK640uDkdARw1RVUgIGO7DklEXl6t8nTFyF9C3/P
2QS4OzLncru/oTGJ+b+XEk4khbb2sZMAkeWgSeYr4lHx7zZ67Wa4J7QbQRWFpQRmlhHbaZMhblTC
mKd8t1z52sQRLADCT/Ek2eV+AqVeoWOVlO2fXQ0LKKSc/PCQcGoH/gzc6shZFyQ58sI6JWm3vdUk
vCUNnloNNHo4wPlMGf87fZc6kcjwtGGZYMqh8TAkc6MW/rgdevEXT9MplNKZIsbzCWwgh74G+aL2
eltanAjCkRawBx/TP+uwIe7d09+sU8GEWOB8H4atPBSBP7m4cr7YLwEpM1PnG9eVTxVJpoGoUsUk
e1gPtWITsssbge+HGavGxpxoYX77KXCr+F1QVOnsfwYJCLq+NqcUvuQpa9LCuY2AsI9XlIhpWDEL
tLnHDk85fNAKqXfZtHU5t4LAnADDZBdkxnhZxN9+FJ9XaHVlGUjUpE+emnBXL3+ryYIHA7LZUIuu
mMUFx14xYmq87dJm+FzKI+83WoLxhgYxcxtEcLpDZjxEBYT6tMwxehjwgGp94CCOXFGrhRXwS6qY
Hc7VJkkHBtFmSUQnheDLDSuLYOYKm7bKKNrxFJHZS4kcN06MNUDs9KuxwdNNM8Z0Ae8KPsoX+NTB
wDrLFjWZquAMGIIp410h5m+VdwhrgxHMdCD3TMvPvGcllZq2sL4dWUhIWmmT/FXJHE+wc8/MuL8/
RRrvFaiytXpBPZbnXQYA22HLMW8q8FtgiH97/zasESVqIEqRIPshcCTv7l2yK/a2l4W+F3TlUrY6
9+IMMIxJ/1HvrNMUKJdbHpx1eXptvoWQZsbKidSVbtb1G27qtczu5AuP6HYYfVgCTDNjHDvo4wtN
Pcgn/wt3I1Hu8Pgyc4HfN4bn5wJ2Psd7RQAYejpY6qSWkl4QkyBwFY2HHFjrmHyhYNiVIZUQZfvD
dTpurHbjiW5QRjk2wuPlEEXYwjDH6EgyWU0eAwN7XSsFosC6Xfvex72BTLK0qQMZBh36F5llIwcj
6+Zn2lsL4WtGbUB5BAcp++2P8uW7syKbsr2MBI4ebozphKEYHaihNtRnB51zKfEhz474aBltURXv
lfl0j7COuB1JdUHoHcAjwr40MxAFmCNrGVX366jYjPNWzAuTYNBpRSxWlqol9YxRTTXQWQ7vABht
AZA7LsMxonnRuK5A+iDpfr/ycHVXO429efz2GoatT+0PF0OSts357mXFaBWjiOq2TmEaykqi/Qai
O94Hg4gS5mgQHXmW8nheNF5SThD6URsMLTYhzYnjMEpS9MNGsTAqT0ReQ0MOUjx9d/uEZRA/sRwm
PvlWP0xrf/IUL/xAnFlMTy3o1fIRODOf6C8L1o+FYIKd1hEsYj584i3IaOgxjdf38pmpVlw/nnMk
jEGPACy69hUw3C9IruQeIN1Lj5z52ccKevFtAnGCmUp7MZHxJesD0ENCFYE1OSivGpnnSBcZHKay
iRzrvQcRuoyAc75uCM3NQqKGS626vpCP8MdN8QtUNfgDW2E3D/xQkf4qkIWU/SWx9JT8egLZ7NzZ
rSe/pOSVWUYHAVo1XOHxB6zagHzMWyTx8654JHOgr4O6MDbj+RFfnoFuMh8R32Mro3SV0tvf27Xg
+5mbzx0Usegq6iEt9vzH2CGL3t94nz09lFdlu1vNwoM6fNrXJZxG7A07jtHFjLRYkyUHYjBaUif5
yK1/BwAVcqVVU1G8+BH0WrawaX5HdpjlUcuVK0s4wLN8Pqh4ToXZrXHi91qdf0CvAG6iR/jUJmUe
SCA/CRz75ZieDjjWjPkjnUKJb9pKdV+QKbLTxmdC8O0UT5Tq7mzpu/YGDKBABFVMLM8uWbgcGPSD
27Day4L4QgZKhgt/HPxvkcj/Qn2sFmliKvvG8LqkOhdaSE+zaXZr/dPLXHEYa1wSGUMLL9hOuQnG
AU29RUeV6zmbN7sutp4T81Q1og9KJi7E0b+dcwLBes7YXWoUKXcw/KtU3rUd3oPdu7Me3izETSHY
xekukS59cM81wXMxVwnpBmKTyyVRDSR3f71gstkbHnaOSwUGuNRVavhR5ED62KbtA0++LqR/xV7T
L6ekrEzTyUBg3P8SzlxFM09XOq4a774CLIikD9/JJGnKQ1s7gmxo/vRxdg6UVJUGmMQ2/EPWsWQc
yysNNzI0UJRmg1b67im+8XVwRVAEbK3+eBJhk69DDZRtVc/JQOmITGUjbOdAHYIrZfwB+QliKzQN
UpH4MnqgAMB2h343OLjf8X8SZDTPOY2XyV+2VpBj6Il823460SXE9HC8KT6wbeGR622VZ0tkv0h3
pf9cQu5q5Jz8DpyHjH5tOp+n8ZajKYuoCiS3zvH8AfVOap6CTM/wBFkqaEcOQw5rD7kYYyjz2DLQ
LzHDu9ExWIGFf64rHagmTk5ysZWQw3l6tVduEzTyoKEkkOKjRbyKIsrjPbuiuymvI67cMX0Z6lOq
JvBCSXMQ4wf+gKoiPmCyCpJHHrVrpVhFfa3jNlyoxkqIRsCbp4mbpMFXA2bqsF5NFB8keZx2FMst
c+H+IlujyVAcGtSQ9ZqeO+hgbW40oSEt5IxMIaLw7TCKDeD8k+M0rzMOMTCZENt0aHaqtm/myrH8
OdJEU0ExSFW3ppux0BuZufW554Rh3J4ml/jj6wzpiOqaYfbGAWI/R3gdMrhWfVsrN7SaAQRlruPb
tKPY4pNiGtMuHlBTwFbcSO7lvxxHtGvAtieoT9urzeTtWi9ZY9u8Er8m6YnALVJL75DM8n6jiu+T
nEuuGki88d32tCd5XYUoT/TLdB2/COHfBx14wk8W851Dz8RRpuCwjamTfaPFRZxOUD3nJt5A7NZ3
CJXQleu0TxC/RhaCwQV3gXzXTOFnw8aIgHR+suPZAfbXwJuU2d7W4Nun24ORy5Ho+bu7H8Ub14zK
s4s9Sb2YPFirXQfNk9Cbc+rU/4Gh+noA0MwbByBhRdfP2cYIspswz9LFUcV+NCfeNpIoV1wN4tep
e9JUdVFZEJySQTWRaVPwbyAmqz5PwcqXsL6durzGxZcUcKRhJaQVx+3KLGtij4CDatvIutMdciNj
dSvXpIg72MLrRyL36cV892B+PD/n57sosdDk8UwJKiXZ6VakguzBji+SWA8pWtBBARSJENsl88QN
msAIK00wa59/RdaT7Vg1jrsbQKBMC0PyLC8T1GKzLJgnQ/XBWFwlCRA4UHCClFSzmBEaAcjQCKIM
EMe94ZLRWUJzMS7KyMoGrZtNF2y2m1tgo+/Jx7MoPJ6qkoCd4Huy7XCSKiqauWTMXyS0LQJ3yn2M
zAfWxSdGTKQ7IrREv0cspfax9/9Ll/tf47tBgz+gIXi3rtmwGNOsZ9ZMtNlvrklPkzfQM5QNrVxg
1hT1w5FTiWwOCSbn98MFN3o+RwK+ERcs1Df0sUlmf9QEBWHMlvCkiF05PiIEcQoydy1B6CvB6SFP
V1wWrc/m4HGD0I7IHGcF3dk9O0R/HwPEnmLgdlQouMrezzAhWtdTMauhjuC8Y+2q24Z6AfhpqEAJ
zmOADvLURdJn05y5Z4Kv27TmkYnasRTP+i8b9EbfujM84R/c9uuUiLAy4CK/kq4lQm8oUgC5VOAe
9dwy2WH5kByDZGWKxnhHD0DJ7OHBB1mT1QCcHHQB4wapHgG4Suv0fbGKKSnjDngRrnxPR1ssIS2s
0FMIkIXsWN2m5Kg5i9dRqbQ6YjEVmQjrR83koDZ91voKliCA5oNUz6mdWBYtH5xr1sxH55uNgu3y
VAL0WuAcPnkv0+OUtkQj+z1oMbC6B7Y8AMtI0tejD7qd/HsZmDzOkfQM9E9AMmC2D3iwtIWCbp1a
2htAINXWuLWzppihoSszUri0w5Vh5vdg4KXVl9kyQtphpkpvlnMcuBJXUG98udJNz8lxgEqUihs4
bJfkmu3swgIgUeVgdDrXhQZeKB8fQwrT80ukbdj/gv31WqF0WDyvwlKAFyJRbYCDrTWFWx4Ahtvi
RFECofexPc+ghZGktG45xml3pBR2nBiZso6Tou8bYcYfI3UVXHroRpy/F30K5scJhSZtIPFKfysH
vAVb4uPuTp/T2ZUkt3XJ0miBYeqjHpb5a2WW8znj1PBpZDVMWxF8guyPw9+3W+urnA88ZzUXdc8q
rWc5l4IKYkpJPkgl/gzz92p3lUB58tOf3AoFOPrJc9GQhSYefsceY6g366dToWl5MUZjUy3uXDYc
eIQY4S4x3pwtfYGKsZJ9pkesH1o93yWN9Z8soT7pnY9gdjxbPjf/SGiFb3nqzkT6qwSRqmQAZdiE
Omj9on3ow+shgpB3Jq9rCbjGOnIV1MpIy9TjJkDEyyqtsoeRDLK4lljeUp38Vu7+RRCB6rIjI3g3
clEjmIWo3EF5nHSSJKUsNgRlPjUEKIarwtrdn7HRQnsswbPxolvwfE4k0fWk5lPmjZgi5m6X2wok
OHu4Vr6hfwMp3EQ4qM4zz3ljwn8C+7+Rv+i4ZWox3F6MhEZpCU6w82dJsCDHE7xL61dFLO+IDkBz
+poJkRvyiGqCDreLw4x4/CnMfW9ISjCs/GDDIJYtJgkU8K9cio1DC2dVDoraywksJp0VGlXkLR64
gzFknPbyWdS3X4/2cpn9rkaGGgpr4VlALHahCfg6Agww9mTzA2J47KeNxDVEhlU3NNm/q1/nnTDz
oQv2JhArohdvT0UxKTcUyA1fkX94w6JpcQeVMmstIT0RR3fj+0PXREXZRIQYt6VxahhVOcopEGrG
ClgVOd2adIkE0SNhIpw6/nZOzPdY3pRFm9b8vQLOTC5srjW5YOV4DYKoP9llB4EAolXaGP/O3MaC
7ajaKtkyY2F8JZiIWGDXh9K5UJ5FmN0y5rwHYTIuzGCk8AOF3S7Psu/vkBEwv3Ey5ec47CRwr6F9
AHdH5t+xxRaUsiQ1nb4IXn8OfTs2YZqg1Gjrv4GmbZK7JYM4A6aUXrwWm1v8G0J5w6lnuAxakBA/
2irdlyUyOX+xWmWu41rxwixqw8otx9KJ3BD/N+VSBMTPVBtTMpkuFdlFSQJXBIV0wRv2WMtRrMO1
cBobZ8/kxxj+VGNU/RlwtiQ2Olq8GgYNudIauDnPyMYmQTUM4uxRdTDtoS5mW/OZLF7gMEP0X4e3
cSVBWD+lGlSD871+ZeaX5s1ZqL3+SZtNZ91JPPUG9Zl7wdsZAI4hnISGTBLNlSy26pBDfp5/hlbq
GQSG6jy12PnXf6Q4tBbeOlEk4fl5Dw/HtTCZZr4488hl70+YjGWHjyjqjnFtyHow8nUI+GnQT328
ChHDRgkU0Gja+Fr6CXk1/8tmKmAQSvwHANaYnEZ71/7O706Ia2qTgigBJZ70DGBCaRBfKx8X1yxf
h2Zwnn+RzDsZk/IZjZ6UHeHye8Hq+XKbQQT8LHTIBKj1Bxft8K/uzuj5IFr+UckTJn1pBFo6hCq0
QHDRMCBcHQRiVZJWQH0YOYlzVNuCV+7OWY163nqvPq0QDDSW0ZxNfFAZCG6G7Ou/7lEEeXp4dLBx
S2OcutrqpX9JcWrmt8cEl/wAcH02yq0LVbchdSnBso+YNrKx7D6yUJxxxST2Ro6RqAkgAmKpHmqi
UHaMP+4BdCjoWqGrir99XRcFqdFKdYrv4PTwpzYyYZO6YybRhT6LBfNskjnd2d+u1stslh7aAXvh
zxyzhsfxzTksDi7YRFNwL2iQlPfKqGfoPtiXzptRyBW0nFYWbvt7CSWotufXe8cKJRNif3uXEKVA
JF4YgIkd1jGhnS1BNL/v0d7LpyTgaOuKxmEj5TodnDMQlr10KAM9riUTux3dxTecBM5I8gfYunR6
H4D3YpGy+eciLK2prTcnLKlWa3kcPBfW4jwDgNfLIDhtUjedMN63BiTPBgiBRSoN+9lcaKvoVW9c
XOsv3tT4JC2HKVq6hOOKiZF3IiqBFRoEci98U6mx61haL0S2VenEayxzYXS2QKl7SQEJCfRE4T+M
aWGi98mCJ+UPaWnrdnArFyh072qtkdsF2xKEhn8oNBUej82JsLfl248Z1NUTkmblBpjwDqmcBuiv
6Ox/BoW1UwfgZprTE5SKDTziBSrFexnwXOlgHCU6hNbdmxnqks5/C28rH7Thy3meoVRL+r1TDe1x
Ayv2sZpoWfGDzbQngC2hs3LhKC0jDtc4kn9Hj3sKZMFQjOHZoNHmJOvQr062BbDWXTxPZrdjbBOv
C5PF0KGQVRMBSUwmSjDXoj8Vju3c+oJMKycyVhHqtCtl/z5Hb1+VYBnQ9/jtjyBX/+rxfCd2vN5j
0Xi1s6rHhxKu0YY8QknwkQ/ckI72AbbkD0WnQbyjo+btA+rBf/cvgflIvj5tumMkAexnzU3loxxQ
El/9BnKBYxcAoz5t2XURhFo9tSN6n4Rv5JeM7MmquNphNnWR1S40KsjbVNliORGJMuEozOzjPmQt
Vpt5ymaTGqiaYduJs6D2MEfwH5RCvUBx4mJjjiJHiol5O7DS+Ig/tAuJAwfgGng8+R6hOXWv3O1o
tzc0sPodFLeO20CWnVzNSkpx4LJkJTWKHMRjZnS2XIkhqlSgU22gZQCpqtBiHglSjz6Eihm+hMN7
10ncVL+5AZDkt3MOf709B4L29KLuZLUGG96veXZZVZRLKr3ggfqr9ghTZcvpT8l8ERv5PWTDq9UN
5B6nt0050Q8jF2ZHUJ52Nyq4wNZAMKxQHPn7REnBtCWzP59HnEtrcR3HDS//COKakMcSUGWc86L1
kVAqmzjC+wU3A0VBNNOtxuWJsg8GiFD2b1bE3mrSmzT5qORCdEdI0JY+N7iRBpvb1ubTIhDGGQMP
8ioZSWk+WrY1v1/YuesIbdaWaZbUYMXAaZjMCDxZjxcI6TVatCT9DMvKakRZKxpAtdadpRk24pzy
NIoBOB6+U+Aoema8Fs3ygvieoyBK5/ikn8Oj3w6qZKd7STnM7AJBB9JAzkSWO2us3Gdx5JXI+jLF
kgCQSpfqRxfaXpxlrN8+u5nHKrMlLsTjUzFrchEB0ricnFDOwAgaOKv1TPGSyezmTIwxepU/gXDk
HP4W2sL8B+jfgLGsy3WEF/Jfw+GRSDAimk/3ymr7x+qtOh8M4M19qnK15RsLpv0pyVUF+UN+zhV0
0aQALW/FjbezjeuNEy/uiRjxjS0ge1FmQWSELgkvB/9ntE6N8Lg8lP/UK75JzPl1HivqSHC5km/K
lKLF1QpMBWuAC1oxjrihwk7JZgAqED2EBoucr5lrzkPaxZWOcvGHCRafHF+TkKS7JHoNFFLsDCFX
K0A4DZ4xsotGwh7UbF4I1zoFs+QQSFSWmLG/qVVNqhhjwgezn50KT7ioY8uccFVjofk1HVSXMtno
fejeVzzjrNi7JT25XoDtgyo9iadASFixvOjhrjafZdYhldxow5w8dBdG4SL31CExUFwmSDLBIDby
jDCVGajWCzds3M56lCjqeSJ13YEWHWw5kkrgRZSPUPfuDF0mtP8470pKUl+yYBMCwI8pHsfAbGJ2
SJx9K4a0HLGoIxUzVBOMfc6nbvwFBxqmuAi12PWg9EVxQEh6B387Tv5XZM3scooL39EOsOVUkQg7
MQAvKSRsRFJ2b+LMcx5OxL0o+UchR8yCAsPdjQlohedpgvLXeOfjzPkVo17jx7vCygk418kNDI4P
S48iaplZ9yF9BK8jrgYUie34VVeNdKbLH/o82x4vQ0t0M8yqXMkqLRfw1dYtaHRWXiigg0uxiZ+n
1gXgy254PslhBFnTUonagayJe7aiw0+/l65qtt/vVhZE2dNq4qGmI3NttGj2BuAo88jhevjP7VO/
hFb1avT2/Gbhf19HmwEJlCrmYunUrCFRCiRto5nofaaa4d7G1G4NUG5RPjHKUiEIpjcrEmDbdROY
7XHKSkEjZJRwzcFg53Nu73HpZedBdipCLPExsUcbN4ztlmWnkjkkmhISY7hCcezzSN6bON1W/h8Z
ld2TNflaZdJ59PDyl5U2PhbgFRgBr3jUKTvBrSibT+KrHEizqrR3GXhDx5hU4mIFOxjuXBIcg1lr
bEYhUWcJVCKUSkFoOFDYFXVVDZJuyOzVeA2dKvoKOLJvki0VMysg+75Qhz9laitXWZi3/SuDOyoA
WqvlP6QvwRCRMaA7i4UoquQ3Yjytp2zWZOKOu2KQW0Tzw55VJRqafzS3VulRQdkjA3ozO320YgTc
NIRtMjC/803tcY8pkbwQeukUeGaUSkVHYz1mKS3fuXVE/16NKAKUc1p2wD0/6JPIqDk4YwaUk1Oe
8fmXlFs+V7Hje0VgCWNYpshifhZTMuUjT/JdF86khsgotC6poBcrlshkuGTmX78iLYR88A8yvmrP
SsFObvSvMrTR7I8QK5kn2hzwfXuqr1i+mvqNnr6lL8Oowa1BeISu6GJeKQsiYHWu+Cr81Em46qMQ
NrK10Y4PSk4lkxSUQgqBQxiR6IvLOcvhvyz/wwfEqcgmndNlSJTqRm7r3izFL8NYasdknLzuprk7
n/M0s1jPS3J0/gPbzto+WqQH0ADjgs9fcVD+goaYXkXR/sx0Ez0XSlf8DPwjGPQVCas4bZBvr2F9
/1JjaOdZYNM2hUvby2ZXq8AnxO0EuY0Fn62yHw5IRs924b8VmtiK7hxypHRVHOjE/u8qX5TjN7sG
5/KVFNXLZVcSAIMK2WoqcWZPP/5X2GJieyV9G3kwKYgR9gDWKlN3Y5xnOF2pQlIdZjY2/hwQDX5s
CX4u+JKu9zy5B2FJ3nbUnqVeAQYhc83Wf5Qof5jZ753bSi2uvyt/qtU3z8hjwaq5GAZscqgLmm4/
RtabUdRfuFBU3+ZW0teZgYDd9ibmwezR4vmgRWaNibni5BbRkXySkAGBUJChQZKhjKaosPVaZT40
1Ial+nvej7icugzYvE/NZghnkoqtynAaXtozqHgjPIwE85ux+YpihfqdRpJf9BrX9P2HRYXpRpXY
2kiqu3+ZsV2wRWRAZSh4Q2Ljx7m+BcWeu1bdRhaWHfrR0tSO/Y8SsaW0JOIfWL2i3z+cNCJJOtqH
s47x2zmpLICOmQxdh+C56eC7iNfx953m+KUt8cLX/O6A1lf9abyuKndx2ZsdkZB8NngOrIZGqPPh
kT38fRkeich11rLTKJAeWOwjV2iQ7btS7WnGnvmj9ohejkRSgw9h7swsd/JtrJm89oIcDdfadLoz
HClJbi/M/FMt/nuecySd314NeurGjxsPg5CJxbi54KgmufpRm2pt5VwYrSe0KBx9dM0Q8/F4bqZT
GIdLNmH4aVAenv/FEyX7Wsn+ozJpr4YL5P6gxTjbBVKLwkNKcahadA7KMIwdNVANdVKRocech64J
3Eei5WeGhwWfWv5jFkw+hq+pgY7EncukmzkLfGAOiqvjfL9kKtAEZ7M+fh5Be3e78WvrCGASE5VB
aTdAuM/ZWYYYHHjXTZIwGYerSw03cIk/sVDIcnnR/I1eW/k+I83j7uokw4Rx/dlMNEwBNw1PyDnI
dSnuS29eCDuVUhPnWNG154x1eN3/blJxaHEjkjEkdA6whkwFzbgMO2oaemyX0A5YS3R0mFCoU9Du
Hs607tka2/cho2AehR2X5R5NHUi0Cq1XFAtvzuENNyUFWsf+YW5u5nlxP5RMfmUgmmtcT+Z63ydh
tGJeayglSDjnMytNxMWqrtWmySRc/x2McA5U0PSo0R7j6w/g1zOps4J3vQ07MN7y61m8l41qMErd
Wj58ghy61zECnun5KUf9z6B8ujRLHP01D1PHeukLJlwXaHaklf+W5K+D1vTw1Yyl5n9eAtXe/zYS
rvmV7Gagcct8ccu5yjmBcXrhCZWoW6u3BNevqncZh64kO2IKb6g6xxCWHfkIlVAlbnbjpcf/21JZ
eddVWJXw6PzhHDwIJmIHso9MVoD4/WeAXh2rLz9KJ048WTJzHQVj91sdoNCHEJr/GylC5A4y9esc
nPmr8wdd0gdJe6QmTmhdfGZ2OHuBbE98UWuOYXB+IWM+DSJ3lwzmtzDLp8l2T4cf4jEFsQOBng6B
xppDX05Lybj/5pZEaz1bL5lSVsFzegp+n1DpFyFMq2I+T8zU1O681QnDoaHLC5ug0qOlemff4GTv
am10+kT6sq6fF23iF1Go/QvK0U7aX49uX18a6WfT534kpVXPGvvmcEXo4i5uuVd6jd/JelpleRDy
Drdg4txzUfIu0jMSOUN8Q/XDV2xhwn4cLxPGgRYS2ezk3fx9s/VNE3HAoq2ew26fhuU8fLn9kgMw
DB7y8PMyzPmd1pvpX6WLZvGrfW/oZrt/otYQECKbvoSvBQcTuRUYcRbvPzZZ7o8cvrYkBB8scRo6
aaLNmt2BIiAIcHgIk8oKbPGyF2EN6RtJZLA1L5S2MAuHjugkueRgMCqIp9Z/EnyT1sTeyyWPb4K3
uZHEq0M/ryGkwDkYeSpSvFGdL4OL8hX25tl+k+00r61EcTUD8U1zBGj3e6fac9+s2NCHS//JJp1z
EnCy3D5FbuYcCsMJedWUo/fy6MxSJ1y2PeZZYG04KqiDAd2BYN94NRXD+Km/tesuJJprUlvQrnG2
NxOAImTAT7hYoiSE6xXmj3PV/25R2efOYWcpQwwjW47U2PnM4zKV98h3rt75Vl7KftwZWov/L66C
BMmNnD7RmTkTbOWgsrFGSpDHfsd1BdLA18wDXhG+Kgns+26jiEJLnmwnLB5ZF7UvGQReVISTOfRC
U90DaZGHVqPg6Vo8hPGZVKgHTdPuQ6anJ1LmPpc43YaUzWx1jyYf0TP/Cql2lN+qQy2pdIWfPLPL
1PhkErGGqzh/8rwRfcq2j4PEtEyQ1JkIk6ki0etLT0zj2WUIKVNYwRE9FoadxRur3iunBqSLiJqD
eRLMxTenDyTI/m0xpmjCaxHIQv4XuQ3Gqn2Ht4113mrwhRdJShvsgDGOrggIGB1knuOL/tmzpBHJ
RhE8ULH1R+cnWmsph0LDyzO95w67yuIzl54HfJnJk/VDrxHWc/uqQRlVX6lifuWO/N9c2KPzxKTd
paZOnQMhzke67J6oFVfPuaOZIawHtMz73ICJ/g4dXuJugueFLZ51wnO4z/j/dxJ5Mm7ls8ATOPaU
vHI7X+S9iEyxRE8a5B7T3FuZWkhYDHIPiYY6LIzOA07htbbi2tdWCCQsn1yjoBBG1wiG6OCbs4BA
AAuIaM7g7tkVmGdHwJXjwN/AZQ338OL4KgOy+DKutwTMiCqKZMAolZLpH51C2wqm9Kvlc3MKjnTj
DqNdTzDc1LDCqW4+zF1PSgbP6v/wN9FXrCeDebQ00ywa9Cs5cuQAMy+3JE46WXiGYEiusUKVrtZT
nb/Uh2fhkmvD7WyO0Htyz5B0B0dpxhKPJMY32EBDMntkxtEQVLEtJHlYe/nrQyBFzo97RhcP8qdv
yHsnbWNx1iwdz2utVeVXHPpta4f71DsykeVI9f9pRcCYCHyStaPRVss99g6L+nbtXdQvcT7aJsn6
GQAMo3VdvUMaCjbOLqujMI1wWnq6h8hsH4heeJLT0knFqsLxq4z4Aw3AlEmbpdY80wb+99SX7rel
ejBVDhXyxQbaki/Griy/ZevAPU82nTumKZvIkq8hxTMXkN7hyLIRhk7ADZqlqN/1skRMNNP3eVbK
WwxIt7c496Rf+w7JQpd5e1eHprl6VuKpGZbLIxFOpeIAOAF7JJqpIF6mhYuXzmNUKSLgNqGk03l0
FwIWXlhWWYVjmXfqMy5mKbMaV9Y9tWVDH54a3Y+7uJapiUCaZKmhE0Sln91EuXWhiHGVNM3R8vmI
kHAtnTFiJVpZVTfUrpqGKTFCxdZosUAHDvoiAwTHknCSFrkdH4APqv6Uk8JgwWO4ubxat7TfnHdr
CuvGJkjLCO+YEJUpMoB6DLq3xtRIDG36KJ3M/cU7Zf+1dTw2wBTEmDVBNux+ObTx3ehE7jr6kfiS
I4ciIuIJ5Q37P4JcBGUExjiWWbyLHs+q4Rt0xhs5B0xysgp96jmexlvfeejWCftJgTfa5HTL7fj9
1L8+Ng1eXQwJmu7osiI4kL6cvGh28QAq0yFyNcW0mKsc4cliMz4A05SnPxHIxAqMsCRzj1S9mCjq
wKDzF9UaaU08KWj3SZzctMZzTgH13+qVGGPJiCKFNiOSqlGzoc/xPWyrdE12j6bUm42raRC6V1U6
SipI1X4+0iZo9g0xKwD6mkzWYJ81ht+3RhnVAQhIaU0gGyybJKo+zZHaxbrWqbFuaUz3T3eEFWcU
SlXuiWlzsJ5jaD6KQ2MvAn1JbKEC4yNp8bQObxeTyOsgfVTuwjIs7d4+WdWBzJ9R6jKTDURKQg5X
/ECfUsDD2lwRDXI3z9G4RoNWqhWufg9sEofvP1g0L6QGlmt627Slrzzto59nzoZBry9cRwkfXeOz
H6bGQPv0A97/9kFxz+qOnop4lc659n9ejLQA7qtxDtQXBrju0hZYrGvKNjkeye2MNvuuOw4F58GT
MmTR9lyzGU8M6HmOBW1/o2Dr0AHeNjTuTu5Kph37G5d65iM1xQgD7/2FBmSfD7YUY15G2qvha5Vh
3NMcLx3ztmvIEkTW+fWHBNRTXD76YJwk4H4DfNpXpiY4xKeu9Jb1RqfXyHdQLBMeVkkYdxXsarSq
C/gaCsDUj1ox97wEnI+AbTeex9BD+TutWQ+SsFiKM9m3QuhZKOjQkX4E0DDEOwdqD5hKNOWKVex8
lxWa7PRi9SJsQfH47R0ikdqUvGzJxXoQ6dr6Oyo8Ru4zVPgAnSmMZ8fbYYris8gBavHFikP1A4eV
tcd/LkfQIcQ9yphGMQZZF5KvaDoK38/q7mgjCQxOlNfhrf/n7Lqz4BSFjs0GmIPDm/UWu4WTLa8Y
r3Ea/N91mg+6sdLfPs1ljQiXmnO6PlvyrEduZKc8oCH0itmuD3IItOVBBeiGlB9H1RLhuIVgEsTj
x8lBD/XuBmPyq4BA36xE3dMFuY3C5TPlWoiEs8RCPW4Cje5+dSfwyv13rg2yUM/A6dhBimdz53R1
euAR+RZAILUCLEiSQThEy/lbrzSoMLLoBeA6+GmG8kOk6lPo26cGH9Ecw/nzFniEU3R0mOIvQ59U
AoykKXbxkZl253THMr7+8lRCZ9q31PkA+VYUR2Ki37sAYE4HBWSWAPaev3D1J6ihI0inoww2bG+d
D9vlbwAgfO7o0FjU4KsmBasqQm8934LLGR+BEHCL8cFYxdT44ZINSWhU81f5ukABxXY7Voji/QQd
tgJuAS7RozViVllkkCY4aHLq3YKYUsiqNwb5eZPb1tH0AXi1OBgvxvTew9F8W7isANIUvgQth3CX
I5rlrHzVkOStgRtgZYNcL1dQBQEf171WvmZmvSJV0ZlqRbZPsCqZAGAksJX3FO8VkfCKaOD/TAmW
ALtSdmKlx2q0I7rxLDrbukLQVr3mMUB6JEX+22EuGfW8I8yc/L1GK+o2mYp6HVdkccUISqmYeJwS
kOok4gtlY/A0EwTKFg3E5pdfnJ8sG28cVDlgu976K9otcT30+9XWST92xQpClYE+tsDunfxQHnkP
+j5jkTWsqHy4rypLxdcN4eIJUFQyTyCPIsGSfWsxmCcXZ3G7Yxyy+fng0I0oeMECJjpQk59OERjy
uvLDFgpFFPMV0zTDZ3JUefB1h9l26SqSE8eZsHaKHOXeZoVw48rdT21Bov+6TXxeujrpFrlQxTPO
jOwaTVfLoH9aGhc2+vfFtMpJ/ImGQ8yqwFw3c8c3kVENO8h4uW+7jB6m3XytleeveIsd9JoONMbd
YHmvv6a5fmyBeE+5LE2woKi3TeN0YYfzvutRQuivOTh0WYXxjkyCnbFXGOXcnmtOMHpYnnzTaq+f
+bBPhC4SVEvox+tRRb9QNt3J6LHc9reuYjmmiI2yC+mV5185ujppu1/CVEDmmOjF04CW9+oyD3LE
zsgZDW6xI/AxHsVqm0GnPn0A1vRj2ikAtsTSKCj1unKWbHpdNVq9+wVUdegZGQj4LlnaqiFiD17m
/lycBcBXS1sgtW85txPnwCycNlfxHRpS/aj7ObCq+YiTKR6xP0kamKAkfn6/MmYuRJ3M0QQtbXp8
0BBM57oJ/+8tvJEWE0NF7YZzFov3GjR7t9+i2IYwVF4tF4+EXWfJItrl4ZbM2h556aGV/dcbxoGG
+HRwfXGDSoml2/8Yode0vCivoDLu6WVMX0WbecE+CjmHyZM9w0gz1rYSZBYia6JjcaplyETQwacG
2sGl2GzzsbT0Ks89+nWLa76fTj7pmsLtKlnxh+CgzGyBR3AJSIIeMpaVgpjEffl7GNmiojEBuSRx
Rf2DN99nlVPOPpVwscQ3JIVqy77psr2tvodh25nVzBhbcJFtrQ/weeESl1wo3DQWwf+YGPQs4xxp
gzLe/MEw6osWSqRyQHpVh4naPOn37iQFw9E4YznwuraNQmfJy1Olr152ZMuWB8gTajoe2ofCXXDQ
wE9v2/+H4fjZRxSwy7tFZ254C5QSzSgjsY5mQIBtWKXCeDNEQ7kKoo2vymQkKYBbncRwdYQ1zJZw
WtXK48HoO5vVFhpdsCSuZ8juidmXQY1XtEIVd1WEgE9mXoZTBMianQHn0UIKa8StH8NzJoMUj0sy
mJZtPrBt+hrRHNu7eIMtwqGMVWsrNRFCRapFGvCBSzEumigAYhghBtJoCeASxWutc1OuLPDpXDY0
AfzZD8XJuOn5WiusKWHICmtMoaP54RrLxyh1D5MkDZfXR92yWzReCYShJSW0xedx4laRK/2F9m+B
bm8M834K9YLgV9xNMmHX97wmHLFi6gIpShzAhcCTn2E32xwxAB29aqSyUhsDlOh5vUAN3eyL6c4c
QKdYu3K3hF0ymnNCWft4v89YJKtR8cUtA7bcpb8QrjETtdJ3CbMr71iX7UoxXCMURnqqajqKySXR
VZUmWsdBYw5Jehr/5yPh+ra/HYHlAqGJuiwHxHVdq60mC4/v+Urc1+MTf3qnXo9BRu8ir42uj0IX
vgwxyBvSxUtZSJpdEL6jX9klswSShpq52tkoyPildjGcYVV44WvWWFQJxXRZD8Um+Y+TUpw1jJ7p
Q5MCSwC4V6398ZhkcGFpuf6TkKRSi5Jak2cKxUeZ/mi56RqbXzW85PlQcE7TaJpRECtN3fFVHKUr
raoCDVw1gAlSrmB5e13MPmnXnIRM3nY87C6s3SR3luy7GcbmyU8CZGZ0uiPuioANZm96LYjGGlYl
Vu+ljMWQA9TSEZCyZYPLGqIyCrWtpTGnmo4ekuf2UPHOV7Ol4V00VNncNSFazHD5X8k7Z4oPDGMD
MBn7apuyiPE7Xf3pRpPa4xrvumMBv8WZWQcce4ih2OM0ItOIqe6VhB2oJuT0+/96g4/UVyG7WPu4
uYOZLkMMqdo/46BcOymrH6DdV8Fe55JRtobfl7qhmEi75iBc8ejn1O0bwQxRxgl64+oWMzYSQarQ
p0fi/jP8FGRUUkslj2bcx9ETfMvogijOEi5xtqDjnAzzs9iEeAf+n1ZgVxnTsz/r3mmKjKACH/9R
RNUpcco2mjTYkQf24nRNUejEUQv0onFxVRzyuj306G5l8/yHN9ihaPbnY3GitWUZa1JIgJHd7+R9
av5TC0Wxcg/zVnZtU5++EVETyxUGfBLDy8MzMN33nz/ohfQzZGr3ddS+TqkNEm4n0/tKKD+V2i05
WgkARLceDwnJXjstLTjTvV/Ee9tYYua8EqG6e5cVtXMzvgSSFAaqKbhQDOPdIVpIWkTUiZrXzhWN
vb/UgIgLJuJ7vjDteeb0kR2skGdM0Lg+CO5r67VB+7H+JOvYojFmbneFH7AL30YhTpvCZLuZA8VF
eiodpJzo+3Tg6/TA545ZU7b+zrLSRUiVLE/lKguBGpLEpumE0b3bRFVfk3zlMey1h5lRGc6VFWzr
w6cj5zqMJf4TELRLgXCqx6HQlYCplA8RqIFct88pXJExCe3VbQ0BSUO0kmp9LM0u1Orw2w2MzbvC
LOnUIRBLaljmFzEJVWY9bSoTr+aZwMwz55ihDmWuH7gph7F5XfugZARa3eleGnJusnj4GBQ/4GdG
c4b9WXvbtpiHRM0pRyPSYN8WbnYqa0sgXWbEk3zv5X8Rhfutjg+qHbeOPSBbJ2NMCJ46aw906AUT
RmLtCNA4vMrXtkyTirlXGi4JY8vDfCSD8t0GFrtbC8pd/UASAaTMlVkgaa8Z4mmsLcyC4wfSI7lM
MFi8VjHF/TDIvuphb2kBK2/oHpoAlzSiUiURrdukSEvf+i2SSULfYKRVfJYu9a/Hfq6aGkClQ+V0
DQGsquLNp+twccNHZiSX00kp1NFz8qlSIdbJDN68ONmx1wSoo3Q/dOtuR5HN/AsDAqp+hfvSu7LN
p+g5jCQSKYc+RsXhhJsZn8jVW+CPUubYHr74zso8tm94YMIRe0GlwUbZYu7/V1bEp2WjMj1blpv1
Emqc+zcO0IkYKUBjlpMAcoHGOWrpGCf5kq2ZETIPetuAp4UC3X4800bqD1goSz+ssIfRD1Einn/P
MJM//zC2kH9uvsFluj02xKok1H4b5saUE2tqu/OLkvaXTLgtAVPycau3nWB1I6Nm53bpoLHiuc5E
5mYMR3thzapbtbB428/4HTFOQPQY/lKf+g6Mf/A1nT6eGLX4FxDEAIUC+C+q6JsL57ZSzpjYD6bl
azaTdFHEloATPLDH8XHor5iDDUuGOWbbtcma44jOjV6dl8WGKDNA8ZEARlq7EZQk3jwr2E9yMrvM
QWUIVo0PRBZz+R//DBfs8SmohOSWGiXyDOYpMYETC6Qw1oHGwPYfWPaNIv85kMtZJyR1hHWEBg3S
H4kubZaB0WBM8fA2lM4yK+7QuyEWs2f0olWj+++yofB+ojPsCf3orCuQ7iRYRo8edf/pXIlpAj5j
rbsdx6/8xnijDCqrgLqqU0tV9UVAwkjfI8cqnbOICY3PA9OYfzgCPH0v4u1SHj9Oz1ZZIoIeQQdY
rt2Im+fy6eBVRcRs53N3nD27YzyMop9B0hv6Uh7tqwOnQDcmnLE1Z11YmvBtBui1C273tC/oXw6B
ZJ2rEtH0ciHP4ZDMQaV6SgMv5pzYBBpfKDxJK/+25L8ctCJYvmtvN0Lr+NaxN6lpNZCND5ZO0kpS
75rYjUOrinWVk+hi0IExm8kfxlXDPEbR3/JYgUDiVYgZaXQ13FuPG2NFxdAUHHrc7X4BdcaxQ3td
q19mGmWsIl4Q7JHWeo2LwCmjF00oTGpi5tgwdRfqzH+PWpSwqd0934W3OZWJeGnhXNXHGiIRy68X
Lf+LfXD/Q9py7E1GQZ1h7rT4y8eTcvbChn3zN60FhjZ2PpX611EyI2URPVywk4C++SnidkdYP8Lq
lh45rzE8NYSH67aT5WG0xLwqg3wO47xW3UjLp5e8fUuz5tuEH7olGRQvxtSDLa5wBmhHU8KIA7Qd
ictBdiuCiQNIz5dnBW3Da6WPZu0wStZt0MDM7Mx6J5GS6SDZUJ199mUe/5Bibv5cikaT162/0Kc+
Y9WEV25+3nvk/uODQty6+hxujWdLko+0xDXTHj74I2wgB6ix5XzpXUPAQbhbR/bA5JLKsFFtFGEN
59jePqU5tI4iEdVrh0R7+LsG/KrD9SO+cJ9pCt0aC9aGgTxLT+QO4JLGsmSXPvc9bfGiieFet6G4
J1NjiulwzbCPwJb5NLpI0TgQ6tJWLtp8dV/ka1IaS4t8twonNLqGdPivy+Yg+RMYm6pHwUTgKIiq
7yV8DFjFfL74z18/vq20ElHDLyMMdvo7P0CqHCE61pm/2OEVjXxBMO4Z7gs0atzG4FwjhMHioloi
ByFGOmHIoq29QvHSKf2rvcWthf4OP1ZoWIXUEFhNzFlTUpVC4TSBMmV2xsbR+At64VXIbCYRQ1LP
1J4xdHdi64xJENyVH+RD2CRo7nlUJNM7KSkqt2ryOsaQCCREW6M82NXRRWyjAduTeYq5bkTW7NAc
8tPfZ9tEej6UCRccsf0+cGLDYZZ0vW9xKZ2Pd+hsMqeGNvmQL5Oi37hq+j4WmjNNWcA3m9731u8Y
M0hCxRU/PWBDLG8XKpbx6Ph1MaGsPkNHtBOfRuTsYLlZ0lwgmV5O+WknZNJHNPc79Cfj0QyWUbdX
RGic1/cfChdDU9MqLpl/JCiVcFnn4sKhxIy5FUk1AwS/H38Mkxwq0tAnhCbvBHL/6EqQGecgtIkZ
QsO/HxKtkHoQe/YBsbDDmfBXIJbIf+3xISJJkuB8aUz1ngvqTmsW2FOVyTTdZ5YK11xNw9EyzeWN
IN6ruehasM0/dJZwLvISR7N52mlOL/4pianZzKSKQ5xcleH6mVGm4xbme3DZCQH7Uxqw2xvXZJjA
rPxGi4ImrA5E7qG0Q6Fb3wTIstlfMknK7/FrKpyZ+tKGUfzPNTzy7bcLCH+N9OFO78Rl0vd1RvFu
CQ2WV99dY0YOn0IS0o8okbGxs/x8t8dyO7o78k5Qr9bNZj23OR7tdReCBg83tYCUOXN4u36jrvr7
U0z5aAeBLM6oyUlASbHbWcEm5crlHBq41dSsmAwJ5rkkspvOlOPZ7CR5b6hXZAYT/Gv7E/48jR8c
dqiA9VG+TgBV82vHmQux51vgBOOr2IfJ5tfOondr3HQG1Pl03ynI3AN5KVsN3cTvuHQ05ZTClx4m
JVwsTNVZbStymNOIKrmZ48Qzyb0meV3RQ1YGPG/XH/Plxvss0gVD2A20byDopfPvqa5CdqZGwfPp
MUOfuvO/8+54z8ndafkEcnXUp0t2ul3YQfFQ31JUKqNGbMeEo7VLK1zPnHnK0QLv3LMmn/ygbllo
KdS2ttk4TU6vJXNBN+NdWOgByx0Up3cxae44ziRgtdCn7t1LY801JwinNRFDvaNEkQC9mOz8UDHi
c0SfJwg5mhCvLNG6JACXgVSQvKifetWUrfjGJDwaqpauHSwXJKCt19LF81ALwAAky8cj/N2aHUvZ
aPHNyEHwAsnMOLgom5JXUV86WmvxHvm1zqjj+YI8EdEHc1RA/SK6L71Jm6RBMIRdQT9CZfl7WzlQ
g26FiMOq7U5N6RbNlMdsp/WttindHzD2ResVT8X5xm81ddJPgj2o7H+gcydahVPATWifxO5JHRez
92ni4kGuCwsWiT7I4QZtaiKUgZ9rbBCv77kJYl9cuJtExdZmdDdjnAN81KlEiN61N8UOsTM4wolx
1taqtcI+JSwHBJtzMdqniy93x/Pi5qlNZK/udb/ZG18N8x1V2Um3YGPHedkn3f/h25UVoCKkiyZU
Jvj92g5rh7zNiLuX3dsvt4//irGJk8wr4XucY3qnaYgtY/12kNC5E3CwwbI9pppfZ6z8LCV5j5Ru
LRDdMkVhsAh4iuGike3RLR2tC0cQ+y97PUC+8Gx7z2fDCvLkSfihToBXvz5PpmMfAa24cPUWN0Dt
4orhfJbJU8YlXO+JUOrNJMHgDnsPqOJdrjC68zI3N4iPGXkOFwbar6vfPZtDtMSzulPncJZ3CztG
ksZqUBzmQXYP5a4iJriWyRlHwd2EiRwPjk2iOs0dH+g3dgr8Pwnc57tnWDysc35s6oSgYbCaOGhJ
3J2NtpQE4Ff+0awRpafw8Ts9iCSb+MJwB80fqmbf9wBicAwyabITauQ0IecJH5v1tyhzym+oFJ0Y
W3jYXF2uLmA68LHLRpptpLvYXPZxWw9v/d+FsQzTGUCAK9O4tdOzP8EjhoEi9S4g/LgtcyN/yF8p
Hase2Ihgo4ZSDO5XAKoAJl5VwQyaydjtKa8rfRe3Wr7QQ1yJK5ecEL7ITSw9RpJgJEPMKw0rs9XD
jabNa4DOlEgbwmKD5Wun3rnFY0BXSRSo2P7IPquG40aBEwWKDv1sQiybTwMGKHWuvp1HNHDyGNTx
iciQa2V/9UDeKeG8uUj3qjdv3CIqykfAvVEyo0vvS/kRxbI39OScuJQOHNsArlykjSsTVjaIqpXw
RKyvfIsHWCNe246NBJevWFgTM8M/KoA+S+e7kztjRfCthqvBZipo87Qif9qQHGsTOEA9wWOA0Py/
boMhSaGQYPWRcybfHjJf7UqAevgVsvjRhBxziZojRW4/jDlTjVxxJTOCzpE2LK5ZTy867FWlxVYX
ye6T3NWAnNxjoHBbInGDKD87Nr8PR5Y3IQ+yMCPEQNJsCHP45xWs/xiwRwNjIX9XrRw710RXs2OE
pTe2a6BfI7fCOB19ZWLS0W8B8mjkHn6/EX5ztvzSPTT4Yt5ozmqd5is6YWdRjGz0vNydypadoGU2
Oq0+XLGNIDIwyGNl+82Y70LHbtMTe3xSi24k9ZAwRtWcRhySGYg7mriFPW/ySwYjqPuMcbhe7D+9
W4GGio0D4s3wYBQwAYz1IneiSMYHCxUxHAu0Xy07oHm3mOtD3k5FImABUVPz/y71y0ntUxSYuNzq
bn6eWkzB/X0/pwz8O9yFKmyPZ38kvNgGJ1LSQBwgskanHa1bCbbjpVqlOrZ6r5q3Z8EdDmznkQeQ
CAeGdhhdqVUL54o2SJPs/esL9FxWC0yB4St1xct16bW7ZYC07W8C5okmiBbSGgfQAntp1gPkOA61
KUvKIjcbgX0NhjGNY+qg9vZAf9uP3UqDVGtPEhqWh0beETFdSIdsepFN6yvCZyU5sNZFnn7Xh9iG
IadgTXxS7nc84lWx6WNrLtFtwhmjntmUdKIo38/ZmefowUWwUFWmemTUOgxpbkHRu9ic7pSQXyXH
Gp7HRHf1ruBMwc/qVd19M1fOWp0KGbiEnRxp/ppS9Wi5axj6XJ1mvUrxglpxojGhFvC5iv1qLslY
cJKFUIIyJxm4/KAyL1XJOAuQ43LCaWLTBHbPTIGVaO5lhqjwPBt9e+z0ZPfp/KzFt6zbIG7Jhiep
Vt7DhgrFS9GD9vWZ8+Uns00LEr0sbp03v+Ervvjip0tr0Pf1SEcvwdfy+K2BRe4UbSs1Gf2FZ4xl
iIrl1tvxx+MElOmVofOeuIeNUW/H70F8LzgPbL0bvMH1Z39/ckdPEnN1U3GAFePMekwlo+YaNN2y
e8CyoejD+JPoMCt+UozthquwFXZVziDUpfGD6jOVmHXwsvfKzcHvL3UeqCzGgzW+oizrJ4dQdbgB
YKl99P/50oRKny+AAX9VsItspUJKXqcC2zG+qjPWdCd4WbXPikFrV9zP7nDUN0d7/SdTLcDc27qw
42/oMLzjMqEiVB3k/8FFAd6F9yJ1MN/42BKQuXXF0oZ9U8RQHhC5HaOnnBXgjecRPcDIOx1N4EDL
WoVuziQT83cmLme+09XOu1tICNgmuDJXFVPedTBjl999cpcfn8xGHL5T3ZJEKrqG9ZdDQOSUfeOI
MWsyKqowI/R6p1BaIo9jKtPNGL7JAV8dRtB/PTAF4k/z6/xr0cQDNaksniVSWkA89z+vFNTDtJDl
Yd/lsPb+gG0XK8jdL3iH6XjBmlohBAwCtYDr5s7UUuLuP0r1AWAMnIiNgQGfGux4YN3zg73YGrg3
egSVoMej51/Hk3rodDhRCheu7LFds/HZdZyhdDSQMRu/Cgl+pH4FoRrxBZ+WxCEcc6KNeqMCoydg
SE/mDTLw1q3IzE1mpH7yzBJZiHR402VCYC6BM6Is8Zh1HrRWDt0cW3yzopQqawkvJkvQ9R1F21eL
nZzQxwUVTag25UJ781WTSTJX47N02CLQTUt31yLNQUETvno0STfuE4kZvVf9r878H3zgD/M8KMqf
W5A9oLiB5+wB1T20Vonm9DyPM7ihCeDv70BIqx/wpGktUhrJpLdjgyDjPPjNnXRKtmDmSzwHkfd2
xeT9gbB4+73K5v9OHUDzJr4OEwO9s20vjutAKOZNAKA2L28BrmHPTcJ2+5rDOS1TvxZznvUntmfM
F3c11viKSjfdJHgfvsZY2j9X+oboCjdG9OAYq0F/S+eO+/T2ZLMO7/HL281f/b3Uyllp4qH5XYNx
AuiT30Qj7V/HyDd2+Wnf6mXZ7JJ/kbir0e9WAFv7+Vp9Nr605sIcEUfqiSJufMyoziQvoczqwiQw
tyhkimtcv0laxsd7sqs3cZJw5KEB5y6WU5C6s5O+z2nv7GDg1PIm5GY2LZ+KrNNLcgdcznBArM5f
kXNMhJ5DGd9Luqq1TEXlvQLGZ3Oc9qTKZwzzb9StLJzRfhBF3mgnvHkTQ47YpI0krnyS93oXYCfB
Wr4fJHba+9WbEq1E+Y9pTnsdUDjqXSRAmU3hijmf+2GAEl+dLk4X7eiPeiAPPZ9pR4VFy4SDPuNL
jLlKQ8Z3TXEwJzrd2BqODGdhI28iMzI08I0rWq6OMbgeMq8D+tDMLsEPDbLTcNusT+dufCFrDBrS
dIiPg104TKb1E3+4cCudcioT67mDIxGE7UkSkDn06c4tRk45abSzVPpvsqClO6bn+EugnB3e7mm6
LYJ4c8ARouQQ9ysVEd7i5wnvAU+U9v///DSAh+IOY2YbPMWYplkDUpIAfKjw9O5o9sJoDAdwUyrw
dRm2HeLESokj7P5viXEy20+BpQ3C+8qa9pYEOwErVgja2z0yCTpLMSOO39gyYYUPn43wYFx31Vmy
oj4JUr/z1k3BNaiMnwc6e9MC0naQE4MhTMpyGvqXkU7aC2n7Q8IPrfiss18QIibywONCDj90JEAb
k3+ChSygCUoJOEK66VLxf1eBO1zW7NGL1DsVNSWlexwTVy0K2uR4QdtFC8+yKfUJrQCg4yMi6Hs8
HAW4WQmSy6UPbFjysyDzhG/EnkB28w8NuaDRX8XUAF2eA09Hp5xnNzwmU+ILFow+0jZcP/zkmAk3
o0tS9Av/TzBMmlpR5dYs22t9oGfwn/A5Xb3hW4V/jmbkPjMgWYL+FbfLyaywqj9BevtYR3Ie85qw
IZLzYYXtUGWo0i4tlWCY3Ccku7cbm5D0CTFIM/yCDiDhhyxY5iiRTI27bU3VlUjcjfbvfpyZxWtK
wbYcc8DJ8wuB559R7zvFMVRE7uAd/dg5pE09GIHuiiBBOT9nIIzfxNk0BzW2YmkBAB6ALYRAUplu
nVnUXkbe0e05qFOSZSunKBz8juc13iZ7lcnug7BpQXzHvtTyESQynaXcrT/iN8TtJK9UnhiUxwAM
ZfaNOjSWkI8O9WvjU6kBwSPEHmo4E0ofMmNqvDKejby/MjNw+oPQfodSL91u1mEjAcof3DtkFKeq
PHNgFxKQY50mcTrlk7sAqhTF97TtKyahoF28pkDWZvG8LdAKtr4cSqcZTELGxJXdCvoL7BuFDy0i
7mIb1c/Lgr4hDYWvVtyHCf0Lbnf0XIInP7YGhyUq7sktYL9ri3OmyiCHuVl2fQqTSv5QAX/7PgsH
+D5KBhNW3HGr3tLUnVjPtXK4WCQ+9GkoG4V/YMLNzBL5hMKbuJlqggxkwlf2OaC54ZazNH5Wm7ta
VuJdG8DiKRDdAlG+J4lTDqqSrMzScMfPaBtm8roqOr6Oqg2WEbH/iL9tBlaZR9BGFaDz228kdLhv
WQo6dURI2NJOD++Xs/XntNrB/X3kgDzNTq3Pcz99yl4G5WSVhZtHA5Cs4CbvkZZUVJFaF2xPHMjU
jcIAS9V+snFxp/gMi5V9kU9nPiyb1F6iCDp3BN4LSozgXoS+dZuReRgi36JAc59Eb+9cscRMq85H
2bkXkUWGz1OQk6s5BzJBIUhqfi6e2VmIlMo9QChVBlFKo/feYYha/JHMAgEEnGbzBxa5RFAEYuMa
p4S9TSWhRRl6s5bEpykMqMuv+sZjKQEtRRP7bkGQ+XSXIY8BgKv1wYOyhTlyBt/wpReT/nqBdTHs
9Ep+etCQatI3iB0GUJlzYWZtYxPGQGqgaIJaTOaj5fqzrC4CgpvSIsxjltG1646BM2mMBxetlG0r
Y6IV817TvFo8nOnDe+h1FVWAnPSm39A8UWZUtuypcLeRwfNgtCWEWe3FE0Ql22WHQwEeRNx7uso4
1EE14hGls7zVrltnKapfEOggDocRs9CAj0rPXQyvtpICV11REj+qRKNV2zFOXT0Ig5NGz6Bm9SnV
j3egAcGH8PsDX9nFTn48ic8ztzszuiPUe/bPP0qfPJQfWBbqnWgE69UMh6kJCWf0BgombVlmeyAB
HFEXXJT27l6T3ubzfx6WbtxPjgcQ27vw0RlUuCZUViFnaOfvJWdwYM5YbpEjeumurTl4WcQWrs9j
A/28L1R138hHlPI8dF9hB6ByqugjwfxEDzrszaSV7YuWJUI3W6KpKMk0ltFwaePkJnCAtCGEibiw
9MGMUVOAuz5Dqg+sjG685UvUhSL/Am/zGsgWWcN9uYsLdka16zFlcodjAyJDX47aX4mGtBEH0NGx
utacs5B7aDsnxna76XpXdm5lSvLSjwlPDijuO48XbKG2QVNO6Qs9+7/9GSU0iksMQO4BAchBUTXw
pYwj+8Kk/+ayaV/o/X0TsPg2M8yokWuhm44tCNPvWoaJPP20AluRnstLOLr87vZPMo5ohFiYSOAi
dzwiZH41wXqtSdYB9KM38L8/Q/mgImOXcstnSof5i+3PCEWyk2lgp7FApcmtD4e1qf71Z8gYEUbS
ZTeq5fDEQaGNX1huOn1zOSgVATSvFdHgsFar8hxoUmRSHz0aFEzy5chezUtv3DTX+jzVHwISWnqo
Qin/1OD+/IW3/5gA1Vl9Ya25p+iEPDcTvgX0omZVOTvi5RUCupRDkCXTQ+Sg3ambLAwOJPFQ+6t9
GQh/4mUUbprn9O+337WC6Fi8JpX2rdGop15T6MKB0wkFkQsd0DrtRXxVwC2ngYa9mgOoG+/goFf5
TjpEpVXR0hBj28lu7TXjQ0zGNZLFbbP9pO/Y+2yxM56fLfAl3cNtJ1u1uepVqeiio8k+ktr8l+WS
q1rLB22+9PFEOEbyIhfNViolLN5hIm9TdWhebtV4q097LfDy+aS2wOUTuX5esE9fJJ1T9skY1QX3
Mtl2kCRoKwt9T1EYdEgqfkFzUJsVtMAvivXPLPlVvuM6qvqT15XLsMpwt04wGC3ZxmIddfJ2deeO
S2LACB0ivGUhs34R0yCx6qkIfCe5dFnICnl7FCcuLQitj2YZP+9oWmfd2lCplDXbHkq+nJDsE82I
s9Td8UjiGNaLBG29pDf+MDGuOCwExyJ5TqGbKcFzaRliiNyICcTJllR+y385xWMwB1+LKMkqK7Yf
Vu/dTArqX3KT9ogHs9PeMJXnQow5BUi/H76+wFOYKXPgruDpzjx+Pf5/sCjEYc3a+IGRCto1CFZY
9LqqJorAJumSLpBxDjsx6c5a1AX8zqcIw2BH0BBRcfGwgLRZKiHP8MXCfm4kVJcQkZ7eWPeBlqAz
TdJVDb9rp4PEuU1yKqN5s1e9OFWBkPobjANhUAFahjW0ctg78Rz7cXxwvnz1BaTkDdH4CzwaBnDk
6p8R9sXKXhERIK34Op5ko/WKP9V2uHyfq2EJwNXXpwAO6oe5PW4jTjr+adZjxknqAbs9IK4NO5+h
ZQ0ZJl6P/opUwKwmF4wLj1B+NFB8FMx6uPjZiT6nheeLCJA9pjs5EbPGjXIYjqIvh85ugHYuozLc
8vsLFNef2nMV6LhOX3HIuwUo62tFBXCctXTlvmdsAB5OWZEGXwW2VaYfNuR/rfDZ1SAh/BhKGI8b
dCpwT24VEYM0EZ7CoIPQ5fJItcLroRtWqTWL6RNfg5h42ewbFRRoMNIvzdbJFDFiqlnvYxOS6fey
dl566ZOhw8e0o/eiiqP6qW0oAMS26g4rZGVahB4O1dZ2OIdkIvk2flRQWugojVMUMzYcYVzk3fMq
Q/JibjcFloNQLJ7ncvqNH2oiz8Cg4FJbbCT8mp7Qq5XkX+Uuf6s1jDXWuiamgY4KW/znZVvNw2T+
03ZijAr2i4+1Mr+TXviHRdeXSQmfWxjyAm2kze7FnRNbORKoGg/C6rLDnSkwUkW9h/1q93sq9WT/
v62dL1fib6HNd8GlVTp1cUJgGbwOlJY6uHC+nSyvVnXYDsF6dqIj/kBRH3MeufF/QQ4e3nqLvdzb
IP33jrmeFOE+gFNvxKJqm+QhbfY6sLsXlWpGcTURUpmkNHrQS6jo+MSTqbBLQ3t/7soT5yIUlAvX
7edCJaYFln4jFZTK8whXLVDBLUp9cYxAxaZ35Z4KmCPT0nNVIsaMbJ6hD/M0YqEQBwp7OmtdlpSR
yTWxfDy41/2Cb9hQvaHbHaDFz50yU+JiGDcWHPdeMh31w7BqazEUTLP2H6lBVK/dvT5W87pzUsiq
X2qsYlSmvXiA5vCvk/Ss9PCNFWiJW1MopIxGBwIhQ2RF4tDj7KeQCGE8SV1Y0HalV0uGTRZHEnMk
oyjEEtP9ekVafx7LK4/b4l2/MrVys+RKu2MuV1wprF2aFOHZfubkQyURIwTM+2v+qbCvzltWdrT2
VNz1lsCFrvV0QBaz1sTehko3nTR7FovQDSM9HfKXnuv3iui/xJP8Wj1ZBtKzrNeJdKdyygrTAnKO
3gM5JzjXcNdujz0OSqXQhwsUpC1p6kXd+JPVlEZW1PeK3TIH2fLx6XMqVL7REs37FCpHzUoUu2/P
cpHHzSKfwG8+Ottot8HVLqP7os1wDy4/gfslHSoA4fpfbLXF4kBbBwWs180MlYsOz3k78DPppXL9
fVX/iRU+dZFRamHUq4zzdCrWM/2aSB0ueCdqdadUuBAuDdi+uEAq+lowrs8awwe7khhyK7xgjoMT
rK2VLzXVxdnBW/og5/djDE7FchrRCopO3ZhcpoBzP/gRxamFnnU4RxJbzFZv9V5yY/W142Ou5HZI
gnOH5p5b8alwjIiJNYwMw37In0WGquI6sEYJr5evoDCFnsGxYzcl51ho+jc504NEbdhNCgEskLDN
KjTCceyuxFrzcyREWPZBZrNE/SvZKOcIdVXadYO7rfdzIArJWCwAFqmrKGngNG5Aqymbfvn65xZW
Sv0Kes5k+VWKS2a3oFXmFseNTKIH+oMbJHpa08Odg8YXR8ENXjASiy/dkkkPN8O89vwq1ZMVoqqN
zoyihQZJCvZEJoTQC/ialbOA1vQZhH/Y1spiKoDf+2Zfl0HQNgwgnbug5XUmhY/MrTpZFoJ4d8M2
VQMvsa5Z5n6MMrCMZJQgcHhEThmWItGlH052FaRFp7sScW2F1DNoC43mJK050iCOX/JnpqCfrKYO
GC8lCEiySuLic/o3/HNATwoEupomyj5Pz+ECB33opg5f/8V8vba5F+7LnARnzatG9INRftqGGUy/
7qwp4nh83jBnYo4CCSbgFXkQYqhfSENeRWlbhr4oJFUOrIJ/2HihPh55VAuYjT6j3KTyBG6tsxIB
D/6gb53WrysI+NDhws6MsZTl+kLMChTTxsdhuhw+5L5xN5xdfbGy96mekjDFl2Qmk83uRaXpxTEM
cHPBs1EYB7ZjozIXw0z9JYt8pyRyZBDbiPanObPiGuiT7t+kQuPbhS237mh17xB1b9KDfGdvQUX1
PsVoKjFODETTEVRm0qpxy/W91zT98z3kIa3yefT4svdCFtXV414NbHa3VMkMA/1EiiWZIlvjlcwn
7Gph0zNvcIlaHldamFklVxWzeVuvX4fxN/R91bwuAMO1+sxt1QFJgg4MqdgyhxxTfuTLIdB9veeu
NbSZCz2o0jSaPsvclYtD3QjASxNPCJCFYtx9dcot/b0pP+F3p6pmfSj/j7wvv3GZoGNrYyx4ZBx3
omkx2aaY8v+a1WhAcys2ZBb+y+Mu07j7ENyh7xGA1dUSrWGBv+O4qYiffykaRFht/7bKzyLoKSo1
rZFKdqbn+2tutDMTYzNWlnHjFUKEpwPshL041kLzx7nqGNUfd+N4SLoVAhtcZtAS3XaRulWpNj8Z
VdyFFs3hwz/fj6mrX5b7fMQBfYX+TQoI0nMyGH9Z29y0cX//YdbkC5sBmWfA3vfOi61ngMmktmZu
20boNtRjCLP2X8jU6FbJgIezoKSrCuAXGG03RcjUKGHg/GT+foSk/E4iENOEz8r+3jKhwVX7anTN
JFO6uHBbbhgv70+U3a058vrMfJmQO3ou8zTADIBpc4lJIdajd2f6lqgSS0zkTcx/GShMUaECx3Ld
SEhcNGAnffLmLTxvKQwfXb1VDJHlL3l0ZR9S4T6d+iZ6t2qsbgHIDBp9if0cyDajd3jqUUQgRC0V
Gb7jfE3lYaszHxOyBb9BmVfZNeCqPy8X438Kg0RRQFs27C4m9GNEP7pOLxKa6bDpY7WgPl8kV3uW
0kyKy6N36QqLIUlFw5ZrEh0oknieBPYZMWpKfGqt2TEGcmZJZNmvNhmosekd30eezlw/ie8r3mCr
NPkrhehfPk/DUyYz4CecKgSJAAMtOS/nvancOH8Bq/Dezm4dJEJn66goJW1IIPymUHSkdZMB0i9Y
WLGwtJwkKL59KARs18mgJkBpwZFXMF94F9OsknYJXHN0NPg+b7j/RoXzjWECJiP1bkCpa9Hgrb9t
xXUbZ1cdWqz0dtGpzpkGM+2axwMzs8SVw/Gqqs+l2UnyuLCdUVZNujIIpeYI1MT+UeoxVKnKsKw9
p9l53sQen/DESIV0hltNBmYxatNqCGeSgJGyBKkoHuEzCzKYuxatwoZraynlxogGbBF/STktFFGN
4jIolRW1MXk4ipN6r+HgOhX9cEDZ3h1TdGWNIRyWdvVwi2Fc+9qqkWR5Wos+xWfvcd5BaLVORyyy
/1u2bEEhmpyp33Ww3dsoP4pToUAA54IpCdvwXQhlJULrZts1Ko+nn4+xTI/aDpjwIXeiKTcA4tSX
751odzHPP0cBM26RVQIBB3qqy8XT11xA8zdrEthI7zctLeH63Z80rtoQ5qbWiHC6xaM0ybtgZZux
jH88qnlvlhj8/R2HwHy8IJXdrFN5skvpVS/t4EiPGDgeLRpy6OxsCykLgbQUWc18rwJgcpZTuiWg
K6vgL+YxTwgRRrG68p4kevNBAjqzmMtitQuVOWEHxLfT+nlhrOu0ND6jugbSIxuOFlb4gE3oRLwW
VqM+2SQbdRUlFDKpc46gQ4HAfXjwDV9+oH8nzzaH/R2Qg8MSAFij/k77DNY7k2VYYbCZ0KGLxa65
VDzXZ5SNEEWw+zhFmNM0DP9eBl5fUI3QgXXVdDahvysbtkURDXjINIF899ojUpJ2Rh5GL72fSXhu
fSWuFEMyZ61NvLtncIGVrqS2f15RZlEwrR9vV5+DfwI5hkX0HRMqtGgNPsR/AMdh+eGOdsoWT64F
Zf/wcY4cECSyNjm7+EjoTzvPO4p+2oqjb4yOOUF5Vc0OUHg2Nwpf0c/SZfvmRsG7bMHs4Q3xQtR7
Jzr41OLLZdHyhacxCQOPSGPEpPgpopnA1Et6qXrDLLZqW3+r4gbj6rH1VPNi3GX+ajdSUz6HvCUw
p7vtTmG7PQItX+1iOQV9ti2LQn1P1vusiln/xeiJ1ZHoxmCI/IndR2ZwilwPFmV1l3+tdC6BZ+RH
Htuclt8O39us1didC9xg59/hWc7AQc5Ac28z7kkvsTTiD5cqZESn2cg3TV3v6XhcieghBoSMt5a+
s6CPSLi+ZrcKT7Zbv+0A5Jsq57ixNbdugq3TE8O7UJZXfyVK0sfwYJYRJeSRbohp0OQ2ePAQPALM
JX9LT7abUyKnBkdbsLuL5WbMBqiRRSQSHojQLDHI8ZCSIzkF9ubSEHKhR5GQWpQKamTJioOJEO9a
P6xVSCfiZiwh0jypzviQFCDzL890/OPBjTBu/tfAeSJIMuSAHvkmP+FXJ2d0vFRj6zfPg8bqqxLG
JbVzM2DMWYU5CNIcrhdBmcRi40nwLYIP0IHgUitSmdZAd9kf4Eq3G/vBpSyupLq+zMF/TrUK44Cy
EnWqhb5kWp3fdZOriWuLahO8zlJvOc12YSuY4OjSaHlUWGz9ya+n4XX2rZwu4hA5PGzCyWp0ZTQ4
LtpF543xU8OLPp4lkOebzAcdQE487QQR6bn6ljgiP+jwizZjPdWleZnLkTywl4C4tvsS5t1wVEF9
zYeUeR+5ctoV5iganaEy9JdmNmwIqzAJOUJUDJ1tHWZzI/i3D3u7MFJjq62zMMtIGXJd67d5j+kE
JJpZtG5VOX/bnSgpGc4n+gs9y2Y4F4P6KOJM1tDlS2q3WlMk7CKOFK4qxD5lFXpCobIvJFU1TWoA
OhgJ6zH/6LDqTvEEH96WAruObMOHVTbHU1A3Jy2LnV98CJld3PotC3a7VY8iozmodeDwdfh+FE9N
hBO25+Jqfua1ITErDA8W9b5LmY65qRL+4vz0iNhF12kTbBv0O7kciBzXK2QGZIwvSENEX5WZTU51
jvuJ3g/W3vnCcvDha7aix9aXKaxDzdlQq3rJ5hyHKYnOu8+YgGcwik10x2qgsixA9t5nCP1bJhGq
FEIYDCQx5r8OKF4InUk1WssLKN2NrhAErdy/8VtwU3oG3nx+1z30BJJYIr1ynhjck604WIwwsMzc
cStqCnXfxWOfT2a9Xn3BmRSxDFlSMd1bXbh1jxa6Z8OThH+7Ew3/gq2xunf+I0/A2v8nF0I1mH+M
/gbuY0nq4A6F6dvSnAwGZ1+FENR23pMStMx8XEdy6QkVORlgMVF8E1ZUfV9W7tRKF+kF863LQ+M1
5nS8EvYFc7zYZ6lqCqWtD54yJ3iNM1lepMtRoEM2r6iB4sWY7+SGAhSyreBxwr5wJT9rAGzjb6va
pfwrUpqI6ch74esAAKnXMdRfBXFIN4Nfy5jDmFJosZVT6KINALTDtEJyLLaU4YTjOF/QDfXWjQ1D
Fz+par3EmhRdaFn4DYMtVGSTBLKYIT6Pht7E0u+HKU7u9TeI+D8E41Nt8xZ0vq0Rw/hyIB0wNakS
WX7U7riXI7sTQx1J4PiIzvlw3sBL2FKrs3Mp//Y2Cpm9ZFgYxjqEGHSWqiIO8yH44py3ITc7LLxt
KFmVxPvy+FkEOvRjaueSxUJSJtPurBS+oxl+gCkSaJtzMxHknhcgqBf1WbJOVjNjm95DoWdb0p1N
Wesrs0D2aqc/0u/w3fGv9JF4w15B+bt2/e157GNS1SE0viQzVPQk4RMnVAmgDA3ZqH8NzqgVCg+8
OeIyvbW9EAy0yflbBfZVbVaWdRCaXz4aArCJrxy77W2Yh8gBoHXOV4PFm0hVnEpuJiXCgnd9vhRy
ykRKngMCXCTsIluFitliDeulYDKOBvVU2qXI0cBZHrN8I+ndiZkpVaY/F4x29+e5dPg9FsBCsYGs
VA1f0B0tc0atDmq0nSprC0FsBN+y3ljdf3VQr8MqG+TdtQk/sH0yOfb3/aF6hZnCfs7nUhKe1+sm
EtgCEzdv/tzv3IaGb2bWHE0W3p4nYrCILGlaepJ96/LlzzXXC8nl0PPvBcCmoT7QHTe4ap3rq4PS
Qgm1X5p0ak8t6wXvnwWFQd2ePeWpfU0a7i7kkNc6m1j2LKWLqz4thWAog+iqwyhEuKzDgM426u+B
plHJsF2v4nM7D7cvkgJq0HgVZQCbIW0j9ZKRXkfbpQT7F0Xe/jWOKs6RiEURbBAfEtylKWS1XM2m
ShgTMFHT3kc0CKUg3ZLpD2NFV1ejjDrJVlu1aYGz54l0FDCNXhH1q5wzDx8ks2yMjz8cepQwEkhI
smOknk1WY6xqc/bt5Q3oAtqfC9LyPZcOxdo3AfK0YT+i3F9PWuEI+kNH46PqCQ+R8YqfF0bUZK0k
VJK2z1fHsGuZ9n/9sTHYVIUgU5yCFw6wZAWrsNQuVy4OpekP20uX+Bh4puXHa5ujKQOltbpZ9V93
DoPzr3gJwy+N3TWG+SOlimZ+kLhjersupN80xrA3cLUgP22lH6on4vkbXSoKcPy5aS41oU6iHvAh
8tY3niI3MydOZS9jntgh6kV6KUVlMbk7JFkTPkWKexItLD5sv9VWlnYvV05BOvvDeOWEbbT819O2
1d5DGfD6OywBvBZR3xYhx+8KGF6PNmpBvFNILsX7cbbTYxstDSlsGh0hq7bvzlXBV029168mSZRA
Y2N+0GfwS7Zregqz6D+Q8F0/8ra7A0BMWRG1wKQGe/WDquL/UyWWIlzoIPDQjV9BD8LPOh7pgUY3
Di4ReC+GZ4FS6pOlCHlagoK60f4JjZu0XlzLAnBvLd53RKIIBtYQw6UtxO7cT0zfeEBKS60Wpa/p
AByVl4mbANR+y2dNIjVB8NQcxFLla8Qc/U7Zgk5O9AXYXyYC+gU9BvhUi51uYyOxPAi6uLzGJXlm
3dyD9CyyVJZGNAjAEMNeTtpvURDxNk84HOfm7iguGOLQmxI5UQ2g6dcVy5hSLmWggBPQKwOj96xD
1dgXb9t7PtRNWU0MDcOuPh5mBdpqmOj1hip+ZccI4VMi1eUYtWidtaNmt9zqvmXVQQZP6BLpO1Ik
vMPCJSSdAixp+bbjvk/AF4VwZa46+9BrULuuu5PA4sf7qu5DBM+anLmxK7iDjs33nXGrZvqGKasO
9XoHiK6ea75QzcRSofMZrMqCqoFOxp81wP5ddcQqR11aS8E4GqR3EbLT4PrBNUm89Gwbsif+vJ3z
PrLPz8CSpLFgxE5xpYHVxA/PmDppHFho7/8L3r4dk4WcIpngrk/8oZrt2u6rRgKQQ+zvE+piidLj
BhcQ3MhzcEm46K5hCnEX5K4XMxZr+9CzoawUiwUmyU9cLiSdgy2h7TBD/rMP95tXMJiB+wyORPUR
O2HBYhXPezAszRnP9JaZZZ9moUODwVSbI43wqhHDI2bQOyhszBFzji5XgYFOIhwyj3XU+yzSpXma
GvRhHylhvehEiMTQZaxytNHmmItjRnCIy3K0xH8HupnvkFVNXNBxEPyQtynG7wISJEnHe/BPeAfN
aRK+lkU4FZYQDNR6kQo4RomOGtM+c77otftqnwm2HTrbsq2lhneJmbDfZoEjoDvik7meaFuqCVl2
c1d4J7IvO+J/ENCRldraIjlQI8esyKq6aguB39Zf6C6rNhS8JOnnGNYt5dcq3C0UquFRjJaI3PGZ
H1f/9nH68EFZscszj5lgtAH3oz+N3nttlGts0dcfzQSQ2nNzO+9x0fI8lmyV6NqGts7i3PM7Uwlc
19qPBFYc/bTXbo9tyJJZMe+3raUHAMsew8nSE3EEcPE+xiks/Lwt0Co18EPGhFJhblDfYfyVviCE
ObU8L7i4GTEGMnJAD98FDwyzdnCbwkviMqJlMKVW14eSJggnc9gXJ03UC+VPWxvLdKOUMC+sOn2M
AV+aPMeW7kHLu9deOTBxyssIL6YljoiWc4q2s/FKUuD66n+9B1hG4lugIh31uPxVXrQaCJ+rl54G
UgwXuwG/RvHa1fHa8l2FJkdEkSdftqWaV+jY0+2xrV1IiZO2yZhq0QDGb4Q22IB2CfniqHK+H+1+
xMOq3y/cAaUwPbYjIaaFo/WPx1FiEljAEFxI1W/nHtyvfuPlDm+wXNOMinRBdxlxsuuQZEa9s9S5
pzbPF/72WnhU1pyxVgJLftLHxjjHTRZtC8vXg8iM3JXyNLYLBMWxY2ENICvesci4n2VGYgFMtyce
uu4L7AsLEQw6PXKjE8zPU06C93PoTxv7iJUQLTl5owrh3IkqdmpVEqg7A7zyGX+QSvXMoJ5Szqvu
hxKiTMtnpGU86I4v2N9tJvQB35pDxBHh7HYqgXALWGfT3QyHeKncRI47PTWqi/sziMjzKYkkyBkW
WtonDoykzmei6G8CrgVc0vQwLdOfsSLYyz8OuqEm6MPwjUpVArMV9X0dXbkiI5erIdkXj3xlTITa
QIv1YwPwYL8eHDc//X4HsVFFbu5vkUsABTkarTwcAuoFT7nMMN0zyzL06z1RuDfsmK0fqu//bjiV
bBXvSeiaHsEjgWHIUGjmGxJoWftbYTmGitHbewV547JEhMELNvDb+B3CE05AaiFjfjOR6/uoqwGO
l4FQZ4N7MR9o/wtEKd2+GJCdFQNFFa0zpERISXMn1YpAhkGQfDJpmW58SvZxxLGO8YXopeQLOKFa
fl7uEc6Z42EdryjtT2Rm5JqS7FU/akC1LYFfl9htHWxoKRmUrkc6YbHGdAzcSWXenrWC8yG1KpG3
WD7w6wqZsDcdqnq+8Bz7c1D9hLwQWRzGHGhJie4Ddmj5TJNkEMAPr5MzAIMyrOg2CqJT5SCjAGUa
uGdCbVWFyHYA2qI1KH21SwE1sxhyhgEqfm21X+EQXaQ+LzZK0N9y2nZshcbZDldJFrAIJD5c+49s
Z1fJS3VIDb5oSKh7XlWfEfgBPJKGUFbcQaIUavTVSzFDXkRNR3GnOm2CC160EGTRuwxP4uZWdNmw
OtuCFOZAPlgwWqXhTgZZOlc7F+DpSHXOXV2M7WO9yB69NBMyJolVAynah5/C0g9Gj2auXodeq0Xt
gEosq2GJwZABdvouvCOCLP1/YQ81y5A0CO1qwomQvdiZ33BJ1v0F8eVNl/fmY6RGaGBL8lJf8hgm
qc2TQgSc73N4claLLCxpJWL8CS+zBapGwDDeaQiQ0y+REYx8fUXY/pohJaGkPB4h4PPszKxLBjVF
LcuDhofvkhaYka/VyLfQqjzIYtAJZ2R8UOVUhRjTd2iXbhnRhDesgEfPJQCIZUQnRiZB8ncPPYqM
9q5WhytuAqtg2u8gDE8EY3iPerLvBmVwpgoNfFk5OhIkNe4hYV5S18ebZHEOHPOSJpbhRptKI0q4
4AGTaWVmEdRHPMtiuanhYOtvzNLkvitmQOCcuyOUYmipQCm/ko/Xj70YxzICUHEoyhhyzsUWviZT
aUo0fjRxx0DFCNZd26WRgYlW8PhLbe0RPGsbp7KLXp5//TpDpr2KhueMZtbJiz+p44FoeXkzheOG
ZwAXOQzEbKTO5oQZ3/lidNziQLUQedLGFz0sE1r1Uc8cjmw3PcT3ZN9FENH9CbLiHHpFsFGhEEiu
9jlQvsLcs7iCxP+SO4acirsrax1zaE/IGTigZM7ZzWvM1s+qfroUocqslsEmeKlKJ5kxgGsDQkSC
PeO0vOkzDqsRPj1PGsiKkomaGaxVnmkX5CHBt99TB75PVyJB8wmzNFMkxcSo/X2Swgbx7iqLlGeK
JlA6/k8vVmHOkMnL70YWRVxLPvrymeDkLuTZARe/RzlcuNyPamruAmQTYIZlU0GugJHmMi3BDOUH
uTxPZ/xNOl3JGRWcoW+SZ7AZMYwJoL0kdsGjT7PcpE93mItx0xowtwus1gEDD1FwgndsApqEMmgb
KiQw1EdISKGDE8jl/f1qAEiLdDDQ+t8svV5J0eLT4SkRFKYrt0FPVSb84XrDTLxr+9SV1bAvq5Ds
ffaTome3y/URKoI+nJss1ZVo89t3O4yQImcg2hOvF9S+5Be7CKEcZxs1NfBNgOTfsbYydLcknVNL
Wy7W01nkUAZ/n5yGeqz1CfcJy4QO+j/onqlZ3ytn0TvxzE15jJ9/q/jyp8V96BtwPpmAqOS9Y+2l
8jEX/i3IvqNDsMIHB8buXXDi+msoZmTxJnxMbdOj/WVCcSFTCv2aCt1WEEjrzP71C8IVSs8TVh9Y
5D+bc/95PL0Nq7hgdAT9yKihY8HxkQC1OiZGhMeMAVauWuSPdfZLJHFVNM+luDkOC7w9bPj9DKTm
6TxJw/Zdmx0spJQ39gnkfLOIkDaTK4SkzV7Cdq1qjxgPvN4Jn29Q1zjc9TBQPrpXi4rPIteXGd3Z
+WaPp96AX2Q9pv0cnCCvbnzXOZi5rGsZ1Tw/KWAe9QU8SdqoQru5obhGV08ouuQQUQFMN3RbWnH1
hZDicboTpI5eJC3A3aZzaFNnuhjOzI9YNyejeBad9H6YiD2auuCPMjy2haoQPtSLNhCuKwsfHsfG
Pemq8zLZDcFXnC2qfIzpkdC8VxPXSpr8rfaCeY84hQSakiN3JRSz0LRsuv1c56xKrHH0nBTUlC7e
9SJ2zZYVlqVzqVdTj0hsrj4ZSPDsadM07u5e3Aag1UtvncgLWU2zsPD69vMRPh4ISmphm3bw0BQU
HS5aWOqU2Mevrd4fiqnUL16qx07ei1XlJLCRvt1C4NL0ZHF2sGhQEXhAKKlHZLUVskHcMhnsfdZ1
qB1CIkzSA+QFdmzXWmhXUOw6LK2UqN7CWEdyUFKnW/reTUjwfHFJqmzSdk4DTZ3WlFvja4Udq6XJ
rTfmiZmSfa2X7t/9kNShlp9o9PgWm8bxbF2opIhxLaDWF9BXzs7gSdTZaUte7WqqO7sk10b+7zZP
blLPr+ih2TyvpeemZbJ8oHm7E4Bvcw/8XTDY9yyhIkG2pgPVtpjGHyu9jCHRLufVPUAvts0YxSU6
7UjZ8KQGoMxuJpiEqilznM/Jn0G6R36uIboc0BJxTSgxfrApzoRF+45HkXlBrNDTuQpCNJ2qXm8N
o9N6UpZO6QO6KvtfDlpBz8azXDeApm0G3cJFlf47UMoyPXRGIU3OdtVQPBORAAJteoJ3MJnExL3l
8p9Q+HODNCIX1a7ZWovLLImfVq9shbLut7UeE1tArVE786ICORsrO4ta3JnJ8+bQaws3TeBrWPRR
EfwvTda6K8/246vlhx9XYXma/VZtQARJR0MiQGJQiuoxfDzImeypLOePzQzFkTRfgPs5vpqEjA8j
xjI9G5MXtb31z/1iYhWZZB7G32TZQW01x2C//aHzRW2yAyQIPXaUuaRwE4dNpguqn+jGxoBfxOZ9
NfG3wAj4xYPHl1S8QCye21q3E1nZ7FNQp1zYtDjKwjEiSyD9KXMy35TipNNitCDDBrxwHG7x+b0v
VAVy6B9eT08l7Ob6JvnwvLqpqszfdrBxqGMYdoRqFcbpZ/t8kHKdET1tmFRAITADKf/QjTF0hyrR
zNkU4zx+/LzfVHCom+ckCJQRYL64qR31xEJRSh49hMLO1cCMKlHe16bvuEPz0z3AOkZ081UMXdnh
QYGBhgyrPJfr3pOe5lDrcF7PpfSAG4Ylh+9MXAG4BQVRXnLkuezBOuroc6Q8VhSy8rP5n+guVPgo
IlzVtyNOP3MaHwV42SFY8VKX8ajg+igptH8orwRioDTZHQH2WWu5SivLthZ9Rk3lIgLwnzUe9cKb
wql9XurDPdTlO5FG8wbLMDHwDl/ACvkiFvfHbZIev0yXk0pRykr/AEpSNEDowOFfdEwr3knbr8qj
4//N1tepqBZyGKUrIrvP3btlxH5DXl45CUnABuLTq8u1WGEpYz4T+nCmZPb/0skNtV3NOAEVNfz3
iy2Kvl0TT+SVfQ+NSooVE5Fl97a3bI28CCNAzrr2SpE0D9Oax2AOlb/VQMSaR5GINVob4yqQD9Sa
FewYuna9GrmFt2pTLiMB7BkC/eP8hYLCyoqVAl6SqrSDbRtCBLLwU2mEn5lbP+cwJ610dlaspCL0
BayCN7v9RTtXIvLl5gprUBXft8rkjLDMLxRS3TsqymJ0kyHhevUnh9jnWBgOtzHFArzjLY45dhE/
q5+jW+OxTLKNFCms47JTJaIhOit3y7Mn6RkzLC6QvqWVwzUKyc6QRhB57scYZoX+5fcJK9UWzCyb
Gc5uQhP/IRVuLgeAIfA0cF7eQcqGaq1eDSSvSPA5sgsEfF05yTIbMvymmhLwnwHZto64hovMMIJ+
BDxjNhE33Ep67VWN/jC0bsEnDl1WFAxegr7jZtHA+49Y9SJzyH62YXSEwiYTsmokax7XNmQbRoEb
QPDWMkOJYtK6Ayaa9ryN74QyZeanz8ADTliksmFIszAfLfXM4cDHh6qBYJq0f1xeggB0Hn+qYlqs
rW1gRCslfOZKfpbDzA3iAK08ouvHHWa5gC/y2XuulSDBLiHJyHFCrvbS6SZY6JPDTXTDThKLl0VW
OKLnjgGD+aAT21lM/5Vfc/tV8euECV0FeLlfaVev9+HEwWoO+atvN/LUJW59uy32T6jkqz8cIEME
qZiHRq13wmS4muTluGy8WXsonjVzrr7LneRIAV5HcvApq8E+50lhFqqJxO5tHBI5Ue9QYl9YNX35
woR3tipHQRMPFiFnGUqj/vJLdAiG3Uptvg55Gu91un4sQLSARi4rjwkfhEjMJV+ISGaeVEI7WMml
RsaBNdKY8zwxxxorhTjfPqLMJiCdHDjN4mblMyAc0/lBOiLfnx2YnhCPQwP21fQ2EodXSUC9uTSI
JjsIrLjylcPR9b7WwcqTZdOzU9T2f2+eIodCx36CRsBkJ0wZmVHy8tRcXpETAs4WWFN8c6r8PWY7
oElqTVKzxEJfy+PSaekyRVhZ3lEUN85kDkxeg/YjIYeSEQwLMQHUeWvSGaVdQTE8e4tPV8AysVbh
gwUFIsq7DkWog7d2gn/U1aYIHmik7VCIlk6bEK3llKKzOC0T1k8RWvBL3WYepzFgR/x637FSkPQY
L+TMibOYDEGnJ3LwTcwegMThO5tOwxIl60SB4YBxansZ5SIytsLwkSADFM/80JevZ1LGi3yV+tPH
h/36g2fvHNHYL5tG5z3aHQ/uKBsy0JVe49sV8bpze2S/hRDLhXSy/7hq8TJ1gvLXUDWJ++mIlxvf
q/ACd+t3N4/pBQq81yNOwWBtfTRnCyE3oLORySbQ1onfSAfIn4rgbcoAzYgEQSLqasIz/gEb3nkH
fXel5L/eyiBeh6dhg8IKf5YdDL0pBKtJNyuKAKSZ5KWaQ++qopKH7rICjqk0AP0f9MkpyoW1FFW2
OSh4Ad3Givv1NCwn/xqSjmhJgyXJraPRRHSoinT5v/DNddj1Q7/zOMHSYT06jn1oFLzJdLsXxZPk
EMdzZTispKuokRnFiTN16XQDpcBQAnhm41M9HCUy2x/3/9yS6Y1h94oSdxJ2moEejK+cm945XH83
4i5YQbHten+16uVV2KfX1M9rhRi5FM4RXljZOVSQkmNVWQvo/Ikfl39dc/aqL2EgLl2u2GCFXbUH
KO1l7kWtGxex0IxVQHmfBmJPHK70yxGeuWDMQwh4jYd6gz/gWt/SyQemWwVC0z4ciO+6jrEciOmH
5APsG74BIn63z4XQ2BlCdcmcfxsslhi6/ZN3B5AR1L/L4WzjDucoKmQOIFkMfWkGaQ9NKY+9M/in
CUfV7IdkHCV8t0L5yQ5WmFXX3O8L47T/0vwca+UmyUj9IQ4sVqZ4vG4I/7U/fbn4AEnPYteyCT1/
ODuFwNNUjMNvuuBxpylFF2n34Psxj8Gq6T3Pwav5wAxm116WKZupkox1iB6tX8+XXxDqjW3VYHoa
ZBO+XHZ0ddeABArDA9jcyTqRqrDRBhOvjZvwiWSXJXoeYG5MmDSZKXaAGEsrBv67ZoKUvDyBveQr
j6f53m3aCoff5tEpJC7PwL0gCm0NgsWiWi/xH3lyRBre6+EuN1CsSr8m8CjcMkGrIcs9rC2UHP6H
+cQmbY6EfSokhaBQuEkv+sUfuetck6PJ2LgzFMwW7YEE4RwhmzAOnt0fEc2LLc4OOk5T65gNXR3A
Tdsf1XKWZSxgNKZ9+yxbRYC6T9CbUiLE0OJTkiZQgl7Wy3NXXGvQ7+KcxaPe1vIX3O9p+kSm++S8
dXeVD/WV1+InBq+IrfhpvqkvTZj7boe6Ti9oiWHyctsFhuyrVEybhAVN0hnLAAEdM8XPiArDtvu4
+UdWDMD7dvanigQkuD2ibaBsRepOslp3B5hFexfjHkBpegiW2UUFRdPPotP9c5CNdjpIRwoj+ECD
mGHqynU/MnwmPmcnQ+Xk1tv+GNmDo731GQspZ4SJ0Qbvpb1bXQVMs/C4UqUhnE2wLFAIZXlwthMM
zGvJjNhWg/xg+pw9GlAB8y9olf20nEeiSqlExnCqerbUDwo6M7R7CbU62AwaXi9gDAVWVAAOByJh
DO6vtkrdmnTIE7GBkyZkFmI0uLE6jtX/p8bFOz4vZCUqAObTRDHoKo/718hLRUxwo0Z8EaaSMu4I
qcXvCZGJQjQ766ZC1+uYLK0yLSObnPcUo5MAQDrNs6wzgmnQaSv7fywx7fUGgBWiJqslvrewyRBE
Zz1cgYTOOD4wOunPr8aRpa8Px11lj1QrakTjR18jkhaVmHcbJnOxsUaCfrUsAgJ1wUHPfhB/Srfi
QmAc2qER0A8pl3PbYRPG/r+niJFI3y/vsW9Y78mCA0VBLe54esrsuw//dgobYkJir0fdAAUevzxE
LpO5RGGi/GsJjYKLMg0WsYZ8lgzxv5E8vMOFyixa3/MQV/CARn+ommHh4s5pquid5jRKQarPYKDJ
2S00JslJBuKMbZrVt87n/Mwp5PYVG84FKYhBWdVGXvVguOVj8WGV0FesWEaO7U6hVIpA5pA/3sDN
8nEtouAcNB2JO3wbVp7Xg+9f4ytYHyEzVwRt5H0AcQ4SXd6LJrkHaDdV56aQxFSQRYbUjA/BRUta
YZet1WUqONJR0SiyT/3AK5BBSQWaVlaot7utdIdCV6fIpqiZZgBpD6rxpmWrPyrRbVJO5hsZGNBT
Tun83rLBj0UaA1fGH8yHgBUUzFFfjqQNqQ/E7dZ/oYpKzKcbZATkukBqzhceA9kZw6+mOTbiL0A9
a7S+RfNzrCuI97otrWklh6q8YYZ1SpsjPwl7rGJ2MrCFjbJ3ijjf0cRKfoaXD5QoaaDOH3SxdZbr
LXkY8pP0uhs5pEt6LsXlfbeCpVFm08JTkYvhyIrDCDUVC6F+agxcIJstLDBQunMfTBTosG/+FlXo
ZL2B9cQCoPbaQ+OhlV2XlIDAqjY0YsE3PNkFYA9GGuKC12Agds4/5X4AVMtg0tdazqSkCyW2A3We
LlzLkFro4WuORxZgbwA3GE2OKwnmZUykFnlZZqVx0U681nFu30NN+nZs3b1kck9uHYBhbXNVHsF6
5D/kiivuJEDhrfYw8AR1ilcfqRs/yPbeS79aPoaxQoQE9Ow7SVlq3wkV5oeyGdjPutjEEpv2/8hI
WFHTwqVWJ6gh7CngygDvs3ukCYpHFq+/4SZRLs5cwX1xmQOiin0z0TrHSAxdyqfheEadRVcjimNC
+jPwWNarZgcz0r6bgMaUdCIplBchXMXb3jbe2s1BBHtf+/VODvS3cAEIfKmyn5fG+727uq9XAukh
vQCf3mgnDQXWCDfhUZhdy2yIzlvDPtMscoktvekUJEqh+Ly54906depkpTvUh3l7cBvtNNUVP1qx
yIGdYWveAxjeV/II+kJGsPMV49IZd+g+1dHipgGpAWkamjlXn1hPw2WyNSWa5fvDZ0qu67yUwO7P
Yj2WFPr5HkuegBGaM2Z5LD0fnvE7Azy4FbA4iK0yQ5TXh3qh4OmJXMBDE0oLTlFk4GgiQlrPTPQi
n5/RJl1UK/BhNXACEzEHhbSZNhYo7C61H0YGtjC21uW2p2r+IoiLzTpFC0D5VN6VDwGfJYAmXQAh
QzdgjnsvLY6jg7aRQUqn6IICas3xIr0sRBtMbqSuYV2KWi3WX0I0Zfu9K4y6zoYtp8WwVg5zEYVU
dlAbW352UjZuQ+LCLs7GGcMuhJttgJb8ckSVHGP1Rms5t4+aVQMW0XGZkPj3CAI6NVGvWGe197vR
SP+q2ZpxCsEQSimS1oTEM3cbJzJaLL4HJi6spvOaHvqBhjVcPQJnCTKVZCAc0cOiEQAg+3cp214l
Xkjf5992AxLij/SuFrbTELI+oOZ+/wlvabZH0oOQDkLhwgSSYIrdyE+BXPLwVxJanjE38oyQtf+/
yQhwVgwMFhvZ/GqOaIhYwLtIMPYPUnKKcMJx7cLElI3PRfOH1Z+0xlCxw9JlyZhSUVebb4L63wpH
FyhYa4RyRqSbx3CzPLbWJcPSfOuSUodSsFX00If86B7arhO4VO6pypFO7EhNQUzDfD/+jQFSvq8q
xm7mFrSkR887Q+A6WN2YSbl8MtNcMas3tt7zScRtXrBdUfxGMJVaUYUf3sgLk0GT0WVsM+Zc7kQS
mKtQR/T01e5lNk2N98UJDZFDrJLi8GEx2tmO5IJVM6Netti4UT4ahJcLvlv2k8mn38olD4jfRexP
JpDquj5qTcar+O+Qw7EMXPkaISYQW1KfMqzWvId7Y8+OWzSV1c+hAnVj8dz6xiB12aANn7oAL6/q
Cow0ieRj7mxx8GfLIyCHCjyy1BBiq45nCjMQP2qJHkFhyiUU/dVxMPendLRUYQH5ax/fWA4uIaP3
FEvodocE+uQqxiH2o0LCAR0bX9VyOI8NCum5F2N1Gi4k4aziz0copCI7JYSLIRBcz2HaXGR39UP8
PIrB4QASLtRFQxu4q8DITho567inO5Gpkue76U2JqaiGY2qoCi2pNLviUgCZavPGx/9UubB9NJoY
BaYV/UcybVukub6FVjykL6xvI2BMx3ZomYc8VnLggVcAwDisotVw5rCzCKmJd4Aieze8A8s4RTWz
Qlp5Gl7JoIWTrN244XUZcUD4zGD7RMJwopGPwg4S+XdS6pQPZ0R5QnFY5ctzsXA0sXHNKOih2YNI
wshopAFJpDDJ9QcYIeo65saZhD2fqbvWNlcX0DPFOb6OKXxXF1ar/wXARVXzt0ibrsOsdyI6CNfE
4jnbd/JlzbcK6O0ph3sZRqR9+HGtUXGwVAKwXV4DuAHK66lVqSfyXdvExx6hklWpC1ZA03/yTogj
WdQNfjfTOtuWRiysxG7NsMmuQIGYV34fjGgaetUjzTNNO7fm8g3dm/H8HYKP6C8onfIAqVFuKvH6
EM1FSCRJJ8k828/TMvgAknltE798H0uUBgeJ5NIUJo4Iwt62FRioq3nNZZiEb1g8vJDWeH1g6Ky6
559c27xp17jsHxmtBY7dkZMMzRNMMq8qYraZQtSBZZP8tVa+RFv/qYrVn9W+ndKJrSPOGPmp++9X
Gzl9J9ud8Wgt4FWVWlkSxuPA1IYsMw6qCE2A/MahvtJJf/URXjIUjWqi+nlHcIjxWPmy5lvVVs2j
bpaZK9iI5iVzUHeBwseFIBBO8VRAbyFpXv4mdaZ8KFZfvhZ+PfSZBkmN1r1nfoiG3qVxz7aUzbUi
7CzD1StNsSgdohgSl2EOnTO72fsG2C9/zHFHxFgMOzf7yU/v+iDJ5oFQKZkIi4XOOYbKzku/4LlH
N+KIfkObmus03dlvXwKwehD0dsGbqCPcgIlQWw4fjgighVp/6xVoCKLPm9dc8avsNzXpLVtLML94
XaNpRCsSAdqbtZ5hf7J0mCt5u6+z8P8jV8dVIoKJovDpwoOkdXPRMKLVVwLGzHmkOOco3f+6D3yU
9I/rGV1yYO66g6FXac9wtLdGARXW1AfLe1eQfhj2NAw/WqzHbpPzwWTK56zQGbWJBrgjBDChHGO7
vC0ULdsKDXznKt+9aDdGulEnjXN3BCpqVodaQapeLT+tOsOD7Lr1C0wvzZbt2Y+Dmk2H8Tlp5KX1
b2RBb7QkHh+WrJJFhjqyFeyFINSEaf4BYk2FNFG+Esoe2rjsrg8q2ySveZzCwKVnkR59H1aM4Xjt
iI+KA3cSY6gw8dyi0WXivo1skcG6zirKROuq0hWK2hSxQkRlpz0XoERHz5Ceib7IZ1cMHk8H+U7H
ycxN3j4ueMrFc6ikHEyfau1WF+b1pCc4BKG2qEBV7GkKwikO+cGRTGQI7m8iMm6F41QO8CZW8UwB
U+8AdpJf6dyv01YdOBrpewjIYKZY0oU/MX2IPfx5Atv8mYycXzlOdltgdSUlJpLXXtKw7fhbULAv
ol5MQIChY70J+HHJMGTrev//Q1FPH0Ag9G/VmyeHZBO+cowS9oQKEL52MyHNu4vHWcsdWXS736ho
TukM2pAxakyXVZ7lZk/0zoRZXDWdQCFeAs3/FfRpaYo+r8t5AYqV+AsqQgpxwcfyceLTSqppJZrP
Wx76RTXnnuUGbJoPw5KIBpse/ZPt+jfS/oZyu0XllHOVH0YbnVi27tCAzQfNUK5qwn9CWZhLwAIW
Yoz1gIg3IkjBPYzpifAVBg+WmqmnA42TCbPAMRZuPd8vIUOW6TyG56bkqWELpq16Y63pPWlmqNkt
i4Mndoki0L54N9wx6pe3mRdB2Nqd4KovqL7Oev1uSblDEftKwI7+v9tQa4x0O3Kj11v3SpgAyDDh
AAx4a7K6CqGilkXjn/dw5/YJplUxzB6sMU2C8FnoiQ58FwAVoVJF0VbUGGnDgO8XdMGlvBQeB91Q
Ua0ucdkfYt1pwwqIwC2hhq98eX1z+B7XLvY758I8LzfZi96LMMVnAJqw6AbNtOpL6wOkLmUy49E/
bYbYRKHv0LIO5QwvyYvtYOywhHlrF6jEKsgHt1vQzKNl3cfdPF1EL8TjKLeR2ba6YqH4QENA0EK5
dEEVXxRjIIk1DPhYj5B7hKTAH2yzYcMN+NnSV24QlV+AsnvmHLmGGaHpkOcp9AzIEYWeiVzczoLn
6Ya4Ch3JXaT3HgdVhnDcz/4ZmeSFwxxaZ3NPBE0BCD9xvman8jnccOUCRX+omvfXxmIT81kswzdb
F2XzDAHEDZGe+3EvOkhafrIJlL373VctpAvY0Jd6JOQtogk0gwqXmUVp5G4mSUDkp/pHoJRJwW+r
2enC57qKOE+denIaIwqBavQSCwjAN/S+gjokJea0hO27+5HIw8VHD3xjYDMnNMo5KB4+LvOrrNcW
DsSXJX1/MAnLaC3txL5kGSrtbI2Nb6oy+jFHoy2plEodCdYcXF1eTlGP/MdKb7ul1tbCqqPANHwm
qkcAtTD0bRJVBUOsVkRTnzkXgo16RzyWB3FVzjawqZuLraW/KKFTusyvYSTSMK78yO/tiq84vFAk
6wvyOxcVKUSCPwoM+Lq8WMg2pqYPDc+xkdMNr3wNjsvYV/zJLeaPXmxwX7zr4nRmh06j974Z/psw
kKoAXWUX+HWBo918rkIPpmjlh9PBJz3x7PLOILNXH1OY+qy/40jwbT0R5S8350o/eClFohpFOsQQ
i3tmD+y7GX5zPN1ReZmHUxk8ehOVk6QKL/Yag3cOIJiwgxB0f+SpURZ8X2ftAcNZRtXAFxDm6+my
2JeigeUu28EaW4Jrhi80TqwksoH/PFyuqt1dyQIvKPpA9EM5bWrLd7yKJWikZ62lP3RFExi85bgY
36VwA5Wf+p4Yc9cdnqylYxOtOW3CVWVoL6yqlOmC+kmpO9cmaAiYyTHxkO74C3ienGaOr2D1OMkj
0FmYx0iS5Wq1HTeldI8AJaQ4HNeb7AmjMVC0/lbOHu8m97XzOnRGtrUhU7sbFQLgYY7mv6tZcbT6
NtVyuFETjNZuHvgzNQc+jrTiOi2nysnyroQxxN3dtDLzollutAvVpDqnKjqq4cU3kBfGzQOeS3oB
uyzpABpmubQ3T/GSKmUJWJbs0ZR6aMdG6s+Fj3rqBlk2mWSyZ8CvOjFstNMwsugHgJVflOLfG9jL
BjmioCPGuyoBssROOdCYLlYq5D4IT31bOOUNkq4u0rHjcalT0pqKQhlcMylCu8TgPvoJ7GJOa+pV
ESJJmg69de7H8SKqy85eRxOAHMitAdHS8dcE/rVxhGofpbCW70vqgd0+FX7+tvPTcGGiw5VJlxcL
2DPptPb3Gbzd6x/KAOgYrB5AlgW6dnuVGdkeTx0LbyUlYOHT+tW/1fxgiYJ6SN7kIIUCUKNBI9qG
Bh5exkuQd+SqC3rnDp08kOoRZ8H/JR/lh7gRmiYSzWe2xZkBNdtwFxji7235byOqfPhLcET5Md29
ew+zcsWbvjAHrILv9yCZhsatomxOyyFLB3cHjoqW6eQrGWEqodWfDPHkDYIi4SVgO+zv6DZv6Gr5
drx1kW8wPb/bBIEwN8Zau3D9XMGE+7ULiYBofB4UveFrin/uJvG84d8Gh9a6aqRzIiYJvTZ2AMCB
xcj9xoiFHR/0Mz2cpDi3EvOPaaBwFcroeLpzknL9EUxi35Ygu9IcK1yJQ8IDzUtFa91pxOmrUEGN
0zrbEmCKKjlHoNTQAykMzWRUq7SoECwjjqpWhOT9R9tUJSF2qef+Pw7ncet82iDDQC6BOhfRBVOA
ve2N5tFODNTLsNvMcuyHescIavpOE94rXtjLuvD5iqdf0NcbUz9gCIaSeBkLg66RxeSNDY7maBKK
DJl/mRVVh8ssm4i3jl2jElZVA+htBZqwIyit6odzKrZoZYhdrf0DxEiV5xM1U1RynxrlBCxywqIT
1Ui3SoviDsBlGeDstc5xVOmIYd5fqM+oxtk831ohGO/wpwte7Fj+KRoD3uzJLr0AfANxmQIU4oe3
pw8B7ycTZVYm20dhKpDZTV6z9XTF38jv70SlvlRtFxYWkURbrB6/rmW8baaW5NQqf7VI9UNTxCSD
ClOSnJkluFVE5akCU64aomMlUWRwkx1UBF+WVghzPotnCjNyTKbdpkMWplUpspXqxFPkORYV6FlI
qaQbg9kcXzLMjBlUJIW5ItMl6i1xfFjcGA5AyMbnLT1rHrOc3QjhoWUYxd6nXNE/WgVWubnnvgQO
kGBIs4yO+0Yc65X8jYJzfKRcbgyYk+r6/SzoZwBex6GIsyfzQzBBLa9Wp49Q8UH1fzQXkMpGFeX9
KbTZZ0eNPc4kheaTYdKSkHE5odWnTgKXu8J5zaCaiyJfCWzUhZxpUMgwi4RwcNkK+Kv0L6c58uah
6XXFR4WkclsuY+M9DaRQIm6p6m/WYMPhv7YYnkNgxW3doSlluLzPTnF8X4pdndIFdItAw6hY3Pqv
1QveC7pcZVOxwpeaM3yXt4Obh6GkiFqR3+drAtxHhlPpbUE6ZXvyIWpBfFnTy6n10dABCo/kGUIT
BWC9oPssKrGzxdwhhZULE0mZNX8Pw9ckGdIgyw+mFhADorX6ezwZU8VrM9WhSJg6eTfv7ZHuqNYl
Z/iEvtOqVaCoUghqfxD6/QOY/C7YKZ987oAf9qS1U2dU+xV1H/rTHP4drBNUaslr7Jp+3V4B7yq0
eD0wjEh8TxA1S2CtcUBXc02nx/Znj3zBPe27lf/0Nl+Dtq00VvOIIG5lR1hhnLit6QCLJLAI3XM0
MBUuqTRjZq7flk7v3raxPJFYFRoKh3Qz/6UAo/0/YmUMuGgBuN1yg5v2oEnkFlG0BhB+ktiODDds
81vFeUZjgPfxuh9tRe7YapzXUfvhbI0mJRH+EcPAiMy9PCDMJQ7/tWUs40cI1H8kv0dA/r3UFnd8
h69SQcfV+I892zs0JRH+tP4Iz+59XBq2D+HMejt1n5YoVtUU50UWILvLB9nzqRAszf9WJD9bQC+7
vbsYktLT2oo4L29Ym+kmoxeMnLPdJlW8qe5pSIMN74a8Z6F0rXb9dx0ixWon9KJkKxqkF8mWcN20
kvSL3fVXTmi6qxOcHcp0kHluRMI2k1epGGK4LoWWDWo1Cc5A9FDUItJ/bsa3+A6kFPfQZkU8UP2w
81G9BBGRz7Yo9e7h1yaaroSsd99bTcuFBea6d5GIAd5s/3Ty8hXUwoN7MYd9tZZf8SQRKNYY+SbF
vIQerC/n9eQOYM3Qfu6Zc+5wcBjGhHnAoJNA2n6fpznVxSB/plMisB3LBDlkx4vtWzZO2Dv5jP0D
Od4bCeuXm7feTYDndUBaYiqrRp9omTMGeKCzeM0J797o6J9RZ3Btg+zIgcXnFGvW7xkMW2Db1Kpd
sQ+BXYZZK0fitQSSNZ1loTPTAz7SwMsj6hv7nuOPjArJ5eRxKsDhHfHWew6zahmkBzX09XLzh2vy
t+Wmz5hfiXLdjBSJCfaV5getW+guAmpd0dfxb7H3Z8quqqW8MAZtLYHXib2tdMp0y0colvPMyws+
9xYoQGSCH1S8hcASatRFQGh05AOTt9Sk2doHg+Qi+peI0/Ean5PX4k9cJn7UzhpHL8Rl1mQDPhnj
kIVKjQyeVyOWMnpydkCG11VaINC4YZ1NbZR0xTl7LtZIJmbSMkqk3Oy/7KwdL/fk+H+sad9i6aLE
kbICKpx+c3zbeZ3v9h8ucJFxZEfz9v22dOWwv/Xa6dWUTqK7/kOKTNkj6ncSRMs+VRvovC2VneIr
liL7A3fYBDe7gFhbVLZHQVrtvm6NAB+RJI91nopL/LtXRulLDrf7MInu8VE+7ToG0aCUxMbMOGdJ
9U52N/+D3Op+1o2yfJhr/KbZRuLHBjpDgJNrArISmeL/nkGGeKYBegRylsjpRcN24Fo97rfAIA9y
bNMGc7wFnfAXde9+r1bljbJ+BW2uTHdD93+rOncNii1XMOqDGJnov0JDtl0zWRtsUujJxnQqe5ym
lo2iA+wdHoeBX++ikfTQVYS4ICvvV6QMa79vAgSkEgDulPp9vdVDoPCGTvxBuhK2+VaZUMRsCTIG
dru6H5uodSRJuo5esPPzeCN5JfrvdoNMS/llIV9dtkOw/IpRxmHYMR+xJ+PUAK7xAe63tDJ0fR21
UpLgywJpWR9oYuM8BhcqsCb5U5m4+PjHhhIhWsBCEymvAvn7J73Ivm4j0wWNZsNabcZ43idSiidj
QnMDNq1Ox+Uzj/BWPW7h8/cHeQGSWy6jt87dwg2gGWB++MW0mAHyYmZIFjBKvi6dSc4A6t8c/cuS
BxDd/rNcjkzBhJYYrbjkQxB1fcGiSl2jzUDpVmr+vm5rXcNJYQTtxch1au0x8Qi6nzkCj2XG2iLX
+R+jkBUAARR/sF+mMNgye1t+Q2C6rGVo3PnQNPO43h9TvEJB7Vr5JxBCQ7dPmtNdelILE+kPP9+6
eTe+cMHdoQ+vpqsXUjVA3zLGSOdTUxiRc3HM7wCOSqlIF6h3w+Z05r/V5S0vRjqAAJEtm0UUejBl
PMj81djxJ9voD4ydvyqp8m6sIdXzYkroJMJCjzwvr0kSmHfZpf9FGcvH7DGrrzvXN/kI1HVQxHVz
21v6uHdBRbQRIe+FiMDcLjoxaXxhfiAKW+DVLCf2VjAvTPoaPKrY9skVacm7AQeqzqHcD7FVWpxU
J40XljNiRv2CpmV80FVIpSDkiDsoQpUg0I0yQIX0SIwWuJvBEqYIPq6ZzMJlE4uFP2NRPMELImRy
RaFl5lt3JOTRo6kGkjIFLjDcn7psLBcIhnYpW8eiC3CGvbINXQdKpYGx5EOLpFIF3HXw+H7lqhjs
Q620IWsRyqmuvgnq1IdGHLRboe6vMV0eMxxN9/XExbB58CjzcNz0/67t87ivKb6gxH6zBL/rAGcX
sbzY0zzB6U0pNecvCmC5/g9muy6BiboIUmPHoL273LN2iQaV/4Hk112i7e8HEd6ksIQVZ8x0CvHB
ENU5djqqsNE3SdunOKGjp8t4FtG+xbD3Es0EmlT9xAqykzQOfkB+UV2SIhzmTE28fqUgXUj8b/dp
m8qxlFND3hF//rIviu3x/Mt0fO0tMY6+BIIiU1MbhWZNyC2mXc2kg9GshqZwgNfuPIL35Xovshzx
AZOIyusHfGNCuGa2Fd61JG+7xmPe6F/IoaLjchaxxJcQNs5RAy7zTZ2Gm4Err954gslljLw35zdg
P9WsdSedqbOXKmwCi9Poms6NHX00AKufUERbtMK6eEyHdU0f/aYVBD9qVjXaRI+GfJwSuEhbg72o
PP5CNUXzZ5ftVB9DsqzoAckHHsyYhO8IvEDaiNW7RTK80YoVoh6hmquaHWAyJ3NQQDwt1JKPVsER
nZilhKIdooyyoeKoYHOZtx4zbCG1Kk0cNB+nNjm+L9SwL15WtpGD8oCH8GKeaAs5l9ijhHyYOC7b
pBrCqA2n1GwrUQfnaa1P+rmKNFLbefn2kWwh7o+0gTNJYaLeJXjcimrQtKREEALgbebqzjdwHuWh
M1Lge4Yw9tlh6LWRxWu1aMb2Cm//GXXO8idI0x7tNSG4JsoHGYoi1oA+SuUzZpehPFBkMaYPpKA8
ZlMMXTWyY1GvzVSr3JYopfQQDVrh2s29pqllFO5hphMH72p/22esPQyyf9qR3ptgmnhLhrIP7E1X
//3e73MDSW2mJLcmjQeNVr0JWz+UST/5PR79Gz38ayEvo3UZCfke2lDN3y493oQBCJk9/YfUTTas
OH389RXzCxKa1N5m9ZTp30U0zgAQZ1KMe80R5GnUvWHAmcd+liOcbBN2fdwD8b/TqaPpUZAIIDgW
hcVLdkINo4HGtBq07zrsb7zdhdPnnieW1XtKcgl+VCPBgQjm0u6JV/1G060zSqeWoWk64n7wR/L3
Alx2T5T/5X+9ZsQld/EngJeo90yIAxktYe3zz15VOHrMfN16txPkH3VWUsSOps7vc8leA+Jrppet
qlF1PbF6f2aIDeM/2oHdpz1f5qxLazC1yw4WtLffcLhgtPW5NrsSSxSSNsRPCrHU7H0st+NOMtaQ
SAXPLQIG4YxOpPfEfcOUJ3wtE6IT54ta4LY7c1VkCgmkHtn7QrqPA4XX02DAYhwFZlVec8JFYzoI
5Oce+35AJdqJxwbyFZl5HELH/beuR2zXDRa+d0g6aNwWfVOCD6YNdfObxGfe9m+NhNbuFN4pnxPr
aD42oIkj4DMb2H0YZtO9J7KiHQCFKokQ/tHx/Gbq+mIlA18B/MaFGvoMz1lyEV5uHU8CT19gp3Rt
ctdjKmHijqd+G8/EBX1sCNgiM7dh/t6LzWzJUs0wnd9urSgi/YFRSH3PT4qqDXlPiPIUiAXse/OI
yjPKtllQaHe3S3Y3MiIFv4U7ZseEgmpoiaaOg72Ujde5Yz/0FV0vZp6PsyJfe51vdkCeEbUWioYu
IsEiI7vCKO+q8W8ROfKysbC+tgVbZ0vjGQHX1sQZbfxRSUFO3a7idj9Ej6GliqgU9zu35PDA63OZ
3oA8USW0XSSp7GQw8QcSZO7hYjoTJfNB8rhzrt22FEnIR8hmLyfRzxzh9wMv92GrSAxYby8+MYP9
8LwTqII/DX9CAEahPFpkQFYzyKb08Yr2E4MpMjtHKAIHTBOtwwiqMaWk7EYCHWl4Q5nUcvf163Ut
44Dv2H7lPXPVHKPOjGUcpVzxPOLnn+iOd85zYARqnXWT/gCToInXN2H3POfUqUeRI6AM62iccJWi
yCXNmV6Z4ROEYGHvdyNStPzlj0x1+w4UF/tLUNizwT+gTTK3s4JfVinZEu5COo2l/xV9gfLHbP6g
c6OjmTzUxfKrklGVo+pnXHmxBF4+AKdpRI0j64RY0Vu1xqHNrY+uhiIK2kFofwvCGL0Oa5lTfQZp
fVDV+ObxfUjudxJ7MJPwh6ChQg/X1jPdZA5IhABe+wiCC2888Dgo5mleC0mYQkoQMpw87uvwTtSV
skbXowVs30I+gGtwqqadCdRUddnkmISc+yGQg1a1eRTSSV8HEtiF9xGysWgFTtxfVMku/wZ5J1aw
WTt6xBMFC7Vba//XYZxAXi9RWtZC7ahqzDujwskMFY1Q95OUTJ4+c1ey/rSnupjTFHh1y+ULjSu8
mzwXxBjZkLbJuJDlZVYOpN0bY1jqfMLWUks/ZviuOfaPHZZTK41/2aPRdge7LsuFMreg1n2IiNnq
MF7aoeLaMYTctKdJZ6/flqOMfc0mm/P9Ms45nJ+cxnsAcf5M6E3wj0w8UqRA0nOKxgdw1wVwpwv7
zUjcSu4bhCeXKyWEFTHbVca1XE9MxQVgkhhNzLQJu4cgJFxWFqDXQE+3PoA2xS8CXF0JHrG6cfjc
0AgtTVHwqiTBSl4N2X1fQ5+J86NK3dOALoyR9csIAHdITbNbE5QETJqIjTMcNxIw30IcLUfQQUQ0
zdl/Hg/9+bF6X0SiNS7a03WqHoDcTwZNDMO4TcgaUv/66vy2XXsIIew1BHQdYgMG7vYRavi5EDNm
nGaT4MoEb1/89WotK2a8iiyaxQAbEl+kbi1YCuW0fOOqSv4Jtw6zREArbbru62q8VORKRzMbJgzN
C5MJcvFpgg3E/umGyde6mgFHNRqxc5n4ZWpLyTKaWNFly8lkcMIXIN0EO3M3EXPb8QlrE6NSSy5G
ux31WLsqwrfiaB/+TDvG5c3CaAAdEted1DQtlBxoobrRgS4aOe5XU/DEndrzUaD8OzEvDNm6yLM/
EdaD4m/LIUmBbj7wSo80dU3V8UhjpqqZqTylzgGluTSsuYaQBc3ZymeYylQGmym6boFx3dwpL3TK
R4EOtifOL5P5P2nflwsmv+gPmKjrVcl/2FDKQlMNDrwntx5u/3ulHUoIwzFBvrHYCyjhIttTL7EQ
oIr0IWWA6HAe+SvihyXDlGPPYvLIt0c6DGuZSK9k4vKYLHbR7JDRorB762Bz9BCXfhGWNiTDPCt2
ZFb4BzVdCgq7HdZIp4b01H3pdKZeNjFnQIFdyHZO4p/8WjeafQTlfFl6p+LO2qIwCjcSv4ONjSEA
10IdhehvfYeDwokcUMrxd0rvEyXu6NhZpbR4Gh5th32x08t5YgLx1fKFC4GDz3GdXPSaXNIHbnrJ
phmfitaiJxBQzU8gPFnPF/lVyGrvdXvDoAhHwK2LRz1jiSF8yx/uG9kdmRBbWcxeIW7+biLZG/rD
vxzU3cHdQHo1K6oL41lDZJjtkzIxH9qJHRhbTLEHLMPVw6oWe+BJXPTVBczAfZtPizFXNgcbZtwn
TdYz9nK6/icNq3KJZifjXUT/mmtTllU7Y7pLoF5ZBgVzbh5wTN0i5dHy+YAG98B0EIu3B+ldnxp8
/jKdb/myh8hx7XEkOVijTdwRcMu+OOgO+lu9CpnIiV0jpEH+BeLteyYxgtl+k5i4tJ5XmdBg4hjq
5hZv1hUqNke/YuZuj6HdSS4yx12biWmX3MTzxqNmKxpwoLt7koyWgI/d83mBppxAi/K911BELmgm
x2uDqqq8T5mnx6agb7myxeSnXhWESpkQazh/lP0xgPLtwqfRe2GsR4n4d63lfMxPgHTd/apmrFT2
Tn2gyAFmlEHfq4BZvhsjYXfoeIgOy/csTpfTy6wQ8qpkAZ6DJu7Q/G6GhTE/XB9b7qfJvFOjo4qV
wGjiwM2TmC5QA391bHONPQSWGGu4QX7K+WP3zBc1xMJAk0k2yaJXIBwwt2z8mZk/MfpSb+F3/62s
p9qXS+cCcohLYSTCvGrPb/BDgzZlET3ZtC9Oor5kpkg5jbJLexvPzT/1uHogGRnnLFK2ULjv6klU
rv20JnrISG9A9Ht0yXiGuG6iCoWVrxIX/b9nhI4VSZNx4FEzwBP+mkNG4QZnEw0oDFOKK6Ml0N7G
gvscn4Z95sWJv/oaJsWJo3F8trhJp36zO2ePeeubEZHcdQyfEE/JBpD2MN8L8UuwUydyU/MQbxxQ
RuaZ2IKZ+ZXhlE3gjNtA6TNtn6WZoOWtKdK/eOdV7J+vC+GT62/fvebnzuCN3z+a47j+7QE131OP
aGMJyGsb5n9FZU4642QL2ni1EKaQ1XJUl6OGZPuuuA4dUDraJuxOnyqlI+DUC3MNxeSxStkR00L4
9wpnQI6+1/hIAWeVC4s5Srgkp7+lHxsMe53IV98N1VV+Dq0DzxLyVJevwcarrB2xrXJ8OidSlTS9
W8LovcFWJr704/dI81nXbFJNdmt2SJTmLXAM8ef7EcG5pGvV7IIeZJ2S3XfORiofXvLWwwUhgeVe
sP6UXiIBQBaL6cqgObJa+n+UcF57VpRmrV0GXPyIUWFRbYSr7YaZ8K9Zuz/LfT0ZBU0rZdG536Dd
byy22BIby5jHnkOPf1tk2Dy58rmo8bTu/QN6+UF6RCmL4YGMDt3g2//3c9RlE8EEslhOD+oT4GgP
PWxL9sgop60CfHQloqrtNFl4ZIT46GHz1yEGyk9QEj6qBEi8V63AivIWP2dSqdPtS29KQpLcwDlK
n9w2j3tHjK384RpTwJxoK1KvO2IcjZKM8/Ga2cTyGSbsgl1rAGUP88nwm110kM1TOATfnaEuZN0S
eGf+C8J2LGKRjS3zP3tMaWkNYeMXgeYDAKnjOLaN8ENGfJ1WrE9NhmR5a0xoVBcGNacAhRQaRcFh
EfDGciCJge2sLdvhyzuODvHLQM5jZJmsmbZgOUSjKUQZS5KNG36PVoljym9cFseg2p3AEYo2WfmC
1FRtE8096NNcu0B/QVMS/qTxfPxqHbMziYX7MfCITXYTtMXIsxyXJ6Q3LU34hdb79tZCNOVKOQ3R
Uxc3DgGlxctCT+Yck7X2Oyv6VOzWqzXGTyhu6muKkSxJD3r0GxFuaOjwWJ58TxQtcXBgisFQvmlO
O/hhmIgRmBPk7vEHzb4JOoahem1b0RzD5UXL4fgPEZ3h7lqNg9cUeuxNsAUTkhrvNQ07sUKzN+QG
aF/f+Td1ZGlGym+zs8tLhOA3WOyxT+T++jeMsU2exCRKE4TayT78wBCkbySd+azF/j2Es/PmQxGm
1+wrBRX4nSqCd81K9zdUCBsR1Pej/bjaCpWjHEhDNOz4xbHnIKn4n/nmZFyG0O92K40VIPlQb6lR
IpCNal0G8pBgqQtRoxew83b0wjYKDBAhRdI86igGC5N6BW0ceF0L8V9tk2t9yfc1lHPHxqhk5rGk
l93c2/7LiaWfd+tXcNmhH5KqCPtQ9gOWMbHl2LaCblHAqXCiFXieJcLKFrxJdEv5QIzqWHrK3Mtf
cG2PtOPVR0mqEjI+gtRO0iQ0JOHkrM7BPg2XbvUkfuy3MYtK8yZBsNUvYP6Hefrw6z4FCT/XrH1k
kHVPvsr1eAaUMkyDkZ5P08NOsDwc3tVYiGGXTm6Y1n+ZPIX5htbjfSGta4sKpDnxRKoTpZyaU7Zv
qlE6R3LpVB2KHXU2V9svCrrktV958WNOZvrmM+nwfb1EfCg3Y6DMAnq6QhhxlV5kBuBfMJbHlo5o
1fjig6s+lDzgCxKy44pv27Z+IgdrDDjGFkAnZCxdb9IY1BX+n2Q4fibmJRtxeRH/m6vXSS+nRY61
nBseJpaqAQ5t0wIrqXlcp/i3bq8A+nPpmCDUE/AzRW0nhCqTBEtUPrTtg9Eq7HUHUGbNDIvPvUyg
t5NaHEsGJRh6GjDE3DDOApzl6m4RA+VeYMHGt5jPKbBBaWhh2nVGBVoglloxm4BLrzxKBHtr1AXj
/krDMuARSkiA+2TFRO+Bn47KYS5xSrmrCRrNoNyVQUSQ/Twb69W2oiM+xzO4Bf9YNgUePBUrebgp
9KO0t/XDU5bTvcQXhLNoUWzVNwqgd3RDTvY4N0MdVHnuFx6a6a5Ve/jLsEhqbWDCtVFMgiWOWpsz
JGQJ3Iw6AQJ6pxK/s/63lJBTUJiFezU5Okg4yIlF8ATh5BCEuCDOgCHSAcKbeJboMsVKRB8YeSkL
x6maJxhFdQr1PANgS1Mp/0g6o1RXPlbWynUfAKZpGG5GnZ5frIuze90LE1mOtFGmKOcteP+CSgmC
+29vfXticbd3JPSz+VA1FBsXSd9ev5isoc1rATmOqCd7dvPuMvB0YwteOtJ0QqCoISinm3DwToUh
IdbrYEpaobVVhjkfAwIj+BTP7IaGzm+zW7YZIlKZTyLwYJJ7yho7fofQGvApI+74zbIWI/t1wn7U
Dbu3lauT5XlIAbQJ5SrGRxDrtsGZ8ZMyE4VYZaXr5/D46/tZNHIndtrYfQIm5EOKJb7FuI96zll4
NAvBJOPTKC1fg66zjxx6knEUE82rAGX3hcgWxlBBO1of9HXlacreYy6RmanpfYapCtYagOCKZp7s
V/M4JxyLnx0dA4lztt0DGfTAEcYHqbJam0aDp2Kn0ljqiaIovLDg2dwISJ3r1HHHHwKARjjWfWsZ
3icszDuRs4UTWx6HP+zGmp/iXpSdpeOiZ/ZuoLE8nN+RGr0Ih27ODvo2xqTbOO5J50pklugbrp5s
yVG74/lkEsc5Eqn+EQD1DfG8kISRghD7TONiKRPjtgkvUng/F8TkSgAdJzBNUPxIzJjwvOYKztqH
Ptg5wGM7Ak9Crw4qvOlyo0dPeVAMZYpG+FGRiL4zvmUAiIR74a/UuSe8hGE+bdudG/53AW4KFv/m
LDY/g0FmqrycAG1FBrX/Vp0nh/NgaCGNxXYB7FTJoENz1JvqeYjOJcy+q3dc4E+Bwq8Ggvf6ZR/P
octTh710G83uHu3IGjLgoyjN4nXtylo+nsRYVpCX6Oep6u3ye40vr+w+kO7WThK04UCAgnDC4R6K
l7pdwWUlPqglqxTM8DbKPe0ceNIpoGGKuuIkLc+KG93Z8I3wUzS9pIJqD+lQnKOBv0fo9A8UgIxP
pF/tXb8SxMBnFYahdVrD3H5t7to/q6QCk1zf51MGGLoG3COQTTi9yQNklI4WTX/FnsaLgDs1JzES
2b+76ODiSxaNalZgcya7Ll1rqWVZRh2ZdtISk4OaLtg4M3ZdrOfi+zDPDgQ7tkU+trhQDrIXji8i
XJ6eb9hglM3ysqfRxKGYgXqssjU3+NyScV744SoPBgfwx15Lku2zVkNNTa5PJ4UFNmizdWYAqJFd
SLOacA20ZldYOVzHSr+JHHKI6Zi+I4od79D+5wg3cqlqj/F/891Y2ngdokZuGFaa5ixV1slY0xAW
APc8pjSp6/KpeRk2x+sAF6aEer4/RoPpcxDt06en/7KciU2JQIQ5QSRy/ZnG+njeRRrQHHWohoJh
rMl6ZkHLjruKJ4ZF2j5lUOiVl9R+fHND7H7S5RaNgG/TyohcipNExv89OMmoh3+wUBU7mvwktW9w
ct/9BLrFl7QmayLNuW27b0o/75RTFaz4MJcI36uod+BotKFPkfcHWWG8xs5tdBP6OdxDAIO6nDNY
Y22winUxQH4Mbp0oLP+XEoKufmk3IVD3ayuGJubOKQimR8Hvrlv4fiyta/Wy+1WA+P4R2vpdyMI2
HSgIWDxj9bogIkY+M75lEzaayMwoV3Z0sFdwisnGSGfgid0wgIXOfG/nCY592YCkxTidaiDhKLSz
dY7HK2CYzXK9kWPu478amRIlkKG/E789SjvuQ0nt6/XUEeMHGy53hC4Ab9oy2cNa154WX5AF5tre
aBt17XYTAWLs4m9fiQ9YJuKd5McRTfBFa9RIzbmzaxa6IH+hvcB/5HwLTf3ACDy8kYOk4ecgJQav
J7tLbRXOtrUliw0e2NCGobquAAapx0W6jed8D6SE/AJtOdLPsblM3RMsbBtP+csnR384bxlykD8Q
ueaj93z0Nw86YSE0WF0R3BSFoknYH73Rd92NhsdN5D27JdURi7dciePxCdiKcYr3fv/bw/UFu53e
WCUkfMBelTirAlr57Z2onxkmc2SERmyfVnfkCGRujniKGrCabx19H0Gve2L0f60ARwUvgMabX8js
EioRjDbZtaW8uZEWp3/FUTuBVxjNlc8JuOuN4fKLgpTbzOqS8s0L+ZSgv3qGKSLi7aXjmFLN89t0
5UUNzGmUlA2SHxeoK9Ur2wva+nxMdh9hMgVUQDMer8SZlcie8vY1hRKTVBilkkT8eVGhMKAcRoEU
g+mOBAnTsZtiwMPLZALV3M4Bj7ofCjFqCPgvw10gpam9AHmigAx2O0T8qQ418VjtLpM4H2gXxPkz
51Y8C5VU98BKtQoRjpKMeebavnqh8awikw6B1kIy9poFIjHdMaslPnSZ9cuibk+6nza0PuyHXaAS
Ndrq4FB8Fwy1ImZ+Y/FcQBorR2uhlfSJkzQdSCWUioA4xBL9R8Va2sc7VMYqw07VKbAnDt3b6Hro
uhLcUNZcW1qJhAloUSCFdJqiLc/JlcAhKnq78G4QBzz0sb2p8WXJPK5xrKCSnfnzT6bpXWKWVhQ7
cOs9uKc8xjbf9ul/nxssnk4ZEEtF/CXSg7vHiZYsWk2F9od7uEFSl+igHSF4RPgLNqTwYlx1ex0R
WYe49S2LiFCPP2Tl+SddcGhWPZHBUEOOX2fPFxe2UgTnXlW8EsdvLv1PkzMW99FwszHOWdG9LSd4
tsSLnGwW0qWYF3lcwOxiczkGs/0TF/UMbglBQq97LIJFbb7p0eEbNKzX35AVktYhvveZael9awYP
qLfkVzLA/mCvbS9XXZ/ORNRanOlA6MjD4YZ+RKYSPPd4m+Y4XAm5yqpJW2/aRfHlEe6q2aDiGQ/7
BH+bruKoSCNi2AbTZNpH3eVvIqUw4186cIf8ErOy07fGibf9PjRBIiQLz1ttw6QqOAU0fGaw97+C
C3/P5YPYhHReMzXKmUe5GhkgEptR3mosUH92EXpaBl2EWkmAlcrVlCVNm0hEOi+dvP8rPUXPDz+a
njJjJ1+vXts8+Q3vt1rfkq4o34tNO1sbjVPyOteFs4LsqUqDUAT1NxoHCMivWd6fiewvvU98QReD
4Aaq4VlXJa6eWNEfdmqnzP6Ckfl/BSGhYDRiatCTw/Q0CdgINzNSKFdwvQeZEWvQ+vDPZzpLnaQE
pBgyGZ/6O31UuJn16kZ6UD7eQ4Id5ZxxGk87lfnCkibJkMyQkIysPf2LuusHJntxhdkX0rKRa2so
NAuiP4MS/MsmI5TuGZ3UkUB+2mw6ewR/6n1pywgz1hcF6khE2jM3yyU7QXKIMGLmTk+SS8wjGwER
N7hZiYjy+EamLLUmNywZlwOnVgeY8PQSFN0GKHYbwVS0LTP/Z0+ZxmatvQYXkS9YKgLCz2jJM85p
QcawKaqFMB9YsC6Uwlh3mKpcrEH7wCwTBDKMabubaKPjQa1mLtrdpyWp1qQ0nykDLfOlkMRp73/3
BuWkek7HQiXa1uRBjdao6jtnKpfI8g7FaoskPLhQ9JsRpFuzb/L6RCX87Oy8Gt2ppXbOngtvRvlP
cXKrCOLc40TZekrxun2WaSU+7tOvyiULaIpFqXQjzQ2GgEngGtTypaQ4+T6UI/8bDPhZ5oHWLTBh
TTOhEWdv+ysjro8Ck8xIkRZzlOmfrj+GFS6htJdGDSMNErooCdP2eMoVHTde7gx8o5oJ0Mjm0PqD
FSqhpeewaUOiS6mUhLs5Jfy1CsjYEjsFfExxPP7UUJePhqPtfdCEW5DlaWKQ0pRIeNZFisDBXjXW
f6GViGu8i3N+FsCsfu9OFv/5HYXcHoVKz0JcBS78ZiE67Kvsou+D9z3ydMLciKDVUeGspaFRWGMh
0Xy56/ce+GwsXFbw0mpiVb3GBQtNTBS2fQW9SwsANd//2GzCN+dwgXnCsorT/FY5GkA7uW8hm9Af
helf5Ot8IUjCpzM3MPnn0jAIpibn3c8eRVnT5Gn2rC7Y5X1KFSfRCp1vYVYX3d9t9N5n5pb8ONA6
GxlmPHR+b6lGFA+tgTiXnPFEIFzUjjuMVvVma/Z77GL8wZjoBZcoBtVyWzoVBfYo+5tt/x/zY/lJ
n+qXxaziq/Tq8U5tG7g+JTaHxyhchbhfxGPj7En1rRKmuo4NJB4SOjUup60sBI6ymGK3Bn+GPNTy
27ynpWeujzLSi2ujOPrI+6rSRSHpkW3qxmnCXcB/T5HqdlVl0jl0jMfrmdQJfnp9Brd4DRNRasPU
tsvrTOb4saN6vVImdITLnhgbWvE8NGWrSuTCBhFtKZjiuQ4vJv35A0+Z2oyl2nN5wnOwZPLmOjiQ
r6Qr4xHVNyJcz/ATJJS8EFxf1bdXUoYzFClSDRDj9Y/I6M26AN3XNgO52BgS143JscABzPMIzgZO
xu6pgo5coSMGep/8/bhByw79iW9zrLOswAjqxOd4k+zxzuLAv5HDnoj5enTIZTdZfMJl9vr7YOvA
rh4jyaumOjniGUsx24b6ygEa4jKPaEiB6yHXRSd032hVyUqNHD11O77gmhbtGA6SaDitedN69lLI
ICgKX9g224XGetZccW5xdkxKbL9fvViMiAr8APnTKLiJRi/pX201q7juokLS0nqXDrcgitZBNa3L
9wcCGfRU+UiLnigVMumN2DzlCbNeLnntkYqGBfj0dsJHAhd9KBibyeEvaTEKrH1CwBgEXpFgKRH5
JqMznizZajihm/po5ONkG9D8CRnB7eDjdGBH9BnjiT6sA3+GhQsCix74yJ/NGGiQzMvVIJ78LvMn
CNmAZ1GMYBjLrp/WUeHX2I98k21w2K/b7pgUu2jhAoROiw7kCBIcAIsQ5MkD3vgY+QGbc1wKmHi6
q7ygqB9zIral+G3+13x+3lHoxjf3Elou/XhL/YI0QL+JemvDKGh+UGgPRGA+Ep4EYXE2hihfWadF
p/zME8cPoYugSJIeRqfxSeNNUMNzZ/64Q+M9iujBC2PISSTDLxkqwTrwOL7qOwxsdVQzPv5mhwXv
PKSIToir4oPui88i6PjfqQdtEKX/YtBy7/I3EfH4Q/1Cor6T1HFPmA+hUoEikrq80IMLw5glDcY5
y8C4r6EWmMcH2UXnh06VAK7cCf4Vt6jL8BnIOibDPhwis+R7BqboJAP5kjRs+G/Xo6rOnXMUVMgn
6VUdrg7lsFaeVFyRWShLBgc/NReWSHULoP9Y4Stb9PXzBRNwryZqKmM6fMTZT3iivI/xvBTMAGgK
lxKiBmJdFgIKdXLx4EtBNbIDgJHKi1jJclKASGQbdE7lQ7zyVu4wnCSveDLDFcjn09q/1qslN8zr
WEBoriGn0K0dOSrrLLUF9w8DQEaI2JpF48K2zWw+sc5KIMkwHge85qY9Z1IlhM/scO6asz5j1K7w
7LdnUDcoUKVL2DdwIv+YrlF/VjgtPhPhr1n2lCwXjtnRMu7ziskoEbkJMLzRARN1L8jjF7skfhes
j26CJBFXG8yH7uDDmukqTTFxooSM8Ahoj/rmxENx4dbDZBIRvF7xMIXh4lacLlkWlkknm82j/gM0
cANxIk53j4mKKwfSE6xzpYzm9CTQgdnmdlhazXwKpNAySSd1bwO+uQs7p/gdQ34AgNAMllXKg692
F7vmPwAYY7rDqtc9vzlyYKDCZXMjKB725UokZN1BbF/Q198f8gYCftI4wBwKyUqFZSdDneEQNguW
Fsh+1HcAryaFjeW2hiHKpJOSdTDqDU0KMyn4UXBegCmUvvxsKEPhjOuZxBwVghVKQPLbpbP72hHV
MIsl6cARdg+1goKlbZXmG6ioDueTbUiMCVfbYCvhAjUSjDaRQsna4OK3OnW6rruUw01RJzbbp9Hu
HcYBdWg1FQNKp/yb8sRUeIK2DI8ZgXv0zNLRiQV1rXVAe2aL4xtP+aTsdDAn8A1iwpy6+ZhcBb8a
r1OXvCrqeziqVvXsCu5Ema+1TjZKI4AZqTkWMx4EjkinDZLfDJP2COXEnZlIEiYzIGEiTaNa4C86
bGXMA4QRvjhcXILi1IBoixfxn3Yl9S24p/siAjprNTxcs2rUDGb3/MkdvyY9JmdQ/K4QI9uKlYNh
0cXGu6y8wDg1SOoljfa8VdzZv/D3GqOIK6SYP+lRbIlendsBVYSfE1eWAlpWqOMxtWyv9m0Ngifk
UbVHQYUqjvWettmf8i3gmJ+0X5nz7xQDqXeTObqcVC94PW6LM8KI1KjabgHeOX5BsTaKk0cnX41F
s5Xwma/mrYoH+0Wf0zgxHhM31Hm0B8sISCoZIHgHtbN1DQR60va7b7n7THXqU8TB6PZTHl14X5Xt
Cgtyym01aYfxUClP11SGR6uUBB2WXMBHvyi3lSZCfnOMjTCce9IaD4I4ObWrn6Ohy0TBHM2kBqBw
hJ5cUlrOBTAREsa5kI9CbaamOteu+6te5oaPV2WOFxuAx23CwFlMJFYMz/kwYPq7uyp53iVzL49l
62O9YiNF6T12LIYF8oBCwwcwfRjEysKPhICuTeY4I7OBlPo4mY/A17qoK1qj9R5odHIBFsnPdpa6
Jidgbqrzful/T0T4M/kqqjV63PLrjHPuuiCaJuZryCHPt4DbrNvO2ofHOc+Qb7hHOL+2utZS7c54
WIAYG2gvFIN0iuWj6Oyb2y/7O05I8/DflrrUo8iWob8qCraE29Pp9862T6Afpy48nlniAJQ+WMDo
4XbHOFQa8M9F8i/dYnoFju9NdH3n+or/TK3iQ2DCLK82GYVkD7epTezsaX5KK1mocyRgiMnqH7jM
+11tzoTDWSGgzJW1XfeEBu3YPOY3jpKei9FYYeiXWWuqBUEj4IHX8LH0xpSnxxmCNmFqU3WWhZ7O
wmLrcVOMDMISXL7Rnvv/xJnAh1TH6OvL0/5ziyshq0165HCTtyis+eKV0ulcceNseMgtdmTI5r9S
i5ODvspGL6J7gDhTOUHXPqY/D2D04rOWIHiM45PURw2xVTRYTyfRjHp7JCcswSppGfM1WCgiIBZV
0vTQAeFLXQRpEtT42Y/QJCRZmf/VvK8GvcJzsf4KdlWcdXJQ3RJyFDf6p4yn1mlXp3rApR/2Q1Sk
f9tlpkWGRslX45eDJwil/ZtxD5Cfn26NKPveLpMwgOM35Bichv7kSVVLIKuWuGa6JWGyH/KcEf+3
4ufVqMRfOi0jZf6SWB+2R5UZ1lepjbEXwODxpYuBM0vRrFMjLcrarhEjv8x9ZAHk9GDIt8ENXuSD
9azBTQqjr11ANMnSmVfQUcabJGMjEImAMvZbUq+Gk1DKHSHNuXIq3NAYzMbx7U3ElWfAjlkR/fEy
uQcB3vYgjkgv2rnN/PI45xEL/o2Zibmqbm5staC1PTT2gcA2vDhvvtwks1ps9k53vPD4nW8+9ac7
osyovFqnj96990UXOE8VUngUPXB7h8Pdr6T90fxz6QDJAKeX4iLMhsTrD2lNCZdvO10bSj16R6sv
kP9uJa/myv3baoCr/pAgOoz7o6glakO48uwTuJXcN78z1R2MM4LnTQZYPSiZmY3tlqznmQFQVJkC
txKdPB7PV/gfVSRZT/bL8p25UJY2QTsajBB81zZzVq0LlDUd2CMUN9TKn+KmDputYLcJBVrxfzb7
J3hXNip7wXEskPDwIj0EmprVoKYFy2rHDRKl1Q+4nk0gtol8TK2bg06IjYILkyt2C5801nTAZ9HJ
NQpSZcDtpzG66YFN29KhvdvcGzYoVPdfHQ97HLnk11rRodAYvvDQQL8w3tqEX4FTxevuwQ//JybL
Ytq4RzcxF+cxxCHqhAx3CNW4AclUYwH93DeJ3GIgpvjEYYi9n6hTYt1p8KtWqRN4sKLt6cN8ONlu
LDPZlkp/36TrnttfG570/kF3VkKO+TgXv2YECIZd9dBYxAsGYqKf8dYWkWGLXCeHu8TLEClcEmq2
EfWRwUN/5gEtfiXYZCU7MEzUburuWbEb//KcQRHlL/ylsTdfXWoaOG9RJCfzbZUFnoH93WKV/sOU
yeotsaO5G5gS2C5yIA/j24MCJ8PQYIqYny4U8t5QkwaYBgXaAnawrha7kKwZ9nrtZOrzFhNNn57u
SA9IzsnzwEwpgVkZEYyqkfq8DOvMpfmJZCbv19430ZOhIeH58tF0RTgWent4biqaRItA9o1jSxuZ
Hq6vDchaFih+IjQJk0T4vX/S1DA557Qq8OFRK5+0fzKYFVD2GAZ5Pn/44FJkUD5BlZtLvuywWZjM
E3vO63Y6Q8my75EtkHxJOFtlQ/sKaMCZ8S9x7xDfolwAf8N1yHuXLh/2+RbHEBJs6WF6lmt0hAYH
LnMmtrb6EwQuL9ski1f5rveJmmLt3f6iPxXoAV1wflkwI/vfjyUFCVa0vEKomzeRqjmTMDcy1XpY
Oqr4ld7pigmpUkGFvrS1FhOJB45Ub3oNXFeK+MLtGeEWatIMW1zD4hggNLYi/hg7qnnCrPUT5M9/
qjEoUqE7OhApe8WDka4lJb0NrxVzq1KUDECRY+0PEwei81QWyIuzyNHRmpp8XzvlwGpSj4y9arQp
5R0LjuPYWLGv66fvajFuRotmCJ6MqP4gEb/7LQuee4wx/VagD44Wh/OBGVAQHCDN7TuxZY+BN8BP
WF9hls6ucvIqNBrA4zm03Wj3e+jbi+EO29epYS3mA51BXIo+x1PwuAZiKwEGISBMi/Cj3NFj0dju
oXzc+ILr8w21/AoUlrFf7bXkC5rCyRK18wwx/g42VaHMdfvtSItNlLDxVHQ9VCx4YGsExVUYt35T
wS0lkRArI31XOX7rlq1CqfoDUa3/6A0FRNOieS1XoLoIuQNCJ+qKj8SFa8jbIsej/t0YFI66Lix7
pux1d47ksvHvG79LfBCrWSi06kyMha7BBiBY0WHyaQnzlt7+MMeM0frsiYPuoSePssQ70O6R5Oks
fGje3wcNCvz+QAmuHizyDA8Ee7df8r0ZGDe2T9lxI9QduytDIZwjsGhUE2SL8qmelyQsV7RY5j1E
eKP+u1b3aRGYTP8Vgd2LHahRawn3PBC7QmF6MtQGc0fqQkufCj0KTAJYCuraG7nFyvrtDUGbYH0w
H/KoVwcl86J6gvY+nP0XnNkisj0zKjPLqBmfcqzM+jN5euyRq1pBY13gCNrYy8uifnJY0f7KGJ8A
0xp1aKoNUedLlDwmqnpTDM94u+mK57HvZJ/jX3f/lKChhhcOBuPqXbgVFSzpF1XIe3gl5g2/G8DO
qjcr04N9YiESIEKD96oFfjEIKphlmHPFWQZMEVgWmhzTshCqkSk1QpdwxcLBV1F4SOS+Y7NeAEh1
7KnUUK9U/WuVZndnzTDHFAkmXqNQBMpB+N1K3YB4F45JgRAFKN+IFN1FecQRhVX8EPQNZsLNucFR
Zs8Z+61fe49p7UReguwl4M3smUdd10yMdm9Y7ILh6Pp+e0UJm+9SceKOPBXTtvLWlBryGt/WII4R
yXSqJFcr5hd/HJ9fylOh9p0dD8ZDkV1rT+nu4/Nv0IjNfNCOdfNwhSUEApI1OcZNHDweuWdQFTKR
1wH5NCuz2TfO7UrONOgcgureyLCdd5dcVE8fa8GonO/E/As8lwcFcUQ1f22DNSgKa1Jvir6NxIaR
Vf07Vr4GVpi17h3GniOWrKSouk36cvs8gihoQalfgxMJkAQVAZVQMWxTyWE9irx8iy4YelzkP38j
jGH80KJGPuleF/J7xcOZ45ehHWhAPUrNPt/qlkfCRC13v4hDc4eKotTbz0o+/Upddh0KvmdzJETn
hG9Y4LWf89iS1haH5GGbfJ8OvvaCQOuNAJBfOz6dRKgoDM21GZlOlTTTDzdzSMmg5LbXO+HTlZ6r
/SLxZ8s64688FLGjeg5V/RoRDcck3iGF3AWQG4XcKHltI1eohJXtiEPb6XpPI41JIgjxkxfbub/J
Xm6od6Ex7bLbu4fPCYgdWLAi7RkPq9BwSMCdDLrItMZcJyTXRRS3VA49TBxGviQ5ptsEFd+Pe1PY
FTISqmDR2ugsx62S3g7xB5DVUbyua/k4Ua1WyPeZ8h3xmqBeV7315cKNBqYWjhDfDyG+lYsTGtJY
HtAN7n07E3XGOkIbZ2KtcipBPcBl7yWdm/hpa7BN3GiRc9Nyw89hPggccHid9mDm5KI/R57+eq1h
6/xvAeqSRbegmUHn6e5rsnR5nSfBSb9cuC8VjMbU4muyt5GkvhX3Ly+EJ/nZwTKWROtugGk52hl9
YPvIZAI0f5CRcu/BT6I4GxhaMkRehUbTWH3j3vi4oUupmE28w0bbt8tsDTMx+GQ7jeD4+bZLI0qr
JWeMJNOg6yIYk9y/bsDgtb0cab7qbfVbS3EoR8k85zoEkccvaD5wlwv0WKkQViVpBXNWbT03h+Cc
6UJR0JBVgM70HZbhIoCH2dm4n21kQSd5bVPmuQUYVj5jPBXoSW5z0D71OIfeMNepQiLePzrnqqeI
05jPTXCSlazjHvgW7jDH0qSt82PM5yUUU4Np0Pr824PL6Cf/UkULhTelEjKwzOd+ZMYBmiM+K5un
jCPKmOdozQ/NEbb9Qc9KF9trO6NLXEXxO/Z4csCMOmGEJB5pAkM8ttWqivuTFCZbxnwpQailNUVp
WMv8ay7PG3PNV8/3kcFD+CXeE8Q+hUyYSxg/AmByPpSVZWJvoRZEVmNG5KFVzjuppS6SUr7z/jQw
iBR/1toWC4THHXhkQul9qHZIP52yVZ+bmVaMwYGrzqa3Cd+3AlbcVnBdxj/t0Hed2WC2btuMiNtm
gX/jq6FhnFi1dB+XKlfLF/auUFNaK07whMv3iC3zuwbbWoYOc+7UFZuYIDE3NEZo2KTmUe+AKFYJ
LH3RJOTgQjkKAZHTiSuOB3kDeT4KqTafNbcZ8d+ZcSX6kYs3DHE1Ccr0gsgZxlzEwWc52poxg1gF
AIXMSiSnf9Bd3Z6WKDEClSS5KSg0SlA9wDAlv3r620tS/fdHzRXV0JUXw+eIRQN+e2yrx1DzG7w8
SHHzJJw8UZ6zL3S6bQ6poQylzyqW2wVaLE5jAEd0BHTn6LuHA7TlKsBi8G4YIl0qYw2pmmtYA50u
gf2yHAXSXEe+qPxDoBProo7POrynWeXoI5k6mjlmT9mlfVLQ30jNjkQFBiEnTRwH5yry3NS0brEE
wLafJarO5lsAAV6dbdC/c3S02sS0m2NG+/ZRrFokk8RUOggYr/nwX/3wD7u/UVOQrVC/KxhUrje3
FQ162TjXnIYUdEj/0dt8znPh/LIovwdsNgpvxK/sOK9c+f6gbALmmiS/vbGkla7gfU5U697XYRPu
1BV2TNTjzDQLezRbd2HTNXuDIFMSIhtPY00sFieAVcvdrrmM6Wns7u2EiXi4JNU4XyLFgBkFr33i
BYTnD96PZe0apjH9/bTFfuO7JAFjOurbvFzFQK5XO09OxyyCGibATFl9+Y5hfs+irU/HSNc9Z1d4
rJ52IwMEty8A7T4GLfDG60uVWZJLScGymssrIxxYzG1a/9V9fg2GgsnekwoJhd91TDpHkif6vhbQ
TbJrCEwBd5o+KNbjC5rSFPsaCrr3ApQ5vx9ODCDfcfA27cLfx3SD0my7SFUqkB9GpbtV+RWtYf5P
YGpkhwmNlCJ3H8j5IjMV/Qq6Y4a0ApXIzpenLJd1PebH73yzZ61PaGsig9XgeX71s+x5gwJdhpTN
3hmNm/cRMO9KfcBrMcnjYSOirC0obRopf9xmSQsfrTtm/wPZqXWtPUh8K/L/yDdnoGfHAOPmIb7v
/1cLTdaNP+t/S4kCcmr4BhSeE1vVVbR0vp0UF+iZGyyE2ymIEuC7M4KnIOMvQLhe/RZjlTz4Vuz7
VScfaGO9TQWozVyHYbxMbuM4P5YSETFE4zTuqY/WGOFagxkZ881rji1pOPQ8CqDgZeOAgojMMIuP
7M17CRPH2/yrPfi7Lx6URNFNLOhjYdkyCY8IQEQa9Dccdx23cbbJdhLLHJKLr1pDsKybkqSxNt27
I1pzJwopjfkqcuWeFIFymOoIwxyMC9/3WjhZrWs9HCHIOm/x26C95XrcPt9GC09Eo0PjBeSUlDub
s5guT+agWofwcoWEVqkqMW6QYAGBVvfl9CR5Arh4VJOQ332FnGnIXVb0tYNp57J2ko582GEZIQzx
h/xsNLmqiOdZwk2NV0Z+ceF8O2FdMVReVdVlTsPghaFKvAhGa5134a+C2J/zVly5yR3jyF0ss8lJ
7NWRikx70GmqVpLb0tb4yqze1f7pxnw6PU/0vOjBznJ0XD9WNed70/Vt0Pg3Thb32CIxec+KccH0
d8ShdDiPK/Ltkgkk4DrcdhV9vb/9FKBHbGMh2z5cv773H6kpMytKBp3syT8CbGL5JUlcUGWitIKj
G4a7AruD9VH39JbnDZ7dTjnoYaDp1HGpCuboqXgLTMEt3A19vHMvN6KtTN3+21fglD5VHe2D3nyY
KUgu5yJ1pkT2Yb+SHN+HmD3i8kgtgGSDkQY8wBHhN3qOhbTkTzezqbsrvm5rQ3kMmZmUjtFeBIn0
LhdxM/8QDMhTRR/1OQO2MkScwevBnoFpat0owUWJVlBMNLnx7lobJBoQeu6G9nu1OOZ5DJ5BoAJB
gk9OR/gQPxJJSZoWGmp+LAWQSvO1+KcmR9PLPr/GgUg/iacVYPY3C/TvrwhKfDhysU6Z5rMGXTTy
zVqYMa6SC0cNyV9z1WD1dkgl9klgU/zNovg9NOdsPBAqKyGYDNS188S4YNZ97gjwQ/ZUsYhEeRUj
JNqgIC7Q94V70X7CaOW2unPUAo32B2cmZm7fNk1+zC16rLylgiaTcYJ9wZiUEacXS2ukU7/JXTqK
N0pF+ovxXwFrlI9PWA0w/icX8yeWE62uGp6S6iV5xQPM0WkKTkv7A5Q7U1PCrM8oyDrVRaw5lR/V
x0rLsp6IznrV83wOf1oulfPoQKbb7LhtR7xQDWuh6etupqwirHly02nW70RRD4mblzuyxEJ+xtTB
1c0T+5aXg38mwfbHCtfkpeDj54whh3gXahCdZEGyHo257Kg4vFF1w1hkvuRdBgtmVJXu73DhcLrw
PeZk8jB1BI0AAKiSaTNAe9NWfN3ZHw7ARmj4LZtBSkFcIP2uogBHjflzPRDqJZ0NzjV+dE6b16kk
a2G8Q+JZL5CgCLqpNDFyDvMM88Jp7fuB0rk2pLom4nhtLEq5IZo5UG5BaCjBaZ84HkpRlB/LarJB
MbtoN4viPPwzIcTLlRtw5qpcyywm0g14Ld8YfxRVQefEDOjNajxqshHZME61/vBJED6NyZT4AHU9
FI03PEgP4zAzyEMPy8upd+nHBBYRmftESNCQLzqdAdJBQGU0Zli0bqspARy7uCeo7rv0ncUSWQku
6/kg+rOFCIYex8sjLb7xKaBrxaID0smRQ0kYaYT1xvYTV58WT+CRlMBy3i91i+n5REqvlO1+SUeA
ooP1HTucFqk+TxamYOM62JE7u0eJK67/DvMHiCZ/TA8+5m77i1xrEEEuM4mlzFOnhxE4YkTniSKN
Ilu4vVKxKZ2SS9u6oEXP3XWU5gXKH0Ap2r7JKG2kXtzT+Gc8mJ2zCPve6YSSwoXkCoBnVo+qmnx3
HvGEXtY0Vim4wP5luebe31LCa4xrPu52qfTGNPxDlQLxkumFUhJl2tC+7vT0xNu0yjMuf4fV8hhy
c4gmM0guAWZhR5HOVVtRvQOPW98MW6fclfqR9btzvVcTDD+jqoJNU9/41ss7eFWZZ+foia8k8afX
8frjhiTWuzYpY1OihApgAmU+awmUawSXQaHed3DQpEGoP08b2zldM+sRBwQNxhsl2akEh9bXo3qJ
Dm9tpQgHVwvshTy1t1GVqfnOQbpN2DGHp7znRlWspuzzo+oXQd2PmFnKnwiGgGUppWXIDOuPYFGH
+/EMDQkdcbc6Q7Z5napC90gmo+UzKLBBUC+AiltdF4iZOFxgx/TyElLEA0JqRXxLrr/wF8Ic8994
2D7WC7wqwNnrYJk7SlkFu7okysO3CoUPr/tgpAbiva9T2Ic4opH+oIyz1sgxUy3kPAZTKWO5bIRI
VxK3A009NFaz2LqXQYNOg2DWHPL80fRP3l091GTFp247sap9nBOfNUWhyoNUpfl9lgqcpiVUBU4B
nOet0Fyf+gkR1Hf47NKXgFnmyUTyk40J9J0S1TIbK/syGj9FuprrotLQu1H8HmRmP/SfO+S8sRvq
/whtBcodgHRNC/wQnr1hHeNvOVCS9cN5k4TWkeuqxGzJ2p1Ha77sxu8Tb0FjfCTP01a1tz8I3LEP
GBMzsqkqo7JT1cR7c88x9PhpfhxCNzz0kymez72ezyOFSORkJ+h2dUWOeS7Lk568VCLrNwjeO3u2
00i4QZwJntkAOKMOEHFLb+zQwNcQcs41WH3SZ9FQqZzaJMcEsiCKrymu9PNMtsRYsZ/hsz72CenX
WdWk4Sd+7m+daIuZT/zOY+QE5VgRS4DjRrJG9wyH7tm1uUFDV3/87oKGO1346GNidNS3H64kjGOA
LzA0r6PYAsneg1Q+rPIlQnOD5tWXg3W5pfVX1/hKmwHywQPO79WZtWf5td09JdGdC7JqKfzduR4h
QwIx5opA6i0yHmDd35Pbjf7QYDizGXDnp8RFS8Dlqyfh6GXwJaSuMmuIxVeNL6DNJ45CAXgAl3su
Tyvo+Ap6NyS8Kbe7UXxdAY/hMw0JQMprHt7tB48rKErwOwzYYkV9qh4CD1Z5049DvoRxhSZ4UoAJ
1J9H3Q4dTTMehxNu66pYMuaCxSpcTLJlGM5qCx6H1n6n7qwbNtTekUvhmTlL+nUFbByflyIME7Ow
iG77o/SBUchLpByPpsFuwKZAojKyhxai7s+ZbH2Fmj59EH3vHmWAGV0pdN/TIGgpwyAIGLu7/BsL
TGr+PdNFZCsfOLg1U66zCs6YDpckPtkzp92wuFPAKJgzxusE4Mjvn3a8tgJtmf/LV3P+PS5SUn+t
PU+QDL9O2NT/4HkpyL9EqPDojA2XOaJRQ94eIP1N86IjkDwjm4RwUxkVTlcRepUViswSwcPno+3f
1xzc9v066+fNqA+YAGFjKCLMUc7Dl/qYdbMmWpQ+aFpISeNwdzptS/Tn2cDV6aZ4ed7qXev7irFQ
H53y7fFNOFbqi2eIeNYFRE1OA2JVxrT0tE2wA59/NvcSyXuaNrK81TlqX/il2NJ3j07Am6xac7xq
od7VKODWnMwpwejgQ75NO438VQJ3X0Vz6w5Fz/f2bxMFx+9RdK73PZHR104c95OHC7gnhKcevftP
MOPsiK7MZi2q5vRVVOE1uxwcOsh6M4FoL59gHIMr9YOEWDW1eiuJufrJft90vJEtOjPD9giSB8E0
YlP+jWPPqz0FBC7lEAII7vlFxv8hogcqbeGvXJCbqjo+j3tAYy/osT3mZrXJPX+wFkwmuwDuNVJi
i1Q2q/lG0yQ7q7PKK2f2nH2rQgtuMUMJSXD0WCOLKSQZ4frJQdEMgy1vWtEEe7bkaGPkcG31eSQm
SZZE7OUHQx2Z4EMIBTkAgKWaf/ULXZGGD86RduVHnhjaR9OdE67GeNodwCw2K6iGXi9c/vJ1naEO
eFgURYCq5AodNCvJrQg5/Lzeuy3VCKIG7O6ZtD7isn2sZaw0GMFO+ilG9rg8BOfW3tYH/0A2BPBV
j31Xul3wccEy28ATSnlcoIQ0eGnKCdBIPqcc6gsixmK+ceF0IPU29UmS1NiURRDFVfOierghlBU/
sTQJpmFCtxtooeF+ax1sef5b1kroK/z0AEdRwP6cYZf7/lkBSEDcRa9UQZdWwjPVG5sJF1JyMyNQ
/JFZOoV5PSyigIXjzTjZK+ECcCpD1f8LAi/+Hn40KFSxNDNh/86hrHp2c2NdT7rsbUqRY+2BZQ7H
X0U5hz558YWQkIgVIEkVidR5PV7uwJx0EZfibtfyzmJHcovcZ0EZpM278aI54TLxKphxZpdUQXFK
ngFlx9jEa9WJhk5HgzBdmGdM6KjfbYesbMSQKO3yCbvEFLRwV6tr9aL9pgVLI0gs4W9pjUId3gJS
W1yopuv97KtRh3+P/o5b3KwF+1EHdx9mB9YckHHbRW7KByCDVsaHdPf0La8ifYhj0NkyMp6WjXnp
T8gLd9xyMfn4YoYrx2nG6Drqoqj6j2srV1k9Xw8voOb7JZwRM+AmkhuLaO0IJlFpNaKvuhAuok0v
bBPFZY8H30vAvO9V6us2eUEp0+RMBSDF2L5cHDWDs0Mdo34Emz1gMc3GmsvUQzMLEnU6TZHZPlC5
KtL46105xwJ/YFYWd1uS8/D7K0kCB10PEU68/JIdXCaBTRzLufxlEbpTsJAV4xBoa2pKWdXzH8DF
so+MldqAcir91tO8953uy3onWwm+3abbVevJ7LuJbhcIaCBTKvvoBpXKUasEnCeyXSeKOgBmjuaA
02QUh2qPnA4uoopAGQyyI7LpKj4qOh33jXKqPMM4QBjfkbh5vCnMaxEQYcPez9hdq0QDR0DwCLwb
wQdWob0BYBu1YoS0gS1HtFMNgmtaV2lvC062UgikHHLivuLvnegrBuPSXcZul5umYKmx/yLmoS1v
tooU6ZN2i/ELMKkwWttLB/UeBTgfpuconDLAYQOstTw5C7DHq4LrLX3F2REvVuZkB93Ed/Yo5/Rb
tl9utqrr1Kl/XNqBCRihsuZezc1gRJsU9kV8ZxVuZemdhMZU/H+z28oS3bWCnixqGzhJaDQh4abQ
2ChYIMUbWp9Yi0OnM33dIJRRTzWhFwU+EOt23l3MrAEL/ezCtE5OlVuvaWTfVBPQLt2Gs9GqLcZc
t+QO0rWL718f9hvfKifHKc4K0T/zyNvNaCCJixmPGGECtxsFfMBamxwJT2hJ3sYpnOjcDcCFogil
6vnXdrMj94GghGkzAi4CdCr5p22VeE/jutUccSjpzWmCT2avYsRQm3JTuFeZoLdtRvwDNvL/2lGM
hNSkzoLv0IV7lL8Wpk/MTuZ7gPRlMZjxCtor6Rh+H1G9643ej1AKQK2e7eqag2XHPssnYfneDto5
cP+3r8uAOaYCFoPdcKjKObPkhHDxUGkbpOSEHj2Ag4abN9Hz/Tpf2iiT7VbyG/0jjtP5yaZSfbiB
uzDuG9093ZuKaDXL/nsEDkyD0wEyjj3QGt7dnqxBMj70ngj9MUhWA4U5YltBHQ7HnORYeazo3XzU
zMir/93P5I8zRN9tvcMT7plXO9i8v0Lraly2KyQQMk3rfpPrjcJeo5BzR4SFAl9WaPwjaezypqcM
QF5w5nmJAJe5E9Ortpv0uyro2/5GL7hzlwcNDQl4ByiaSq1VWjirPT5n1nsxyqAjVsAiibriE3T8
PMFD57XAIZW8NLiTyIsLk/5uAs9Izwmy5t981be6YAdNwNqXHElYT/WMO8zO3ud1lRJrQ1OG5JQ6
7h7TN+JGm4EFVPNpukcbBrzvWfHgAidqqnIFIHPYerP6NmGkDA2A4FHrFYcqa01r8GUk2Et1QLPe
IRHWWQmV+FICoLD0/+NIdV1I++YkBfOc2r/vWqZBWxs872WOhPerGZOcIsatoy6UY19mH13YFwqT
06WffhI6Hv92UlS0QA+bDFgYKPMq1bPUy62hkjdca2W3++426rXcMbUMzsRNJV7ssUQiLpCimyro
eLmT+LKdohjjGj32baqN54R6lxKIUmNCtSQsWVJIywu994G/DkhbqIrCVkdo2jcGmf9wu/COMGxH
uYRSNpYN0Tbv9OsKXJgevUOtdYKtPnDdcQcb75hyo3abnBO2U9T3FzDJilhPAe1ehV4drxLDNpz+
S/fEa6XyNuTyxhGv0jt7BTuQqyLxApQ+AiuDxL0NtyWouIHT5JOoGnWa9eXtDtrf731jYmR4tpom
qyqVCzRd+msboZd3NUSDxUbK1cGlreLr3iSaaSvntlOHCXPozBTKXLl8npbHgblJVQPBBzoN+4z6
DbtCDDfb2U9WIjTX4SszfnMhMAhcfbPN9sda/5YEDDzgZo++xwlB3YjC9AeR40rpCI70J5HN60ZB
bYLLOFLxIe62tEsqfxVWGBPIAerTixmFJPqHs2bTzq5iyL3NVf/xRsw21pHTjQrCzPb+sMBDzODz
ISmilFTqumNOipMB3HRyiewILdD1wEwjPafxQCMuoeTldb1Ja1HXIktrMnQropWZfpTT7WxPbaTk
dl4VXMy1Uc54ZSu50M3Tvp/fkaV5I2IFH2HrkZDmq5p6Ycm0SVYsT1fOiRO+TuZfoLIa1hK3pxbE
zAfKo8xc5aq5uDuIDJX4kP7bnBlAgL6Wsmm7Uo9xcG7OKplGrnc1UZjkFsio+T8tAFCe3ZE+TdCI
MNIasvSvSSUQQKghrlI3ZmdyLaQOr1TD9FchNUSF196X4LNfqMgnmtmPA3XBE948F8x04FK9601/
ObTjGmRS6Jy4tCDkZcoDZDZoxvGAmx++yQ2JFw6vK7osSBe8Wnb0HCzoS8j4n/mEDlWfOZ79Wl/u
k4QapXdA/8LcN/iC/J/dYh/Us5Yc7IWSXvdTxVxuDD99lhvZprT2Qe1cpyOnhrLuQVIrCA8srJiV
ckK0L6giLNW/BCr+KOWBu3lyZ26zHS307/79uI+J+sva5GIFwDdBQeGDfCyAFojZeZzS2rUMNZJJ
CoLaDQwjdK8DmAf2m+PDkAR3MMAXrESz3LWZO+VjqBR4rOFHtw519WR+9LKh/VBhY5kTmkiG+fYh
FqkcyEHKP6B4iCEiCU7+8C89qeRcpYmgws4IrACddke7CSYsQnoBc7Ha98jR6qPwSnW5hB7EelbR
uKJmPhcrl4f3w1dk3/gDMI7O56Nqemm9HfawFKMw0tNTlQnzgJOmSfMv5fMFb1ePNGojt3bKatiK
6l6FzIQZMSuUV/CeIpqngy+J/XMQxbephQ4Ogi79fELFeZWi2RvAlkW1N69bPDCavVQ77CvGZbr8
tCYJHQiWG6a1tO/f7huFS1vfDLQVy0QqePhZ8j1vUTUYzXYkbHa1nAMqGMCEYhzmxdCLpQ6hkAMU
/zLtg+BvXVO3Riytf1BQtDZElrdNzousT+29SpjDu2zj0AC+awo9KKhN4eoAtxpjvdOLzgNCTL4G
DGodH07lebC1CaIFTLnu4sdXiQ8EAMBJ4OZ9PWKkS1S3egKdB9oNqaxmaquWerDxgSJKo0nf2x8g
W7s3bkKV4CYSC7a5SPY9/20gZN6JPgQqoBBj+EW6fbIiJi4oxm7j1HsrKojR8/dGwF3JmsLCjB52
0VjfZlQVElHXp0AmU+3C36DORK6d3pj/TP8g5QGpqSGSQqUTAHqD1FOyfXl8W7LDQdpFsF6GlP9W
xKthrIV0dHobSsRtlJzS/czGP5ZX4ypIaCLoOBTvlrJ5sd5tpGJ2pnW+5+So9dwojYUshz8+WWKz
ntkxL7u8WaW4wNkBjKRUhYnkIHO5uAREC0W6aJPB4kj8Js0cjqcgcd9/+wAME3rYJgwV9YOXz+5m
+wdG3cMsZlrgPsCWgOyGNWJ4su3aUqvPsjI9rV65WM+PgnQyvOgyhE080x3qTxUGVwho6nba1awe
BH3Z9ye5cIRJKalWyw318lahGwa6idrMvuljC4xRYyieRVpd5zzpCnS8YyODAtSk28eD9mPgct3m
goJYU9a/ALR+hcruSu89U8v5Wh6053HvAX8Zd9pw7AIAma1TG9DVoKBLK8FqQBfMVBAvsZVOEKif
jZdoAVJ/IEMU3Nkxw3H205/RQDtBoiu9Uqc9WwWSaezKD1FCRf5o40IzdmsYW+ZEoEDIjyyPH7C1
6wARpLDI0fmJcWTQjklREvwDusJyTyTd9dzVql3ZOJsoE6KiqPiifUM9kzKcBtxf0UBA3UDxZRQB
XAp0VfdM3HYehzeVha+EVc8aL7iqvu3MMxGKMmNedgt024YhSGU/jKM7sb9Xa/EzNBSec7Y+G2H3
aZdFWsIXMRDAVLPvhgeffxh5HWFj4U98g0q5DPsA2UFAzKmow7zp27cTEIJrRd3qdT4c/iMvxe9b
C0ubJs93Z96SlGxj7T94HJOjtc1sB1M6FpiJ06qwVGFI9ONX+pi9SGimE/xgrxYGuTE0oLebCkeF
U5213LEirsR6myZaIRWMw5QbxYOOKBqrYkmafvGwp4Qch8uWGo1k+nkYQkDceqrk3D0o1mOeCF7r
0vgr3zsNO7T2+xRHS8pCCMsBDU58ckMAKpTWpcpO2gHSWlXY6b3UrLOakW2bs4HPhHcaCeoWgPEC
N7PcRcWgkt8npOH8P/OUtX86UKCxf1cka9V3TO2WBCD3K8KhJvrMoKZSxN53I4E22jhM+QmxbK8d
FQm5ODf/5ZAmuQv+WeTSKl0UpyYhO0VvkD59YLNkgv0d2ySKg416onmrx9zIP+V3g8ZTB5jVp5vZ
uH7zYEfiY1GWT42QCZfZJ/QYYSube0fmZA2yR/re0FgyqfCXmkZr7EF02oA2/1JqKyl6RrgO24+j
+qt1j+SP0RHfqjrqk0rsaTT/gdiZSoB22cw0MPEWLImCsbS0sXbBg9CFypd/TxuF2ba/GfzDaIi2
xNcoAF434hw8mIXZb8KOhn06qka10hqS0sX8gbOEdp4I9Gj/Ofz3mWJCpKnp4Th0nxHNgUBDmA7h
V2vkz8cZP4HRGD+HKgpadqEcv/yiMG/885abkxl4KObcdw6u5d8yePHiRmqTlD1aFuBAQp4Ubugp
YWzM6dC7GTYauXxfzya+x8GdMpdMItIwlo/drTaeYy5S6wIcwAnyeFfCK+epOAE6/wfPEkSLo0c+
MEVaihbPzw62ZhdR6Tg07aPuGU8y+BvObbGSMdluFhUn07I4Z+grJaMq5bHMXHQOPMr7Mw+VN9fI
PjYZRB7IPGUOwSzz1Ei6eR5xc9zFR//W09SrRxhnNxfXGtWbw/IUaEbTEAHsyNuUok5JkiCni4BU
V1aYIZAiaVcIKHx3velqcnRdPi5YDiBpsEGnK4dCMEA3nejSfLtv8Uh/XIl/tFGPM+owKjxQzbng
99cS+KTbvOPGoFFkkqS2sWHgyOSAYQ+qbocb5yEdGoAo6dW0Avyj7yiE+eWga3eqNZ4uKaq10i0u
ph1LS1KqvmvhUtp9V2daKzgSYly5PnSqzZ3iqMj89eCbWhVof4mvIlT5zRhwlhDEVzpzX1/ZEypl
17YyEYH8b7o/PULCQL8/nc2N2m3mLsxtvhlxn4LeC7k8x1toJg+Y8k4iD6/S0SVm0O816J/9Ent4
6gskbpFOWb9suwo74/KpQZCkgiVOR0kI9IBFBZ20jy+uz/q6zRxID9tAAix2FYWbhOizC0GACxaF
URRUtbriMwJwEgiFBlEIdwDjZ5d32OZFqk7FXrjoQaEIbWYVGSJGhKACJKbUiLDxbw4YQNA6feVg
Jc+8hnIAQKJcYU7vgTe640LCnFWLWVecCJ0ud4gb/Trk6H2vbDqT2iRB8Avt+g1Kie8z1qmpwCmZ
Avg7KLUmcqas/u1fAKt/suG6Czq4yIUF6OtkcSKoKGSnD6uY15jj/3NHdenKGtahdahbe7hebmvL
U1rsSUiwJy2rRA+qMHQoOm7tS8uzRRhu+OI51Hf79aLFPaBIEuGcrlm9Q/Gasas5bGuOQ1jQhR0B
yraL1Y3uIR8pfZbYVZXenapy2n2NUGklgiDbSTFTx4SojfpaeUtAk9O1VdzJ02Vmmo7+9uV9ajbp
oJsTSyWEobwcqO/GrCyWL+E8ibxsuYn371aGEr9RxAIayymz9YLMtITBESvOdyIZpvuAbm5nlKAz
v3EjHn14RBQnYUwc1AztDk4Vyoz/uRJVtrQfh3Us8QLkcbLQyKenZ0bCzK32Zig1/4kYXG16z2hR
Gfr07lBxhVfqOHW3wFj41cCTEEtxOKeu+MWopAloGjHWBUi7b7MZHI9yIIwhQ/fjo1M1cAEvPVbv
QDUw2qQAwC6PbbI2ZH8jOr3TN0TptWmPjwypQMKzhvlvGHlUxavJ2X/ryyFApJpxEybGsGzc0Z4r
2FNda4pSDjyLFQfxcas++bxxkzKH34Gipt3pCR68bDMr38L8x325N5640rjJvhukmQtndF8SWJdq
Rz47FBKAJfhJ+2dBVn00R8w7maPMNke8LbYcrJG4EodQkk6st2GXh69Kzt7VdCxZzUHkYNgVskmQ
LD2WxsM54porpLwxipzShoTE2jxeETF6ZetvWXWfVwlg/A3/iVsEFrLhmfeAMuiyxkZJn9pqS51z
eXM4JhHr6jPJgBn40TxOOORvFilyfD6C2HNI54KC8lOkwpnjQYuIwGioRumwEt/c9ERUswGunb7r
ieJJNJmZwgB2DFs3AkL7ddVhFZ7qe6qP1D0XpYiIZM4slbU/WZzjQyMz46NhW9nUegroQRHsdTD/
iU49fpkDYj0eEtsuLG4HBmRQYI8IuT1srzQD1rQPskIX35gBecMAmUDNjQvEtKp8Oc9cVwLLRqWC
HrAOTK/XK7hryKvnY92TPZzu0JCBHHAzjuGd3GubCP9z4ATWIbO+vRbgnsWyop8ggNbbpegUX4OG
Qb8Ebdt159XjxiM/iubL2lcdGmZ1MD5+hyXVI5ZDcndvtEM8+HfLjjOzbU5XrvtG6yuTUe92gd6u
guz+O3wqJoPN4jb6gTcP9nZ5zwtiLweR0rYAAuZfZidUjX670j4IonWeEcvFWaL8kQgK3VOycPTL
RcGR/zvs4+IkY6bSnhgmuABsFjctYRQnv9EJ83KnsF1FUU1rCsgyFY0s8KXQD9PQ2Uz8t+IZoleU
DpPzPXkElGa6QbeRfv2Yj6ob7yFYGBAO9OpcTttk6JFXeyxAo38ojBjEZFW1OhvThkNGHifirb53
Jt71+MsL9CVORvxVes/9g9hLITfHGPY9UpSLKGwCLc9DAA1O3rlzsVFk2TybJucO12kpWEjg+GNQ
KYeNXEn8IX0SCyxfmgH/CO9CNMA4K82Bx/AcI8J1v+IRQfU+kNqK7D0UQ4UiRmm0TJ0ehPQ+g7If
kktcn1Pcm4DPHkpG69/qHEzjwXyEqcUeiSWCDZYfZHY9+nQmjhAtf+2g11t17rNEOzcHCX9OLe8i
sFbocK0zf+ecXN8GRvGvsvX8OLnXeuQ9p/8+B55EzH8RcBtVSty3yCa/iVXyKIFfTQ3p0R3mweZe
1nLGP1cbNI6jIjefhiodo+0Veco1RodebvW7OU+Ilz+WhQDxXyK7fOWN6FQM1BLoNehRwEnhHsMO
oNbeRV4tdETpZlnPbvYiNn9qIJ8fFNcHk03f7kzHtxrpZsY4021U7Cat1AwcNcKvamHjBoV9rIO1
UTqPMzyV/HbIHASvpfQ7Fenby3LOrvB9w1Q1Qk60E46zmSohm92VMKbK7m8HCdnrj0fx14hHAxsd
s464tC5wHuV9ckuLEZulNX7alkoj+sLR6Rmx4C5dEdTLznDL6murvLpx/FEi4ldWjk/5X+h6t90R
5jtgh1pRGGTkQa0rvD7ky/Ke1IjA4pLsZ6wTjq+2vTmlDPDtAEbkcVi+5xSEr1y//FVFc+GUYBre
VDBdf8BQY2+8JXPU9896ivkfVkoSHG9X4vhMortelExTf6yZFQNcWjzmNCCmA0bVEtu6iLu32pZz
fxkhmHaHfDksYvJ/I7NdCTwZFYZTxu2ibIyDJTJMI4SE9wKEucWrym0BsFPEZuP8ppIbOZobvzje
B1lef4dWnwGN8voZxGclTKh4vvGPEprFNYu+nGPgGB2ZaTcOXkOH1MKXkn6RqBaq6HKHTMIEe8+f
vBpV1DLS08eV8w6/BuzhpNwsCw5AZFA3cP1ho5gxd8DAufZ6xy0hd79NOQxiLupLkK39nyJepI1i
eKQ94BI/w4uKf/PEuUmPYYUYZ6Yv07TGQoNI7t+YUX7fCdgj0CaMHZZq9TV4Ha87Epi+XMyX1Ao6
K5BN7/dRuqT4PkSKN+8i7Y6d6wVViHr6miRv7bJk/ekBPTwMfC/LuLIMVP71fJH22rNZzY2R3zMh
JIlEGXkBfV60ZU+aQukxnYnRHbxcaAOGb4b0nUYJ3N/Z25lGdS4D2pfZJj9IBSZOvzc1q7en3deG
4Hx4SaTlSxupIUGZTbrOxojwi2WLAh02C8dlB4gyj4ACRb/7HXnEMoAQ773Df5KlfOMpE0xkRpDM
JhBlky++EMfx1sNFfIjYW9rIZTwv6JLBNQ0MrEFPYLP2Y3o5lk9lLmmGsR6pKtWRjh3Pq6Y1HQSe
HN1dV1hZ9AWEmIeujXELyjiutxoO5PaUnM8snzf1bLevrq7tJsq9OO2erOHDchWPUJNKPLBsAzaw
whEezPUPle5+ltkZJrrO6Tbd20vsUuBpgQynclf2Dfktx51V4TSGPe8c5yfP9lVLB40FlLZ4foS+
TPSONAZLfa09gtArRAHG9nFX4+YrtEba3+1zVsn+fdCKXUE+lt1UYc0csV2dHyzxs7BnbaXWlMgT
Qjw+eR1wUQ9FBw9lY4cwZvCxZLcxRzr6c9edaJ2ZZhdZLrlI1zB/vG06tetVUe+Va8Q7u8DcXqLG
5FbHNTMXNJx7uQd2CEMwIJyyjmU1fbJLpkZVrpLZJIhOy6limfv7Nbfl9taDqWBMpYbB4ABa5kCf
BAIN5dXC262iczTrBdzmZIGjIHMEEwL4HukHFeNNEM/qSTfdwdi4JtnfM79MogdsclVLk9qHRD7j
vuVYnB1WBu+neVHZrj/hw5UQSlmXIAh2WdqFTsd4jFXNBmFsduHl2lICDdeKuq5qvNkyvfctIWU5
TlL6eXRrtpknHR9t0DylIlq4fGD+EETTTdca0jZjObxNsFRSh2GisX3EgIXTAoLtCy43y3N+1n1t
XsdIYIlGLaQRtVNDORy2sWr2qzwseHY+O3Em8EDVLmrLnekvWXH+Z/9nhHphCRfvg5CdgJjo9t2f
LSub2Zcm1/zuq6JztcyNpiymgyyFpHHY+XgItfgrxuGOFfRpppa23/XW0jcbzEhOWQU/Cp4hW2pd
IX81rLF2fmyTvBNhcKHHhNolhTWvhu6vQ/SZ0PLWMV9VnV+EoWvZQbTjDDvhBSM5lZ6DZeCWnVuL
apnQJKSrtm2J1yNjRQ845Sa2gHp5yZ4TDzV7EJWGYaKjABo0mH+HnLzZx9lKOsEi/xUQezc+fh8/
//SdStK9i7iNnEscdiUfepw6UrpjjBcHrGGX0HrRjh1SyPw+GYL1KLI8pP0BRDPFzrT6fjFbhA1T
vGxvdDonr44SUAYGPqa6gxxg1Og8dMPzTamidNQ2/cKT3X7X5wo1dF51UHywth7helUcwrLg8dkI
bjqDI3UI7K+58Keg2sW+xdA2JdHtrIczIsCnHQEtCWjR7jblEPugGmR+PWDPAuuDS5P1fjkfPt2V
HSrGjyj3d5keZ/gJoFFj7MLvGg2M665LwvmXEl9vGRkDdeUzNyz98PY+XPgYp0RUvtzUPEHxnhU8
Qs0QtCh/PxqmUqjVkgYjb4QKrg6rI2ZDhao/CPktKwyXlhShxY0oFizdY7WouEArMvvmwyeB2lx+
hKixWHiFfAUozAw7fI5bIPVXiwiqv5G63LQbUympyIG5FDKW9mIgTCUSl70HRFMhRwJU0gVCSCAo
lrjv2wFgFFV6PiGKiu0mlbIRfJjPFTJiCY9HccZpaTwDRSnu5lYkVoFzXz/kxGPZ50bQt4l0X+mZ
WV9BFqhitONYJ28dJZh2/SfzsasyHCmpnjRe/Nwfxd55BV574W1ZSeurS8QoB+w05E+Mg88MeXrj
cCMKnJ+ZuVZXUpdnh6VMgekVdboed/GpEVTfB6zbWlB1prjhW58kWDqgwxxG9x34o7sqtNqA+Tfs
nUXAtouH4HQWsngi09KSbJqY31A/M49zuhLobvzHerWdnt8I+Oklv3/26L9hT5B5k2FbqG9CAuzc
UDSU9aQN4/FGbXA8jMGfju+OfBBhj4z6Hhtr0+IhLfancvEk9sOrcrOmizYg15LZDRpB2d+1CbKX
H6CXF0SqFMnbCtYz9K56QPieZesMeUdgEMMQFS8oz5tVv3o35koVHwEBQHRmjvpBBqJXPgvRajnS
HD7a+RFCB0C4Cc4W9FjS0t9XCk1oqdSDw/R9tyBbl4+lr8tsBunEo4Ae6FkBs+Dvj1Bq4DwydnLe
Gco9GsubjjRcowSXjQpyx8KAxMwqRGDypSXKo9hSvJySCcI3z01ljth68HrurmugsrkjzgEUKSJr
ediaYIYTN5bmtXaQ3rljKFuG41ev4Ld3OjJdO3m14+HBrxRMGrDwCwqJ2JbHdnkXxV3VTEhmbRaV
NCaUuMmgccw1M5TuZFkDxnY7xj6T+ENF/EhBSgVfeAkXmD2Sa6nkDB4b7eGMWoIUsdFgT2HdPblJ
+7WjX3EB9fhDdCMD4iSKA3N5PFptcX36ESp3lf7Xue5AgvWG8rOqaC4TnxZRkQPc9YxKtwB/FSRq
pw+vUa8Amija8Wxl/XqI4KbLBfZXE30lzs6fRm1Pfk9s7/cAnqbsp8IhB3mr/DhvdwK6Zj52OOyF
5IawnmKFEGRpHcFZT5a6NB089kVm3cenC1IWUGaSy+NIj7X16Z2R3BBA9R2WOW1AouWhBIBPhuSf
YLmM/Np5GUpMUDebteWhZ13WLpmSJKpLExZOK+mOLMbbbZvn5/q2376G9Sj0KfX2BVRCS5ZeCFBS
aDf4Gv4PO8ulIUreWR62nqLfXkG5UN1VP7pGIURycB1+YIjMo5I+3oSl+EeR+hgBFXapeaEOlBVC
8c+nh6KXrCSbnYpRG216FaQPmgMv/sfc7Zd+aCUxyibESeuH7CUQ3VJ1TCj/IceLTkIjQ9emGfGX
5lBla3D3Ve++VmpOkgKtm2plLnEfOwrM/vnH5tzRMkbbmGjZt3EZAsMXxHrfdnR22i0abwciZouK
9hE/HVqyAzH78yV9ZTp6ey6KRNlWbZmnVj+OBjzjKZS3BofFA8EX2mVYn/e+FbUcgUirQmIaYm83
1FbhjhOuk9/Dd9nuxJwOPQDrr4qZvAUw+30zbkgkGLvarEuND0N0z2ExKrbccvT/iT7wZUp3g+gh
vsRS1XSYrrTkgh++zvguvd1FAU6eKvR7fJ2Lcvy9kt+RlxGGhyNAqh17k6fWpAPvHdyK2WkAg7Gl
BgyeIe7jGUQAP+994lXwNwUUIaqyj1f9HnSd6db0WcITyxJkpxOYH/IIgjItaZvkuPDa00c4x1cO
RrmyvsZ7Usn6dEsqDKNVYUMaeNfI+Xe9DchNaNLoCsMj2XhBlx0V027OdltDB1EdgJOO8migGPgQ
4EGciKYTvacbIazR6e6sG+7TGkrtQQEUsukRvO+33HaBYWUqx1uCG/avAyzhdFZEbnbF63j64rqX
gz2/R4dXVlsK4ELuzDnQU9pi/RvMQKhR3LXXAqvUBlRQ3wQPCuOnNhSrW4THzkEz+66jtZNxjO+J
Gky2ll2bUCwzxDyn6T4To38bAg3KcP234YvuIPi0FrZPkf5qE2dmaX9CWCoH/m4QntdqJbg1GleI
4oC5Fu2Q/WUil81YdsXx3Yfn90/rVUZ6E4pUKYAEvfgPB9CVwsqFzyNXyqZk5KZMSFEJ0UU+Td9Q
GpqafrtyCmwvK0T173M+LD/Kh2v/KpSbiITcA2jtDbTGtU30epHpGcGKwMeBW+QigoOVFSm9Sb+/
0yQq2lWoms8mHxFJGIkf7UP2KCyxEdTSc53Uo5Y/2fFVDKXou4WdkpCWeq1Ule97dc9+oYn7biMm
ClUHHli7krUmmWFijtDvHrvtVIA8WtDPL/1ywST2MASDc8MZT6tENfh2X/xMmWLgGPQQKLtDfYAE
4hGEx8D4vwkrLqCJLqpgfR/JoV6tGvHteqYmjUAL06HziNPAfDIOudCoT+ETkxKG+F6rDNkdfsQd
4OWpWi9zkkbTk3vb2kd99LvcHaA5UbGdetnFGe68hJsO4tLxcxAC+TB9XGOmmsMwsY74mQQ71Lq5
g8ulEklJsm3PhsjIqgjpqtH+lAdeCrO/ab4nyZj37ayZlNULnL8GdoeAPUK/w2abBDZI2KRjW6MV
E0ANDNEvX/3DJNCpgu25zAjyi1VaNuiDVr0MXhoiK38YELEhbU7LVmwLVbWgupf1/5MyLm2uINd1
/CPV3qxhrPWfWf7GI+yIHqBMYzV13E+vWpeQqMzQdh+MJOJox/2wK6qnMdik5amfDdEjfF+q0qpS
h9RYn/GDhxQ8UjBt442BuuXbpME3NFiPhR/Z1ieZx+29iilFykZuAWiYkmFhjCi5sYu25W70X1yb
5i1LTqQMSGgHvfnDGNDq+HmUtbKizy1XPh0SExxkZjFvvPiXNiFozOuQr66HtVIERjbbY4P5am+Z
2dcI0zhtj0ghJIl4So4u6appukBrUx5ItF+KxqQfdSRRqlYLHDxOUpinYqa6ThhRhcKSZWZfzTR7
4cQaG94/+nyGa0ol8ZMBKw4JbLQ9BJNG8j/VZ0wPxxmVKgsIW2oJKFj4L3fuHj/qYQUVWKE+ehMf
xy4GfbNZRN2TbqsP08swYzbgN4cj+iFNUi0X/WU5JBW1fGNpZomMeMV66H7diF8QpL1hjw6Cb6Ro
bikWxSuqiu0kdANgHfMkoz3whUFUNjKlK0dP8h+YqaQ/IiR/6iSnZJRI8z+zEUCh2CEeEgl67Zr5
/IbGOtGRHhH1/DeaWWbJ19q4LtWLMnYhR3vO2RGowfF48Yyph/fyZS3HysvnbaVMtkAH5yEvlEf2
EYeM9p9EouCgy8rJa9nGAMZUxT33I86OXiq5NoXTLB31r+0QNqMR7lmoNzIr2Wen8iYjtdJxRbJO
MffZTz/lEyX5NKayOxKT+TUmJY4jrQ5mUXwYXKnNXRznqhUdi0Tfxyv7yhc8KtryzY+SuSKOoV65
UqNLSb49rMAmgXj6VQENFvFU42vE4GEkLK0metJIflk6z5+hIMQGOtk5Tmrux5Wfw6weWkGovdbs
Lu3WH4297Ros0iKuGOE7Ymg1EadnFGIzOyyaWt92Fwar32Rgy9ywgHtmNwXCuKHOzhc3PrPxvD/V
Tx8vQ2IJujhtQKEi+HXImOpjZaFPrmcs1e6nZYx3dGGPjsuX08ki+rDiRrbJiWIBx67VZy8TOYwq
J1EoFd/LsYzeniC3+m0qspDfGLh5gw9uiinCVyjQB6jayVjEblQ2egRz9YlxNtI+exsE9T8bzISJ
eTyoTuIa9KK9k43IutVyCTkCy4a7U8iXTUMZjhYbm2MRcPwypm4czKOjzMDuYWmDg47xAIAKz60h
wUhJW5Ikh2aJopY7Vy4d5iGRr1PyWNoXZcl/DsXBLuAZiICbJ0eIg7mrtQyYVQ0nmJ9VZyEsAFi/
fSr5W3WXfb4BNdfCTuvx2iZd9ev8y5TGxhpUcn/W70lFlK9KUd+M7GCuZG5J3H7v/0sMmQPe5L4H
XFx4zuamGLuK10Yq1wORn5RmNLGJpGdlqmTGbj20HAxE30FFf++wd/teRsdu21L6BFZLs6kDcBFf
ZMXmb5hXMUhL1o0GQXJwxr4hY9vx9vtyj3tTzBPxCZnIgSIi9U701mH2/Hghv2dlPeo35D1cROzS
f7fjMpiCI47RUvHR5Wmfr5jwk8ofitE/mFcVhzuXPID5YI2g33s5uqHwTSiuezmeLSTTfW/iSA7k
f+IRXGrSvGV2xoRiZ958UE/bcYr+18WR+xVmqRGKhMhWBMdtMSnxpdLtonT/dczd1pHA8mxrdtmx
HrByl32GR7QWtK1zklKg7Xh9S8S+WYwJ7o233a2gsQht2L9RnPQSOEzLDzCdcA6NKLU2q8KTkvPp
SneQmfUPBgXdiuILlu/LzCwzi0CVmtu0wS/03kxlZl3BlqmEMpxJiasf9rnhQOHpWGPYe1XZ0SF/
1Ki+vY4w9EdQr/1xOLLZeV6lHzeYjIldUgCuqxinAiBp2JPXulXOFRcXSKnMzONAQrc8RxqAVMjK
+tNvpSUL6WYWbAziL7mV1sHzEcoFmI4OriPEaK/2YgH2c23EdeFDO5jdDQFsOaOdFJzBCYYCgZRj
uZxsVqQ7ehUsDU+qu168g9wHfX+VRDU4fPcDUCWbD/pQa04nCCJPiuKjOCKlmTRunQUR4QzeLo5O
wQAc6BIdX+HkSlsmHzIQOjC1ZoKJ6P04Fq9npIvV8YOAtP0ZQ8zYwYSHtv5yP8SpL67EgG/7141L
MyoIQiSaB5p2HWk1W8zaMWV/4Up/CzeO63wCQ6wFdKgNAf/9GDb8pXcacR24Ep2nuak7K8QDY90A
Ywb6NGvVNPFwbsTx8Nk6Oqni1DV2Cak71RUjq6TqBmdoeQBrH2RiYMfxSf1Y08rOhDgowJoVpLD6
QSPcZpa54S/1CWPioTSJTZ/GiyywWIUJnvzTbeYbfptjT8Ifw4IYjM6B0ISaiMmjGhmB08PnBOnx
cx2Bt3LhaZIP6rLy/8z+IIJSu9O+HKXKkeQCDyrqXHxppafJY0dYTRtvcoi7jodKLeTTGMFBEcIP
Uo1yIEaqEOsZlpzNtUD3Vzo4JbuBzl48Rkphr6s4+Ywuxno7hiC7LbBSQ9rqTlDkpV81AN60tcx2
ISqrxORgLRiFCORdeF6imabrK6seJZfgHHp30w/u+W0qhm+c/tLf3itSXQbi8PVg3bINl33qNAek
2vKCYM37Ow5l1lfzmebGZmE57zpibC+bayqJcM+rWdBUxnnrIO/Dusf6JDivg/YvGSMVD6EjghKP
9GGAOLI5D+OqaVScEsf8gsCUE8saTKOb9rrPLGY0OZ+7DDWsqSACwegGUuY3DP5iMNuLgXSmFA/9
a69YzZXuesR2Ex17pVEiMKWycrWiRYsuD4n36NOxe+XuVQ2gADSuxEF5SX3Pvl2bbo+NLxIeHrAX
YOjevxam1L6ffLFo/BcjPQxmHaH9jlJKC1C6OZb7muOVTdYvAEnJuQQnNQCGChqe5chR/2OI+1q0
HJ9/Q2tHmSuCeH59HQaLsfdNSY8KKfrRBqIZ7HoEhGC+r85/5Pyt7QblR/CI7FaEXYbW1iDxMms3
OxzGcfsx1vkLKRQMV7H4L+Ahxq0Dcjfo/PLAopdz6EVgcloUHGihalXvwPACyI9zVDWI8btHM327
ilssNN8lYc23LXXzzVl2vxN8Ndk4HJ+7Tqzk6qngK4xiMmBJxQkqtu1GYSFLLSCQfPEyxVQbQach
bXNvMmyCBTB3TaxLZEgPZFhdoEiXeybx4c6t88wvT89tFa8qJa32ucDBVCNq37aRC/LudhxwLDrm
Kzl2wFpcGXeG7FpmItR9NqCJ7iQqobJVP4ttedfVGOa/nZSOf6YiXDGkRASVwiqKdFkVa/SkrZ03
wCKzASjIQKBFYUeU0CRjhmvRbDF7NZb3FFKpKU0bN2bbtbeRq4cmQ5YSgRYTXeJzqADYuNnESVto
z2wGnJImQWjtkIRVSEyf3EjjDQGq+lDju+Ip55vIOcicT4lUSThus/W2P9Pms3dCAwtHqoh1C/G9
gOllZtyaCHrXUZVdlIvFjM48uW5eVQYUXAbkNyf5zr3G4rrSoED2NbddppdU7CCguCJRc1g8u6sl
p73P9p9eRsDs+lxrW6uQtYd6WqJqtxnECsI+971zExIQ9vqktI0ciJHG0Krt2wSX909jMlxLPDD6
bEmU0eXAT2PsygouioODf+VO+NwKiDsgxGItarg7/cHgPwvCwtbRFJaMopNWdAswAlmzjaRMWi2h
duwyjfIokVSWliy43stWv6YRV+DCj79OBVyt6ehJuEAF4858c/qMO3BZ+glvZFUs8iHYs7Gmad45
01Qz1nCQCCJQKFyYQa9NeQoQO2RLYfvSzDOpXsP+pOPimAPddHsUjtpX75FSQYoo1FF83jvh5wVy
oEUP5PDyYvwqgepNgRWbomu66XWfROHLjLdVGP8RxO0MZ1zwi2mTdPrqLfJZUThP7rhPR3B63LNE
UV/lPwOTlro6R33uUAy2YGedyvMlWIFdSBBNNZniUBlk5Ckg8oPeB3RQDunt5MotbdW+f2yywe6y
RmL84WjvR4IuSyIIiatDXyk8Xk0W1J6JB8AbJkTfAXvm8lEcq/tVwN66L3YQgaL2Jxto62oJpkom
IPHTkx3diKr7HvdoQ/mCzOWkHf6+bdQVqPsQAjIf+r9NbbKxuQv0BbkLxW7kQQsuheW57ikQvObM
Uf+ijdhBmlAjvjZ0M7AiomTWJ2SbOASZFTq0wBoe+RNAQtxYQAReyd1cSktRWLbPB8tg0KLRXRWU
f2+l7RveofRtRHDISNJCoahyA9oAAy4zP38feGGQIFyFPfLHf4JgFipKTEoLMxYZCYG/e8PD4jna
ZoTNSDjQDGJAlySyLxHlKxb4BbrvNDg5aiHTixewWnQLIhuJWM6dUclfH3TC+x8gbsQArB7zJs7D
6n81khkGQ+oFP9yaxguzQnUMPKsGuYTT9Wo/YSaDv3yiVq2RFwSK7VQjEmbFdLwG5UAgtlnOZSe1
Brcsx5TUtG7BBY3G2M7GPn5qhsjVKfhCMfuLLCuBWpmCrxMr5oYYcxBYGXxKZ4V+WBDza3C8hVwM
REvMP1pZMTklBwj+23czFC8p77Mxto1xhkM2VWM6UUFD8SUOe8hXpzjuufUpjYliQWEWfrGvWHwQ
12149LusRis59whwhqRA2NDsqqpGdttVHEBsvBDcjc3rzjAajTgUPVBPnV3xU/jimmWF9le2j2Dw
uZXyW8EJjMMwIC5Gtw3G53V7wFLa8OwREIBxHA/8V6uk+dEJ+XIrzdeK8Yi6aI3tLmL5+gpq2f9x
ClXSMJ6Z4TYq5LCVKXQvMCqu60epTnE7rfx2PpiQCf0deoNPckG7uuEZSgloFcBp1uMHNq+i6ZaU
gO1cddTy0Dzg25dKro+fkuNuHPgvX4xX45+N8piTLojaEYfZS/pW1W+uJHotQny9pkI6Ku/aEm0f
gF9dLcY758COCZpmuUmYh5RIj79FFbYHTvQi4m+nqpMTkp2cDb77vO33HsLkJ/xuCcaGsmc15BZr
deDA/O/uPBChSFMAShwWxJ0attkbsyxjQUZWbD1Y8qg84JUoNnxaNC29naHfi+Q0H5hPT8sUENNp
EXWAVPHCbtNqYM0ngufB/ullH08EwFg4ZDizi77xA1kl73hsXu0hdBDBpsf9yiM+Rqq/y/8Ndiw4
jBZgkbAwakJzrDj4hlv9vOgO8OII/4C3DtOAg6SjhPIXQzmHbLtX5FzLTPvi5mdkboCRESMjiTzC
vyd7PtQlfo4SYb+pTUpkN4GkboD6ixDdFRqYNx3xsfHwtYqHX1WzKh19dYySousEGwcYhjdHMql6
OiTbCObBHRyTbILdZLy/BvHzRadv3WruiuAQL5kx7aF5Vng1tKPaRt9dx3ZbQi16P11KTWJEOIp9
kwp7TuxhMou0Xc6fthtnyn5XynXL9VGuoeYDzhh0gh5slaR6z6g07+T5TlnyeWFEn0iG0JHIa5lJ
uPyP4lJJotU4emJDN/l1Kkw2H7WYa/rnbkHh1OkT939fA/I9Sd+594rAbnRJUcvxc/0hLLfxcZGs
4n0nQyHAYE/cgWAsBjgU2EHzJmSxCQaymMI0ru9nxn2aHk3ChYjDj5/LjakoLNoTeMYWvWz15G47
6WLjXkyb0aKQtsmMUiRFPe5AGQ0OSmQiZodHlg6q4DVnnc9onzAdyVkayZ5zI/w32vyHR/LCkWuv
8QJYTxldCP7LbzXI+JPEk3c/hz8XTnqhZ9ZZeHQJfRmM6RRR3/0FtXb3nVTEH/D6XqWE84LpVYHj
j1DuUv3DTfuH0S9YvGom6aOBNFU4Bxn3rsDjQ7TLiVS2viczMGTLDanDark/44dFZ54H98nRrrug
/fWVyggjeq3WC+cfoyIMLoFH3dZNK7nnY+KzsLcQVhoae35x9ifYFS1Cgm2DhPZ3ZXPKhRVaJ5Dq
1LohP9P02AEwupJvMhdUdlYPk06POqxAgI390mXBmGp7mF93EUUabdRPjhA5BktLTPSFV9JOznJz
6wdmYGSFx6EhYPNwUlZhVotemDh8AV8oSGrGBeBgDpkaLOUEfY8RJTt9CVJ5oRIrFHT7bkToSjJY
DPekvc524EmnBohZVKHpA3WH9nDVnEaigDQUoWPAX5FvO9uAN/Cvu7pF/NL4z0WvqF+uCKoFLst/
bYZPTZoPK+fXVP+RAxqXo49KgnX/DRYrErBU6+CnD/iVfC/DgE5r3TQ/YiRNxHSvEs9CPrkax4li
GEq8g+ai4f0H4M1QPPRWcpHiAcZrPOBt5LRsAx7AY3WlmjPMvGPfYQbqj23GWBCkAY/BgcWVYc7D
/p41YSCLaium5/t+YviMu1lk2Fkgc0Jd1bKrT7RdGvhV/Iq4k+QPMuoAfUI5zkJbcD73/uFfz4gC
V2IcKC5M4yqaWSalEgUVmFLA6DVt/XUlily24z7AumJ07MtuT+q7BO05ZBfYBh39uazu0eRKdIiN
HZI3veFa1HYa/PZhFxrGm6MzPm4joxgNTlcqg/F5zbcN2CNPfQZuhmnPJlzlovsDZ0o9V66zXTZJ
W0MWNYlzR5VEYk99bOnlfgv0v29BTwvHlWKGAE4SioylRzlWeXi30ud52fiB7WOJ+UKU7iKHxfRj
M08UNfgLMPme3RykyZhTTyeNrFtOAqz12lMsrjRCJA+ZhJEp2iV+jPG31c4SIRLyI9y+qIyPkKDg
/fwIDv+3xwundJkbEgrQEukCsifDh0WLW1BfhDR1FTN0afqMRbdgiaBu6XmWGXfbx/Ey+/Phw55w
9Sz1DfvqXuLC0FR8YDYp7MtXFejMU1Xk4akXn+bt69DV4f9jCZ5erhyttyfg+j8mgdVBGhRWqYjB
qbahMKKgueTcQUbV4FcWcWyYZ9yrhUBZKCCroLVI9bgQPqaBABxQIFGe47pZU+W9Tya3mIlgs6mo
BpBDN6nJ343/g7fowdxU4f28WZPKuHWgnob4LaGwwe6PxDMymS6pxPg76hbO05kZ8AsRM4md+du+
nj4fL9x075EYPjJ9Z/4H6d4FAgODmv/oTPzRQISyuypfJ2borLyY0fBgaaZPWZgV2n/8BSrD3Ac+
Dps/dZIyT9Jk4PW1m2qvkzZHfJSvTAg8EOvN5u16w8XvmQXbBsjA+d1njbhMeNbvVRuADRaKf/Zg
8HtqmGHxM8XCRhQK40gQ4KdQtf6NJ+I15WpoFOz3sui8GwdkOmhdqNa9RmxaxyoMlW2wRO9jvLqK
fy3lXYfEIB75f72+JiJsUBxqvTd0o22/XfbEOmbONf17uOwDCmZMgG4aFOISI/JMY/45w78Wxjlm
m6tys4D2XoeCf14uozin5PDcQ2J9m74IQxvNDwrSGrh6pZ6mAE1pOxkLpHNNubZoYrFXQPv+pU5q
hQBZd3cE8cYlLpGekdnFWYGukkdYz10s8rNBe/iGilffjDnltyV9NLw8kP3jx0bXdEKRfKKzqJdu
WJtNoAZNTkYR7fFjLz+TGQwZuYHbQEsNnsFCY2ubt57rzfJvfjrCR6dhk0WDJbEGGj0OcuRPe0/h
caJ/yKBx2G5m5bDA0KN//SPF48XZm0g33KFCQgs5tkErudzM+QUYbtDVOVXSBtaF04ucHFnarHxC
fYDl0YFzW9KtAJFm4r3CqePz7tIVQTdSGaV6hzR9FwTkgEH5JCiRWff1b4Ut4qn1LiVGVhauZtrL
Dm8GBKUqttlO5y8kXei5IDcbUtMUsur3m28xYYJDJ/qOwTD+dxaYNFVdeerbYuqwBmX+cVRyeAqg
FMkkecPwQQplmwfQusrJKhrssWGH5xSx86+C56WXmChGRgy3M3uL+8CbjqB6sO+uc1wTmtQtrCBO
s3cHzXknAt+gGVutPkygJToQgrb5RpkYFWV+AzQW8XOkqH1j5xx33gMuW7bbVXL00aFI3G9tt96m
7bBMrQKyoRs38RObcEk69zvizU1T65D3NuXZDzihsMQgBhx5mnEDncEsu4fJxZ5ve08GpUgTYZdV
qzVNxPq9XokYP+O0LbcGJ6fx8f6w+7Tl92iE7jnpvKscWFi/4c692GL6fnhp/ULoCAUPLF6HtdGr
bHFOtWkdI1u3Se1oiNXW6qpckQYQwJLePmJHOPLKCGKndczsHyD8omDuUW0PE143zhWm/7R/Y1N4
dbA8ei9H6hIIq1Uvdg/Hmknsz9u6d8Ml3aSwvZNgp/B0TwbZMLg05fPHpnrkHPPtQT0drjPCPZPs
Dr3Uchekc4AqwphsWwoQoyWF3k1EZQh7l4vFk6s6uPUIsa5bTgapIsQr0fOWcQmapC9HKLAfNfxu
NxtR5IclbpHj8T9VnN7Qdt6gBsKlIhU+Or4nEaZpOcmA2hL8i+OwHmrhJBVjAlXDaA/qMBZMOqvV
sMYDQ3FaLihR9ffRioleDbXMZ004WK724GWBqZ/VlYr1H6CNuG4gNdF16ArPF3+LJF7rFgy8Rq2j
TJYyNyLP9dk06zLKD6m2RIB0Khqx9EXUHaMQJhJqXT5ldiUp6QhRq16BZBcL5bcTQomM13stWijx
YAZNGideazBY91TiyUrqu7MJnGm6D/0VIOwMInEnSZIfkxWuvFY/Z3w7Q71uTj0OWvH18wg0XFIa
Imv15cHtEe6ZYs8J4WO0TW025lOcizmumZYo4kQQ3VqovKkBMh4YD56JxvY/UTWgJexUM+2SrQyx
3lw7EpsoidefzHPLgmvRyYLwiSWH8CUnUE4F9/pn2ubUKk6f628BLVO+i7RmjxPGnOwis3lJNhUl
SViwGMshxAUm7XWeFpcGwUMdh9tza2MpJhSavd+Xv8qVtc3ocanYoYBGFYoljRNLy1Bm6Sw87Fle
v4EDE5Xz8g4axa1torrHpl73kJjRyMcLiOF1w+LTVDPTdim1Dd4A9tZRnYtnmpmo/mNEhkKqqzyJ
2LtEJG+kSLbItdCheAnQIWfFNN/zhNMnuHfkADQOcoZTcaWiDEreZQxnRvp09kqy4ETMlBs7E6iF
gfd9f0anQeZA4WAFUg15Vs33MSSsDeadVKpurvaiuklDmTHpu6FhVSe6jkrn0HhUk9yjHs4XPH+o
6cPSpKZRTPTlwIWyLTcPBmpfb6zwolOolVYJU6Qrs5/jHxTU2ILxdYGMCIyo9JbkVduMtmnFcAG4
dLDfYRVNAGqzqudpKaMa+WegAUjdoi+6r9rHAsBCPbqmqlyf7vFcNlztRwOBOhA4pcVnKvf4+eD5
DUg1dQVgBdHR3Aa3/5vcfLkcyqLVGLsC81UPMb4fgx/NIx48m3BNVqI9e0YDbHYuJIfZh0538fSD
mZfQqIm10GFWirnPOOkCOqtQH5XdI/eF3jyRorAYQ21qbfUj4HDMznjL120TrB+uBHelfx85FrwJ
J4iTIlt49s3jXK10zZfwJh/CvEKpbL4BgEa7wJb7ddgkCJPjujkRF4qZWKUo2+Yaksx8okbE0/Nq
t/S90hGauTj8fwPYao49fjYdyH1j832Vxih3RVk5PlQvpPsxc7zVgxCtbk58Se4EFAsj0wmtkQ5m
shJzjfxaJtV/LWuT+FJyPI0af8RaHo1t8J5OLIYqvq8XG+W0PC60/9EJTP9wj7+5PZMFsThj1QPz
/9qjz9nAJ5eJOmKbVYqmhZc3gp2ZhRNUgAoKGQRPqX+khbDp9SVmGZQSwKzCP9xHuRIZ60lpoDK6
CwLYCCWdF2D2h5seYP0CoXLlNGbMsCJ1Y297D1fFz5X48WRc3n6yJNjr2Lmu2Xl3AIbIy5Cte9lF
wbAsNBoLiy9K8HnHaFz2IuHGTpDCeNqL/eV1J7hmOLisS/Mlfqf5n6XI22HRa3n+xLHXXBoetmFJ
IpZJ7kOTL1kNE7O3r1g3eF5+qdnSrkiAC7Ny2eBXQkdfmUeN4ICOolf+xJka90o5tu4C5zuGw/Qh
hujXTB+gwHSaS//jtM/ANm2jIR2WLhrTvP/7PF24gkv2ssbYbUqKW/o5blf4E6lmx+MG8ro7GwiZ
ZbIVScgQL45KvBn7LHObpegOWXiZakVzLAEsKtM1TBnHBv2iXCbVzj2kecUgf6aeirQ3dMlTV81S
Mid2KV3PrSI7xpgrBCDyIOF3hPyVo6pSijLbG63a0orlzB8U+AdKdjLVIBcOY5/Kv4AdKyAJCqkZ
ZfeowibtViv8+4aGwLX+9XxavCQvKFS8/9Owddv0zSHpHVFxV2hEbH5Dw5fO8tKX/oEl11MRiZvK
oipxfccsxb6OZ1AdBGmDzOBcyXu+dfz/TXl7c4/W+bu7qaSKTi5JspSDJdZc4/nmLrQcTg6+fX6x
tRVDooEQAt4OWxGnltP29qpJ91McxEVxi12dYMXIof0wx3X4Vqa5/cpBcDIhy94I5Txn3GKgoZpn
CKF4OLQXdOyDEw21sOeA9U6IEhPHn5upY8e3OGw5tCxhM8Kz9JihtkAk+RtF5pfae6Y09S6fTcuF
/Lap3aZPklOYCD00qbymDDbpxK0YhwtfLKfGOcmDTBS+OYVMvHxpAo6V5lFnmey/Pqckod/AkApd
meVGMrnMgxK+gtMDsuNRL8eTHc2nA9ZM0BToEilCkexuXSBJVmwFrp78x+DYzwuYPMWNH4pLYBvD
YuBbr8glQg+B02WYWgr6kLbLnPB4wtOzwrzPw3gmCAFd8xUPyJVIGqKipzEcCEB9+ZikkihYxfQq
JoeaWbJrIcVVV9IzuDrH6eBLmBANcupyCZpK+8vHyBQFk5tg/zchUQ+efwJrKVT9pg+itod8y3CQ
eLw5TM3I8sTAGvIjftsNuyGgvjV2UhdXlkLKHKt05eoH3xxbnjw7ysJmCw/iaGPMh0tcWzY60UaX
olQpj2XT3X7krEVmlsTvDTYtWHaZuq3f4Mu7bUVfWnySX9fPMGW+jtMfaHnCvTS7vvsgbtb4XZ94
1aDOtiHYM8Zc+gfW1AYPUBHf8kj/yNtGrMTuq/gDdTy92TImz4H/cUPVkcO+wMGz0seMohb2Q7Z2
5jXBJjPo21vsLPqVFZdGvPiNH0KYWJKEYflLjZ1Ljz1CtKoKQkNiJ/88wKjxTjsg520eh+glUqJW
Grj0bB0D0fYwYfBTxyU4pLVxY0Eufn466cB5j42sTAQCV7bFSaG8WPYgTtYWckLh/36g8qJs76kS
4QEqNAhS+2c0jhJFplJyV4kbd0yoHUef6Pb5v3Ap7p+d+RFCXnDOz+AT1GSINNaY0kOj3p+MuwLP
ir3ap667rczqtOcVKwlqrS1U8C7bD4gWR7sJKVTTfGRe/LwO65B0ZusiQ7mBA3LRAii7zXJtQgsl
YnN7kilWlE7MyM89Dj6vMQvzz7qujqGKD9B82B8pgz0q9D21HCahwVsDcwtwwWPsbrcgkPM56iWe
LCtmTXb/UN8Nf87AaasJSVmwiTGBSJst9tG7z7GIJH9SVQlPWPoavFrnqZl9oDAJHFkMQWTyWo1o
tGp8Bsll+wNR1V1u6pfGsrSpuTV9uL2le62pQQMgotvQmqewpZ1mV8wHjqGO1OpIRq3ieKl8bY7M
XdM90n9HDvcCrL+BsUKQg8aYTe4EjG5o/EvZWnsq5zg4oAX2UT2iTyg0CzcLAYULJTKBCqiaP9iA
yN57w1iJg/wkSZRsCWvHCf1NTxo52j4GUZwgF0BnZH0JTZkgMHlORwEMkeYsZhmLN0DVeFfTR7I+
3lMv+dbBksLtLfKwfO1Eo99XBtyALLl51EpBCmaEWQXQSwJUmwYk6GduvqX12V2hY+vnEKe+WsZJ
nC2JFtLZpZ2Fkz3Q8mV81u1qknJhqy84/D1viGNsVE0NYiQ0G6QRuFd3BKZGk61eVSCasRFVRoef
Nip9oabZqKTeQxQ1vlXaCjmgSymRQXaXscPgc8xLEXyrzlB46laKWHjAUdn9z60LvCWS6BPuC34Y
qv98c2BHHq2M0vRFslQFUkuqB736rNbBcCjgJagh3l1jr38kQ35T5lqaWEr3LWqVmSHhJcgnFNct
67+6wn3TB0bQSVkOriJgLvheVLyI9I+ffv/IeMlRHjIeLkrFQz9PXJHlAQFY6jCgUinMUKVLu5nU
4t0JuZlE+NPwslQeTlK717zsM4Vt+BehHX5HtiS3CUL9k7Pk65VYcB6HrFvc6QHz3Wm3pYAmgbYp
f7jFOVSOmKWrff+w1CJ3N3RSkxZg6ID9HqStCrP6EyAAJD6lmC9BZa9melpX2DFOKJ1a3QW3Ewsy
nKpBG6WnmOxZTlcn2DN6MgPxO6hxJc2tjZTeWavvfcmW/1G0qI4XnRg6XW6rlPgD8hszlSP2vryw
TV6Ub0lK7y5VPYDVnDYpCH4CfQuG/S9rAajMjMUvNFIBiOjJBKnKpAB1LOOMPnAhfncIOcLiuiOR
CtlzegsnI/rK+j3DTbJDImhcIwUIpyPMP6rPho497YrLaxJp1tqf4DC3vWEaPtNOxzJv62nD5nrj
rjdw2g4W+AOxX1v0O9CN9sNsAO/keY1/stIGUZ4KYuQeS//FzRxGb7a9tSRRqHrTFPHugyoTzsDc
fSxVmQNobeSND1ww/3OF44DMDAUaJbIr/IcCQx2fhWfe5OXsPVIDhlWK9xpG14jWV84Jl8SoXGK/
8053vrJ5DeGCxuKU9LDhsy5eDEwXKvVbOtLIbSTkwioq4mYzugWEIxgHYamlnfLA/NgWG2FjqQh6
NsYCUumLkd6XRCngg6L4COUC16JSJn+eMVjPY5cfiLwVNRy38Un1EZI2pjg3412kx/bocbwx+5QE
AQOzIF2GP+9gX40QVUSEBT3Xyi84seASBmr/kiX1wEQV6tQY/mFPJ9TkB6NuqX582Vjkbu2eMNuS
XCDpOBS/7/ZQjFbOuvZJDc/GsJOXvuTYoMK4elxUENDITJoreaboqgTtva30fDzT5OwQmPOvcyDW
ONcdITn4+NLQDdNQVpI3L0701xmhvsKDmVhiJLLU9JZ1YSlSFZCDVeEozYQO40WXDmd5HrvEhg58
tiipZvlN0lpGiduIHC2S8HicpAWk0yS69fEJN4ltQEdrNZZPrxyZRMad8H+2UBEJlJy6KPMmQ5Yf
XYNQ97cnUSlGuaK2xs6YzbEYalGN4NgnRWiT+YwJcHCa0leOKoGAcWzKUqwlejw9/xqE6fX710WH
Rkak+ofA+bHLmFJNgsqUPi60nf/iq7Wlef5jJz+3YV0DS1IfUirUEeacSWfO497b5UsXIDxKUzjR
qVDAITaKPeMJub0aI3EWaCqpmDY6DyPIqBX7zijawrKzSJSFl8YfA0PmvGEQwKASGbuqLM8F431/
Ag/r7VWNn3XxPR+wNExxwUP/57m3ECY3YQonIBpqnIVC8C23AbajALAtOV6XkKZmovjubDcxgkgV
Y2DkN07aWk9pGQvrwdFUeILay12BKsoB3+HNagBIvhItj6guBtJTEGk/xGjjGoNDPntoj/mKeiud
INohKDH7Mblu8Mlc9WmJXzsfxxCVmZJSvPFUs8zt1Scm2sNx5C9h9Pk5IvvmvEktcaLnnknJuEYK
1GkZzjtPhMPR8r/FrM3b/VfNYVAGRSs5FcjhmLU9uPvHzQn9h7v82Uj3KZ26RyIRW9KbfJUfQKqS
n/YIIulgFM3LZch4xLK/DT7OK7TPsyWQVlyZob8uTkHx7SZR6kyRoK98rs1wcxBozxlJyZBFP6dw
+9beGaQ04N0bMlAR35UaSXKBnnjWxEtL7yYZLrOGultAYqu0Di/yP4a+P2KagsotOqB16zbTk0BR
1xnWtqgXid4HWBdRJwMcfLY4RsStYlmLWeNNRv/e4Ef+vDv2h2vAnns2LfvKMlEDVImuknLlm7AH
r25NqW1NIwVW09iUlH3wanef6BvpV6uahdiYA7lqOaTrBVwKaVBh2Fy1GxbSvMnZOXMTWhUomIXP
Drarn68mo6t/XJzUAvCAAl/AsKiSoS9a8Rlbz1XzwlqmfhqtKiwZwfcBqKMpB1fSoDX+zV34ehza
mqCqiWQFAvWSwy7VrsqDR8+EwrHPwuThVFq0w9XMq3a4PusJMCKYdovhYMU5gogNwBx7pRLEFIAX
iWmrhg5vmM3Oo8e+XPeXvNCxJz8FIkUPGRBUbGXnyTkPU9ZgputjS4R0sKN4c7B6nukTJoHbaNM5
rFNw+75bkkvu2hzQZXur/+XuLvg+NZm4h1MwFyyC4Q7OQFqfAWLeGf9NQ5vq7gOHT8pqdfPoDEda
7QOSD+NFyr3mkiNDQbpwa1Epi4oMd+wZrH7Ih8bkYktfzIOMsgtLTcYHF09mIbYNqD40BdEfXD6u
MByFyV24cV2NDFHvYg3MCbP+F660eZ0K07Vq0CMgPqTTSL766eajmDQi8uDoq8Y/ImrJva9vFL51
+j68XGElseiFMf9R/hKdNrmeKcq1GCES1oyk3FFLs8L5EHF34jQkA9JAypeMXj5pev4DXkH5rqiY
T4HgucAWOnzZqihQu8AY1KluNaAZfl6p6gpI7brOLYdq1D4K0APLYoxaaV/hG+B+vZMo4nDf90ip
Qnad7tMros/5LN9ZII+sdX8wM3WaTvl5mlqMeFxWRa3nFFzMYh8qdN0mE2LPC2PKooAf+oJp5NfN
MSMb3DR2jngqt2kaLjsTk51muzV0Fx38M5UhZQK+l4Hajrcyfj0roKRz97dVWAD06alTTFnMAO10
vMGUAa35Hzq2itW1OlVG3LKFYnLMylpcvxT0Ipf6naGOdf0YjeJr973pJVjesRfwhyyMAlw8eoq5
2tqkSFBu/XIziA1p1AtiGEbyhkchdNQehfsOL728Uwm6Im7Ge3n6PkXLaJy1liZx7K/o3XK+eVTI
AS9nufIulDXvj8K2vq4NG9hoD4877vQaaapL/kIwYzW4e3/uTvo/9qWHyGXhxEQ4DTqqcmE6dCWN
6+zL9KCK4zcp+iYQMvzO5vhcWkrD0Ik2hFXsApBJImukVCJ9GdXU0DZGT3euiki6JsIyhAC290Sr
3OnROXJ6hJd8/4uin1iBh9rZtMnnx4dAlL2XKR8C/EHkZDZ8T4CH/QQgo1RZtTnz8RH4KQJWITSR
VWdBZFWp5HlxShY1N+UdAAvA/DqabpYsz+6UdvR9+H/A6CzY+ML3ZjwbsAjLww2BOHkVL8Dvxvlc
ly0JgW0u6CNqGYRZrPlSp9RwwYoQUr4umQ2vvWQnwxDlSApJvawSmOX/WgoztKXGMoUREPj+M7rH
aPODMnubHcQ83nxtWjOUGpUNOfgIkdS7hRhrYHUUhntM4P7qRrHrFMUypzp2Q9h1ge2t1DaKx+Gs
k1dC9hqfn+wEgdqN8n8uRA7juRkD8jkxrjW66/ZN+wv0fr0VrjCKjR/ZYRmdbTC8GXHqh1gFwo6o
Tts5y6M30r/TfzoBooFiJU+sSHIcZ7lZtG2OM1NccHvcKhVcea5VxREpF523l5flLPQzZK9vK831
ZMAiqFX5w/7YQV6gmcea/lppkMlPm64ti3/KS9eizPGnXOGKfqSqO39YHO/kYExFmmM/+uuu1ah/
fv30Dy4//Dr/lpIkbXE7Fp40+nCXm3G6BE2L3JVZTKRPg3CNHXtBx75/bd9EhHgJ9CALFzkFdCx5
0/BucNsY/G3pRXcWpLbakbKF4KFU6iZpvLd/dnUmXB1fl5gc9f9mjTrMBIAgyT5usVmaKpzEafEr
8GPCKtN+IMyKgt5hAV8UAWLS4X4cUOjNqkFiqvDn1axI0rv6HSlOwvVZRBr517LkQ/MYdyX/Ou5C
7+S9Jk4FnDg20IaEmfGn/slgNwU3aB9Hd/dLdUYH1PSm5My5ekIXGVro4e95a+799PySbUu26bDH
ozFUMHeN9dvkPSmINlYh18ITiCB6iC4FzX+U4UUCHqax3V70kRZXKBff5aamYl/BPWuhrk3fWC/2
Xx15gs9lhEy35cvFySS0OyCYyHotUIP8Lx+hOsVpik3rbCRaxDybIf1HZvpVMsSfpoHpftl49tKh
ahv5uBWsiG1tmOMqruRcTiLtHZEKdU2aF7KQOkawED+vz8lcyuir0O7oCi/PWFs51s6agNdLSxRK
ZsgVKs7RyJ0n7AJqf2Pb46UGjGQJUBZRKuSKsOhya1d7nai4naT7Ba96uiPTT2wqgFQNS1rgDdhm
IzvcCoussTNWmiv6IEm03jqYWjHDxSN/EGEf3/AxgMdHtCLpPSgCy2vO/tdNm7zCxZdxiMxnPN14
1CdABiiqE8RjXJIvXhKLhVpQ0m2mtx3VXlpXj20Hoe84Deoahet9WWYI7VEC15XqUaiKxgqNXeHG
fbwO/403eaD59CaXyFkXEE38KJresdjfiqFAdcC3bZfrxMTckvYz/75QQU2mDh+hDlhmieytXmB5
nM/11S2gs4CNGJOlL+IyQ6AO1S4CXDH68VfF+IroUaCGPuDUnS3mVkIY+mghq9OdPe07XYOY1DNw
r4WMNwLnrggTpXy2f0CS700/bQPbjVPMn2/PX75IqHtvN1IuDo+PY4aFS2AHoK0FESmIrRtEWjcz
mPvNJE6UbvnlAftod1KlAyos0/lScCEITSIXvqrRiV7HVwr8YLqXiv+uXYfxMLfGzsVS5EwrniRX
9+KelS3Jz/H6ukcjRyGNuvm7UfaR/ji1DX+wISQlfOBuyrwVhfQX/JkJWq/SU4EjxN6RYAYA4Vpy
JpARDPwAe7+tH0bwJ2hp8q+MVykIdIlsfN1vYa5FK/EoWD342Bhbo4YLXxmCpaCHfyP1E8TWCIV9
fbIuXsbt89e1TUlF6LHUKpVeNWCOQIy/iHiN1ofA9p57/+WS3K7E8CsJPtXDB/VOJWxyy2Bnbzrt
r/DnUUa3OKWXLmCZFcA5ibr1RuD8eqG+B/SzMycF9M1StXpfc92v6NOQYKMDDKVvq1NIX5t071CU
YH6LsAg2TgWU0TJZi8rgTd6AWK4fZRt6VA3QiKDnvKO4NtRY87QAA5WZzogKHOTl4nOqWPcRwxZD
GgG7/MQWUpXEje18xlZSu4p9uwpILeShV3bMhwPf0eKe0Pok+REm2dQQnQu4y+nWqh9uhkDd7Ylq
Hz1LqnbH8b6li491CZXIONbHkTZPfSIHGgfVxceTehEMwQKuzX3CLS5Ny7NPm788B5xOT8CKJ5S0
RS2TRYAD+vrIsior8EzL8IKkBP6raXc6PGjErD6DyA2yK+2OdDiq8XxZ0jbDYqvNFuzuFtvl1hc2
6MAzLoT0+3hNNULArjhGCwfJh+NTtH8cLCIgUt+11VptoJEn2R9iWNzrlRdbfhYTrmlSgAOEsuI/
8calhco5zSlAXAa6U8lmJWftvD0/2xg2fIxGxOseXU4NdNDmnfFXjLRukFm16OLo4a/rjk7huka6
Oe+n4wKGw5IUN80ExLF9qSz4ZrdILXrWcxV9QypGEvVSmMGx4KdEs16vThEeaPU8hIBNN7iYKXV8
Anzrd4R+mBmDJYc/5LMPFg9Tv+k4PUb8aTTnSOX/RtTRBaNRxbW3JcePeOFw6kLKo4SqyWqtqXaT
265vC7OS1Plyis/XBGAJFrGMoVI0LXnadt3+fiCiyJNWfiaANjALA7TdkSFbmOm4BVCTSVCj1IeA
ikHR4ioKSAKP7oYJWctkRFCn6+tfwYukASuFJobOFgTh2vAvr30PPif1liHIYmWDrOCcQROrgKiP
/3vRokACZ7otmnjziaLBcUv54b3p46vQKxQBVN9y8G1zU8a8eEK8csFkRpxqwfEb06P3GBiHnJN3
CtfSBShRdK7g4FmGyzW2rn8E/M8mdazVlDwDGBh4p8lApz416gBKLZMVbKAYyfueqF6vroWXy1wm
xUTxWETrrNaMplsqoC82p7giZu5mmH2Tuzt/MD2+lV07HAPwpeKOIN0HJNcMBw4b8VAFiXyj6Gl4
Qj5628cx425NSGz5s9/mpaJ3npCwgt9rE3BUpVu/omVllpz4SLI7cKtyT+Wvda584BmkBbLMv1h9
8wq7AdHsMX3xAcSccems0eUAqF19W+Kt3HeWERQP1SxkTvGT7S3IuVfQjpifMWSRKBIQnTWa7hpG
Ij00H4lxVzizhRulv26Ec22z5H2Ym8Cu8+YXixD+oxQPOsl/6DbcYCTYE1TfC4ziE9Yf4TGj0cgm
yUSJabeviaMNfQnn63r838EVBHFtvy/4P1PIovJEC1CjwfqD/nbLIK5JsOHv/53n9639aEQ9XD5d
W3VjxZFxobM990arZW3TWzBbb7fYK+TUni9y0xXheGOw8wTn+bZqXdw5dApTUot2zNwUEy+L3yYZ
J4Nn9bNNNvA14hjAg7IxM3Sd8Wl8RpkPdujvbBp7sqPGllUfGolFYEvYXVGN/mncltME8+jCFwrp
pnBpI31gW0/FBTMxhqNqukqlKrWrKREGeEiNF5J35UVS0SnfYzw6qUsIgaBDUlRVvBxIPZQ8KJid
1TncQ14kGSvI05NzSFbFdhvfZ06ji1Pv0ObDYxzFbXzJVR4RZCXTjG5LMbWHK40wgUiv9UCcFkrK
RyByg+7d8ZSOhlh2xqO1+DzyyQbBNB2SYAkurn7jPiOPmhhSfbXoiDa96faVNKRdFuLA645kpyhF
Jr44PlWqQYEG1B5RttDa7bIToBzYmIG70jWSMtFvrBl5t7HYMNVECsktqps2mXJhQtFFFosynhBq
k2ldKAN7crcEgiBwzKDEVQKctLGnPEPo6LQ608Osy9ab1j4JeHnkjaAzCQ/3x0kNkkoz1nm/44gq
ItRnKXTacN65U4HYwZYjVmhdv58j94SeP61dIFfCqvyquofKZpXMWCMp38y4rM8+KaEfFu4NGH69
2mnD3XVx2/lFo3mH29lmouMqGSKHtB6oTg7/OicaPrHl01qPvjlBsmnDAp0dD4GqNWNYy9gq8qua
xq8lu9unTLlglnwrvIT2EADAJIoLJKaEpvIA8V8U7vju25zG8r/8QnOtW4zzAw9/nyl6lpktFQae
97FKCxMZhPa/3s2wPh5kh1xWOMgv3Yf203BUzi+sYpE8/HdNUeMABXc3lkEHW3CZMZL7La/rSSH7
mhEWNMskJbJvScvyT/m7PCsjEFyiJFBFJSb8qB+ruMzl52y1/ZjDMWLVJje0DI1Mg0lIthkmPLX3
CSCDi2vjEHi55dCyLzriUNC6H54Uj7AIPD1PejSIOY3xfGfWdh9enPaWHil6HS9AsxtCRE7wa/KN
vCQU521tHnNXpxIyZqTm/3mO3GHdoF4QGpfX0KP/4C60vQjvrZCywtEcYTeKRzPERPxykmSG/krC
dm2fS0VVWC2nzLjjUgcotGr+URxQF0V5o6q8YpXNQP7Rz7tzukigCuoiZiN3zUUpS38TBdYRLLMq
GwM6ZXtk/du/eH8yUIogo+j36RFC9c/AIqGfz/W6hMIicZqCRlyhVRjeLOTSkMN4IUbmlTKzDYxm
4d3Pg0rn6cW4VWCvKkyC7maLgaPOPu3t1U7I8LH29WXEenD2Op2zstB7KAl8TM35cjzHp3kNC75S
FS2mqj8Hpcm/LtVixfdV/UQlRD1ULKlJItH9eKtMRR91Rh1za9+2twxgvRPKu4xnQpoTHbtwxQk9
UxSaXFb5HGyW0UoELUNXC6fbLOoS59BvOlWCQvDxHkH9ie3pkEX6JJx+pRnwS1AngcOhaXEvHWbG
jyFW5YiWb2iZgVsQ/eqeqVeW764Mz5znRmfBmBSnOfsOAhi2rEFDa0M2eACgaJCYwFkBaIlRH9Go
qdJYZkKjYa476jxBh3k70K7c7lGX/HNzd6q1Otzcrg0nZyEx++x/i4e5QsmDtnKBhPJWP6Hl5Lv8
lkAQQMMxVSgu0vxhfF/DVwPwdbTPW1W1EvPVia+ma4N4vP3IO2YFSwALs9MtGG0NuNoJejFfUL5s
8SdhmzTEzIwpUH0L3sYUYZF/tgyCGxikL2xBdayNTBTU+doTLFgZfFi3LjzGjZWggl5jQGGkboHK
BCh4+lmMMwJZsT0vmV1S9nSxDHkB3im5B9heL9Xrl2fjLwmZ4GnmjQDsJU3CTu9eyQWgdOXFL5W7
pxVEHsV7Cd/3dods6qA3NajyYqJqUHjN1nXAPwsKTRagZSusTbpon5h9Xj+OTYss5ZdwliPEgLNd
xG/+gXGnZQ/Dk9dxyPbWjBJ8Dsp3jJSJ7p2OBMMYbAW6Wlv0GpfemvcYJB9UF4Z/tPtVs8RD/UjI
kHKHGDalrkHUnoFUIAglpsLa0oryXjLr5HCBJT0QkrQaRGVVm7uoRrdSweDnzR9Pv7m3m7cgBQ/Z
DKlxfF49/cXVlxs0YC8ISdfOrQ7Hux2AXhHNARSLUrL1ZmANkzXMjue+qTkIINWtgkP32VtCMXDv
Z2E2I8A0PdC5KI+TAuPnVuN/Xk2BW+me97RqrQmyKH/bZmfR16q4XsBYBVVs+L6AqcwuUqntsYrP
1fOvvG2t/DeidG8LQEEuhyo4lLd3+JX+AVSYu69A2plEs2wQ0Uez8CkEV9ad8WMYYArpDR2/YzPo
g37XBXA/sdYn2qKlT3PKcj310jpqGMs9GKXWD155eOzBOvLLVE5dJ8PLtODDd48PodIhyRn68fi4
9z03r2KiXziNpV7LuTVLBOtfOBbsDcu41RfLdTfdS2wRKZooDx1bryAaKuDFGum+Y8jbgMjOpSNi
heEYIn2xDLnuLGOhYzN8dYfP/XQ0tykiPpP4uQbN2LSK7Og4+Z3IHYtUmuzVDVj9z0RbQlb97loV
qgdE0n1UzvCViyFM0gUh87XNFpXgSNVZ+5AF+8VNKuK95CkNrCcT6iVfPFrhykLixU2qa6rgxszm
xSyIBmhSJ9NJHEJELjPcWmdivczC6K6VqDrvVnfWwkAFwPiY+u3YOT4WERCLdq8TvMSjMb8zocKZ
7ADiF5cWENWPVlprRG5CgiCMVGpcdUoCXi0m606Yf5M+aWvRopNrWs3OpribqW+xt0iaRvh5h/GC
2Xgx8JVUkWlMzLkPCE/VN4JlnI6CuZaW283ZHDwg/nl0FEpCgGYQzLCRfZFDGoAKFmqDuM+iJ2zz
Q4VHknKR8cM84aEadhT/LpmdOaWTMztMRnM8HLmZ/QVMAnlrRtDMpMlsg+DrcAb4j/NcqSOg82tK
zufaNUtyh93HM4x2ejpAzbheL3TBc2cRnIJN4qOVO5AeL0QJwcHksJ4yEG5NVpdgDlnnBbqEHdve
wCuWn2od+EexCRgNEMK2aov3QNehbt/N6ATeVFl/bxq1HU1wSIOYfV3fJ98mRgSAObQ3OInZ7nr2
0YaTapbxubwuQMs1JWEzC4zNcSUs/rFUpWvMBckFrEDjC3qS8hYsxiiNbJTEJzPze4uK6J1IRuSI
EqO0inNmuT5NPtgjz4Nhv2wmh9ml9FusAVTVaQTQ4Vbnz7sO06sI2CiBp+nUvPjJWBv02Hzy23bj
vR75tM8r8PecAMeuLaQz+b+mBm+IuNgpjeque5b8IjaeX1JBUr5vw/OjbmIVySf2OsRpX9QwbyAm
2+nq4BdrANLHbOas36TT22EOvG+V+Wj4zgHhJfIjyJr7Y9slcA97CVqczl1HLcUTw8e2XkxlD7G9
MQy4j9vU/VDway4WZgfmSLzVLwYt4XrlBEMXgQ8xeS75lhtGk9AE4Kki2Oyy437xkoPPgr57XXnr
FKXhROWIcqlvbwp6eDXDyBh77SOTlf2AqBBok6AKC96ulPGe9SGF5D2ImBLavgomOBqVon9ttwZU
HZbBaiTBTz5l+S6XsRxfyrSXojIxwnSGfMv8dO4DcyFUKjmQO9WQwsTieMQVjB9UJYilX8mBi+NQ
icNm56e10q5e6g0VQ/f5Mi+MK5dtiMjO0kLVaApS+fYcdQdXloQ/qFM2NXuqVeUkifyL55QktkwA
N6Os1ErMWaK/1DHVpe7gtlk8PreZdpElQ/MJRagRDtXQ6nIJOnBhkuyh98K1K+jHlNdxrDnqqMb0
PS3xeJEfnFc0pPvCV9MN0IIm6V8x/cIWjhOJjOjIPIC3ptFlbppy6qmkWaxTt13AgkYCm8a5cpdA
xF7VbDKZeOk1ez05ULPxa63rpu06eutAvl5uw3IzKjqwYzLmhkOYw+qjRucCCJBZAHZIMWIWUlfP
h3pESmxba3U0h54km1jKI+QJxqZdGmsj4wnBel6vGA82JxgRB7pR4SZ7SKaxgAm/S9lRsz7MkUBm
z2skfpK2jvVPs625QmvpEdUqhx1uOB0CwTWbKMp7OlApLxukKzQHMzLk04TdHjp4hWfAeVYiVo1W
DTlSykjgpjCjuhB/Etg71SOUILBlREYDdkNObm+KyaVVk7s3ZMaWjQzjYeZJSxVXJmMUtw3EV2uA
NpG9KKHX7ggbiJrRDhT0l2+sEyyq8ycXSn8LSv//A6R6kdvIB3K2diXbPGImyhHL6b867vgQulYH
/ENAHNwsjc0r38Ycgz9z+1Cy7zDEJIPWpfF8Z5Pe7PH8xpndYln05teanWnFE3+mp6HgEpAGhVI+
wTs/xbHb6cHI5tYG8icwHY2eQbX0BObewwc66LWupKOY+HcQ+GGHme+Uvrwndbzk0WS0AjC8M9Zf
sk5u9DMN4bl++l2QPT9ye5Z0jBteY6GFuRgpcWFe6I5vyb14dMU3WEXxMaIcstkMQ5i2XLy//T38
/hVch+Izs1Iiv4qLErGuk2/mnjcagz4D0KItUrV3PAEuvxDWEYEWcQE155N9JA0EV3tiC2gt2ZeP
jBhtDLGGWbbXlWphp2Tppv+rFLkRkPRNH+AHylcQOL5sYezdMEBaCfJ4ABRT3ZolSfd49idHSeCU
bIRF84/UEbXX7bc/iDgEoYmS5ifrhsSRetzoM3SzaTMaK1ow+VrByGmq+AuXUtHPFq9MKIm+EGwz
QMe9PLRgfClOvnfbflCjRj1v+77rIcu7Lj9kHTWHkVGKqD0Wffux+jMpZJUvJQkjbbgG6+9lBOte
9yuWgwUBbsQ/jw30uxX7iLnJCeZUD8xeT7HCqV1Mt+N3cEscT+PfwadDbq9GWnmjw8JoUy9oRCHM
eh793bCMTXjnSyREFqkpO0OKKJNtRbhmskD0SgeG+z/Vnanhkf5H1taciLYztVNIo251P1/vXhws
Drwxt5cgQsNc345zssJB8YIy5GBhkh0PzdYxHsqMFcWRiPOp+KW94v4DWH9KAyoJzL7H1DLwarB+
iDLiJcT5g05FTzcGIIn/vB4Nafo5OKFkDrr8AlHnJ3rCs+XR9SktKKpaP9Cz+ActuYzRtXNte5R6
btUH12XaRuVETi7jiqkZagnfIwCrdc4uVaSuZlB7aXVymlY8FCxao53iYPuA1ACtilo0zKxPVTc7
mng23kn4UTlspgBO76FwE7kYALiCX/al8AbRbrmiiFVTmsu1buv/cfw8/tIoY82LqKEJP++J+tJs
lIcuteAzpIXptmU/xDjyk0FsPt7slp2+tqmysGtowLhKRPGc+xCffAh2M+Y7c7F6ZNvLjeQOcHdr
KjTwzAYJ/1kYn0Zf73N3Opv2xl6PgBegHeWg7broBA/jaKSHPekwWspnQ21eW/agnpU7xVCo7bAc
g3ccsTRsJyT+WxcF4V4CHOlRFyd1Twe895rSNmy0+aHgIMOti0d3V8d+mMg7ckXHc8RUr5HKenrT
k2MlDGLf23yYdGnwXLoQwh9K6eF069GnnNaos7tmJ7TabBvjavZ9GwP7BT9Esh85jZ2Vd9OywTXS
8isehgeJ/fPFAu0KHhABcR8NHBLga6TDjs2tRK6cyGU8XwLtJp6oVKK5RelgJPnvBriIuFmXphJV
cnm3xGXUdqlMZFem0qQ2AqmMw9mBTmRaqC5UBh2ZutD7FxHtI+sPN9jJqMpD1KrzCzue0QOdZGrp
dxnpQfc7xa3xoLg5Zz4xnAQJ8opXTxJFHvZiXMN0iUQJomiCK9bCth51Qjg/qGmfVVi3hLrW5K6k
1Q157+BeYoWWBhFrnnq9nspJ8DYBBNeU1Kplm3OhSjfleP3izbrCqt42kMMe1oYiWzY7CyJbg4mR
62UODAM78AQLNCeI1/VJmM5ajwRpXzh6m5WTh92iq8uzT0wwMw6dNBJHCCAJNAhuuHDK58Csp+FV
IHYwLPXKJMABzleXOn3TYKiE4lhCoEF6vaqV7zMa7j3Ze6WgkvVregTzb/kgT916EtVPHCCTTh/z
9HA/jG/YM4+L7vn6J0sT5P4He+3EagE2h5yYb9LXmns3gzRfyso+uexPvd4OLHjcqvr4Uxhclg6Z
Voie4VoNiyBZSnAm3RzUzvSa9fKraYrI4fmJRrSgQa6fdt3V57erpZMdfIoXVOPATYcweylJnx//
8WV3x4ItbSIelKTqNnl3ogV8lhi1D2dn8E2RsaLK7sIU1qAzAVqbGBD560szaT9DEXMpZDDcLN9k
7rULCgULyuIGwGGDaGjsYFlOPjDKeIHbsc8MbuomERmUK0V12ATHd4GBAXxP20TAXUzyjskY/sT1
S4K22/LeUUPOVYp0rlEYcmaN4FqyIsBex4Zr9115hwggB99C+6/is+H50G2S3BxWhl/9+xdRq9AY
6TkANr88/2mOwgcdRefpDkNhgWPJ5HPGO6pj8l1+d8ScZ6iGo86bkTBXeVXG2IrOqoZGlD+My3J5
Gt3vnnFcXxndUfMq614cSVf5bEy4PQ/Oo4219IRc3fVzxQWOpsrv16kzEzVh7Bck8FXJ0yB2oYU1
ptfF2Ley1x5q7EnCzywmxOMOf63/paJN6ZD+LsxwvY489mbNtFj2vFV1R84E+IJk4b3px+5JCOnp
7/ypKvNjreAGb0JrxMRaouj1Yfvl5Ktm5Ai2N+/X3j6FjHC4Qq36I7Awe8MnYyJDLEXZsHov9TXX
hmuQpTx03rCBHsK23HYvr2uoD1MKnv0FmdwrQgKG0O71iCMeggTotALHl8jiNZ0RlUBS71l6X2Mu
8tzeLXSQYuA8W9tDMUzT9xTl0Ym6QQmu3KpUEClqPhwMUFtqDrLipax2mnSQ7Rn3H4vVENUFAKGT
RyKKhjtpjTF6pBPEv939P+pZJAhSeATzRmUTEY9602C+BMKkyTfGu/55XgJ/XEEXIqRvdf8AuCXy
doUlP0FrpqPpVmPSiD0JZbzunlAp6PBYHEW+5xHyoDNBHCQ+r4wzPMV79kSAEqpdvu6kBSkyrtzm
VxFuug4OzfMhSrYjBBw3vBy+UJ1Bc4JdE0kSBG2pGvr++cBkTM/QPG+L/44WcBO7ULmnQ3UpTid5
xTl04f3nQVrzkflJWEKzu7U+0mrZNrQqjHhrP9KDvQ80CEqch505ENM4UAKJYJG6xSYE9YpvVsnL
fdyUC1jv0y+r/46mQFJBXYosfcBoG04pdCgJUOchHMAhsjnbXb0GiPWgL5q/CY1hfD4r2cyOCAjG
Hsd95YuLLsrsawaoz+n+u5B5ZeXxcHb5pTmnHvj5qLFU9tR/vQ7lPuNAsd26SuxAiMbQoWZKNlE/
JObIgm/ZHqcI35txRCabqAY3UVyj18vYAzDccxXTtVnPxEpnfslHgzMQrwQb4NSI+7NWeRD8OmN8
PDycrIHW4S3TGm9F4NVXWKEKQpQ2pD6s8OiH3/LzK+OPXj6K0SmARfQspEAWttnT09ppfK0+Ifbu
le6F+O/4LY1rNMYcrVWyuXqzFve++nsH707Er1cKaEooNXYE4U12tJIs93gpF1aC0fFXWahZwuLZ
cEAOvJba9OVpOSVloOiIbEJYPv0jrCcR/Mxj2e3SJnSErbHtgrYX4dKBN+5GbwzNrzxsBZ25Diw7
GAm15BpSC0hFpy0ZCE5J+SPK7VrPmNgwo0IzRtLZsYfSrNAdFpLa6Vb/O5ptxIZONgkIAqnJYXXX
tBZU1jgK52skUZkxEOf92QCMB5fvMms9sj24Tc3pLqBfcyVjJjVlLeRp9va8uxzHO+AZRlBNSerG
Y3FMGf8jK6exmhqdDzoRBDx0x738HwIsGs8R5fqpObsCr3XIBAYxJA3bdaUMxqlQomqNr4T2kqow
6ertnnwgiUDqN/lS845JrrExiw6VvvLJOua13DgfhY06A/M1CVKeG05rufw4PiehMtLXCiyyza0a
xfGmZFg4D7aU+Kc0aXVtC9BJJ8NcXDaQGyCudKGm6/l29nVS4xZXWqMstCF4JhEva5qs0YfkLDe1
RnKirGvAI7IbjNfavQ5/1sJDtttRSyalwgFYypMbaCUFgR0rhyiM8QUG7ZKLyLHoazepE569uwOY
I60Jm8h7zvJobxAGbRCoahJ7kgh4FRIel4zYcB3BE9Dy0NEqOMbhhDz3BBgJpEL0+j74LokWvCl4
OgMrxRWDvacRQvWgYrsRd4rLcdgrPtFTY54pi3dWKahR0fyM6HH6hHnclsqafgrDkDYI7NN6aHos
WOZE335I4/xzDki6eiPe5IdBcvAeTHyopCYXWAYxinvNyD9FaW1ZlW4m2T47nihftAmORuZ2AFjK
phC2wQ6/D8CYyw0b5/tNVC5RCn+5q2tQoyMVaOcVv8/PCMaL0XA+QM4VfMQVQ0PxlRoZFnlGFfOD
HUdZ+IKVaYPPRdfsnY3vfHkI/ErJ/OiUlMq6LSHrcmsnbh4dzYG6c71eeg2bkQT3riXWBgsCQyLr
3T2sQ4NjmApsN9TBPjuahcokmsv+WSIw8rlaml3RIPAMOFgDrxYrxiwqaj2dvfpiwBg1uUSDjtEA
NoIdaVrTTMuIF+2k5BLmx4eFn0Ti4akDpNkfUeXN8aCQMsicFcKFC26uyxP4JhEysFb0A0tf409O
ptFp6TRaBdHdwlxgxTcKdS+wCXDZF6u52ILeOQfm6vK8Npm5ycjcGRp5t2pflbvzoSyMZl8CCV5E
9rSJ6t5ZppGm2qy2zDbP7aD0jaKep3CXizaqGMdWCzANaqPMsvkxKqndW8rU/+k15oawA8KtHmRd
gyLTiCNIogMD5iwwl78gf98LmWghmn0nTKl4jhb2gQsV+oQuW02yXLou+bHUd6ReW70NkXwuJejY
Li2fIQzLOcDYe2Ry9zx6eg2QqZUlFwVMHbhl71lxUYQNlbOkRw7TUTANUmPqJq0kEpIYCQp3pJ4Z
eB9tiHDa6n0f9bmG3OMMOSHfoOgZzRpydQ3Yl21tHk8HMoiDNmL+bG+0RJPGLr+DX63aT6W0OBTM
nT4IhSyMADEhodQYdb+jSYJiYCrvO2Z73IwPljWtd8K8OdmxpIoGd2kgav2HTpVup3HXR9d0o74E
+IjRDZdu0GYYQbhtsYAQBTkkhgNQrsW7VUBFpCCW0Jv/TOIowAvULE7Y8L1vnEq+5hIDGzHQrrrR
aoBg2AHJ44Gt9+Ck09zT+x4cpRZH6stfVUsUvJIkHAspb+ghmHxhyaa9cpFSnSOr74UDNMm38oCF
aZJoQM3l41LmAvILobsZQxdI3+qzHE8mqdQVtNNG3P8ArVGoSPFHYYVDA4t4UG84X6xZvBPW3QQj
T7E8e8AGi1YiMT08XNG/Mf/z7XZgS6S2PPx98FHw0dOrpkwZZIcEgyQROPcEJ6TGCmbwOTx/issR
bscI7hhwjKTEfIDjH9zH0I3LZdIYxRzZkyfjm0A4/VhKCFC1ujQrG/dgHSRs9SO0o8MoWgx+SqUr
AB9vf7J+Q3qKYZdyuKSR+FeEW6Vh1MW4DUGTDY6M6kX7P5NrqtjckHC7l1MDoxaWbQ+XMsSwPb3Q
l7syetHnLvH9gD26efKQe8iA4HcR+w6TfkFr9yc8XiSQRqXKGJFUyd/DHzkUNEp2+Pa3qrvM1KMi
Nux7xcstBngOkoLQrQIaOplM5KD9VAMVeLYV2pd21Ljz0wuPYgLwQWmyriUcV5VjRn8LxWuIcGqL
/ZDQX/o4qkxCog75e2IFoG8XbPJXp4zG/oqudfgO/eSpeknbuelmzzKZIvf8wDE3R1aV7fFhChhe
8x9HWyY004jIxxjWuqr9vz7eVtT+hlSxERHUnpdq/Q0Qz9qPXvTqbmnwdtm+xEWDJhRSVJ5yVwHz
cAZQ0tN/bTAJmH5pf31REpxDHczCrVXjfWEtZWquUSVZbHyr26ccbTnkzA7Ew7hL8FGq6DcE7QH4
njHdPo06sJtFqXKkiUTpt/jHSfXtRy6X0EisF/rLsf7bvFjRy+3ScTUGJ+eTVbMZ6dL0Hpb65ecc
Zgp23HbZArwPbdkj7J2thNifTzJhxw7tcmOpj0NkSL42J1U+OZ2h3+9oCD9ty6hck3nval7AdEL0
oHsdYGxDvqAfnSW8TwplZLreANXhB0GV0/1ngxviIh6+KxTv8PJG4AgWIvCOOOI8Ioaz/JdFMfQG
Hl0hL3T4mPMwEvjyvBk+9Uc278S2cE+RGaNDW7NzqZd7vFFtGHklV4N5Erg2KMffHPO8W6+xG/sQ
5aXhMQ1m54T4u9c0PllIWli1ud/UVZOMkAdMwGoav9xDg5AsqQ3dlyhMDkqezV1UfmFyzWJEtijm
tDSd5rNVlaMVhd9EQEpDuQhSphyjVzZX/Mk28BcsZDYp1KCzw+b8fhCAvKWB8JHCkbyrXHZsGmYk
XNz1Xh0yvNMj0Fu8ViZ2FuBpQ/1K4NjQ45kKtYJZDo8/nGrfG/wY37B5zk+iORub9+dVzZ2lgt9k
afnBYt/hSeXQct6EdZdyvjHuttw8D+MXVa+rzw8WeD3gBynDyzu6ni2nr9UYkzOK4qmS4ASlucjr
I0AxKE1XLGH0eaejnYrY6nhOH0fZYWREEsaaNw5v1kbnYDF8moKJY0rYUtmlaYI7iklM4waPGme+
RUJYWcv9MbapKsN2HZGoS+GKMg3FO7qOhzsJUgDFlhY2gOSwvQHwGk8hEtB86LjW7bIhn89oT9SI
Xvdz5ldchpLD431NG6+7QvcPT8EGMpM6mfVUVv+vtRUvelLBap6BNF4LEL4PuNOXTzGIYSil9Sba
xFmOOK0nUQYUhLG0aundB2niD2msbpE8QNqdukTjFlfMoy2a1cgGASJNIOLNif2p/uPB8vNsyE5p
jz6z0ay13HnwXo/RkW7orGGQvzKtWSfeR5L7KJilcAcXCWkRsw28nuGsmUh8p1u/tf0mdw0/7RRJ
YZdDLzNRQcx0LVrgm+eb4SuG5e/oe4dg/0zyt7Y6+F64mUWf9p3Xxe6VhRflYOjQblTXn+6rEnQ+
gI0u7I12NhTRC91ISXaSdmuZyRRF7SpPOa96S2+P2u4uLvC32k1uXVVV4OGfwL4UHP5v7AdVNZ9L
CSe3PEd6frv/QsJTjy+Wg9frXW9d/Tr/SqXE1r9Cfp2FPzU7qYyxDUdv29zIt82WsZ/3j7+eiVxf
LWph7z4PNTShMIWMHx9kjVEzL2gX9kkS+G1NcFTu9h8sXqa2hkDsFRWJH0b+eeyywnazZCkgzfbI
AQyKo/2erc6rWTjzqB0jQsHNPXZpI6vfV6cHrpDIZCDY5v3W91MAgffbKhx9AxIFvR41wpInJUpm
doOBLeyQC6xaIpNiT8wdxyHSzQ+3VGmXxvHf72k/4acthNM+5/nYQ09+NwgEGDeoGto9fhDTyOYs
5DJmKQ4PzF5ZAqcoKImA+esqCL0LnTiVTslqNlLpQHGmD/1FzkAXpDXaTQoH4maADoq6jnJ6Hf0N
6zJAqIzqZ1lqpQwdUj1rZIJ5/GazQP3PiL995KHX4/bkFv+mLVA4yH6Q0t9Nwsb2Xig4uqEE/W5O
eKU+gHTGI93XyHMb7mez++j8qIjeQvtFAfNlJgsiFmd2Kz2sXftcEEoKG5F968yoP+d2FmogcNvV
ElHaTCmeO2BKyFPfRnAeWwF0YFQLZtc9NFYPmcGFSRoJNR3loU21JVodxEv1TmaXeyXOD0abvnlf
gu1e/ULniICyk9mAbPfd1d2dmnqecuv2qPkUv7S3rRNztFHqXu1KIYj4gLTIcZ30Rrl3NX+hDfFa
l9IsMemUGXVxu8uNr7yLcFm9cGb1uZeEtqGn1LtIKnmz7aYw81MNIJ1Fuw1xBLBkBsXhHR0saurQ
dbCTztvziXfrrbrSxx7Wr9aVAhKhPIV4Qixrl95dp2sjOZ4GoJq3c3+TyCbBksB6LamUVJRJn6/+
bn649Ar/8SVvmZDH0N4eUUwSAOog/t7JAtiTO3su9jP1abHBwwK4J2gYCP9fwYeSYHBDXiAJjZH2
eRVArQX/0wk+rX1sufYAyQ0V4s+yV704zM50NgPdloP4EXZHHm2SBXERFDAjSN5WppTLF9Rbpb0F
k+jKX30tmJcT5kRZrtgLOxSPQ9xyz5CA1r1p8qRdHcYh2S8Jx89q7HX6dLjxLgpCqsVGktab3GAf
mF6rEpcLQGZ7jpWAkGuZ4CqEIH5X3yw3tGieJhdUnYRAc7T1Ch0t4wTp417zfO1CQa6qkt7WVbLl
phT8mVOzK/12qCo8vFdUZKIoLnzyH/noEbYMtcQzJ+d5vNTh3IXzFNamBedTeILlzr4ZdSIR7ttX
tQi/vWC/+FPmc5mAI+7ikAX7Wc9LAJo0mc2cV9q//jPXjg/Zry+b3enzM1BO5Xfjvlc5WUaG3zcD
6fozGjJqjbL6zcQlg2q2ozEo6AScpt/Xd9+NNdM0S+AZquBo97bYnHY7OdzErIgrpSffjeXhokHN
uBpQWdG3UDuwzf95YZ6x4sPj2v766bd7SLkpyaCTTpRJI3KxvJxF36qfQLgdWAExOwO3CGe/Qj+3
qZXs63cQcLLsoEmIVaNoKC9xnfA2pPbjPTYccOsFn3jpFtEORLBuArnlL/XpC3kNDZ7W3EFh9PWv
UhI659r6PsdfkIjT2uNRyMkkz0zWN2FyANxXOOHO6GR4NitHSwmkqUPVVky2BSr2rYplWnDaOnrL
dHIP9/tqPoN6OlbKbIoK+qszjWp0y+OFFvfkWUvuI6b+63D4odBJm5qnIziRmory633Zue4L205e
9mtRJdXH3PiReL539Bcj9YJDMZjNNLXb5WaWe32HUPkbV1z8+IGAOVRo219Mhleo0fpHxvuxmCAh
Ye0fmAwIZGZFF2fVKHguNCS2Olx3P4FEfkRMQFp3D3oI+k/fXrKtoz9uyDA7bY+z8mS2sVboc77I
D+o7xEevG3AgMj8fhHXpr9NFgJGzmkSRCqfFarzBKfDF8nsxIBdLvfW7g4ZM8Zy1/NCoer1imewq
n1+umZAjhVBmt3jdtwrBTT/Fc8RB2NE8NJdZrQIZHASymaesp5LZGUb4ZPmBmnXa1R787DeuEGRY
4O17oPbfRIzX4oIpChVE5H+AbV5yL3k65srKGdgepLfufxvb+bVPGwfFLSbD1efudYjOZXGUx0SK
VUmaiHXKFt7MAjzT2lSsKET8P9Kzl3I8GcfjFTR4KVbO+SmPrLfIxoU0r3GAwx3RbeeCjsX2kjfp
wRHRJyAUhZRd0Bb+N7prFpK0KbVI07gnlOGFugTbBnn6EuKRqdirGWp4I1B7cQ04iIppDTrXGXoV
s4t4Fq1IV2qV9GrEj6T9i9keaI+tVPwMriYJd0qVbWvmvjxMQYbACUk5wgJom41GpAo7NGrNGNMp
89ydLWiCAoO7vYP9IMc1hdOFsG9OMjyWNHZrnzynCtK0IBSsRfAezdQm9ErpQ1T3wuYQlqs/rMCg
NOK+3wqvnNCjBY3rzfG32oVooiE2bw8fJA8GYJ06D2C6Qj7IGtz1XW4aApRGyf+QBlUgTexGInIs
c9EP97XbjIQO1FRx8FToHLaMgqJXT6GyqFvQeq+/awafDok83NNGOW8R9xPgiAjP8TtK0wCZd8Mt
S41VgnSnqEgHr2lvGS0acdloQu7U2+VH0qBRf91uvDokNsYkfGZ1IveGaWMQYD4+lCbkoMIrf+Kg
5ZSz5fIui6xgHvQSeArT1drKpMr3ZTUv7Gtba22NRo9oaiCGETPBwndCWFnGK8QsoMG0BG2q6ytn
4z83iBqBLCyLih+jrCdK12hFUrsMZzd5Wp+TPwTl6hssI8nsgWxWCkNmgCdcQjYbRz/5lhnHU5+5
0jSWRixsE+YKqFHJfBDcetDlT43VMoWs2EX8gEc+YmXA25hN3QLHzN8zJS4ABKnHOaQ0iui61fN9
iHKCF8Xv83t6EIJ95hvZ+o6PXjSvUaZ8TQzhNFbCXMS5f3ad3HUI/D9ubYxBiUY8ZKKwxeVNnD4B
+BhecRf9+nQnQpmB4qn12+csoSj8YdDHKdzRoejyWbIdE14+5k+W+CIxldS1YAv++iLaXQer5+vz
KIAwrtGWo+FZrXa6QUqIFKkjJv/Dx0brLexN8zBsAfo+ppSaVHyS7Rlr5we8x+hyiZ6kGAXzLxLA
2Uw5NcgNvuSu/GRwLkDHC9HYwZkDD4cX+5DUZfdsZKioEjRCYs9E4ljEg7RZ85Nxq0NgKpMZ1y3X
z/2dy8iuwi5/tksbnv2+ESh5GkZBTLEZM9JEU4pRlBdeS7at1FtzQxgoXxc5pWAL+xEj8WYlQioa
0TSz2pLQD4IvLhdpyP4AzvbZ1j9wwpae2L1A8p/X/7wVLVgGWdutCJeSclicRvg4qao7O6uYJ/7o
iglO8VWHsvHxGs7o4gKnU0FgHsJQhn5WoFm0CKRu55SGFdDskcXCoSaEAxy9mXg88E9FBIGSTnVr
fM8vQohlQe1bIGkwZjElK3h6hmDbbapr7iTdhQ2c3Cgw5qO0HrhJ7ZWgitdpIc7/JQo8oBiLurFO
N1hoIupCSqf8MRcKR4miLkJ5P4DEnp+GHSa1fn0AfMKz2xYcFTYr5CH+LSist6UQ71kbnZUcwdn0
EwCjkMAxEN0UPZSt1lbvrdS7jtjo9mUJHBeM8H+iz066T8WGSEHc4PA0GTHRG7U00eXlNJamFcgs
O5G7DMPG0mKeVpy9YcCVLZp3dh6s1Qsaq1Caw1yIfeF7g6dpsmsCihYnFQ7DZEYWnGBpwtq1lpBl
t7yLgfsDwsS8LhCookHJ+KJO/0jwi81Op7KbbRQFyhsw1rd3pts4Fmxi3OVRRgE4OaFVnCh9OKl7
Wl473DOr3//LHhMxzWaHm7fwI0zD/iy8MsSsb/KqzwE6MIlTOFNvCDrk71ztN9KCoA6oBjRiXiL3
ALjOPLV7gcM8IemXDEUDp2wGH2J2yIUGxwnLQXRaPp2oA0YIEu0C/rS9Hb0oaOxPPdvAR1yxWYBM
vGUeGgPtxFcM4q2SCgf8kLKIySlQU+OfPjUp8SCePFqalzUQLsRtqiBt/I6abrslamKocVQHha7O
YlFt/sMXcwQhQCLK3S6SnUSFWT5lb3JZZBpBKHMdtAQepf4rFnPA+bRpsZciVpdEitXFhAgSx/5K
I7dB3k67GAeeQXmH5/ysZ1BOLcmfrmio40DOPgZrFbaG4IlrR/mKphdNgogy/ROmJwbO61ENjfG9
QR4NCUQcBP01nu3/XNzu7InGTYVixno14L9Y/Tw5C9mwbJXwrZRKHZ9itlkKbADGWFuH/cZO+2cb
TEAVEBZKj2Gv8hzIRbL7sa9nC2FDCx2aJhpNgzs88lbIpnFGdkg+5dJ/0S0DnAVMAbVLTkEnSZUw
wAkZZ1vltsIVXPDfJzfLFOkl5nF8F9JEKmOyWwK3DlHYw4x4dQNijDQ4zgsZQv9Q6DvQOenOjU4/
IzpmQ5m8JUpv3cFsbqrVeglhfcrNajN8KDZJytk2XCR/SEFVF7ZGihBbvCnbAa4ME5PsPBHvpmG2
BabdQvaYvKHquKbcgIZ7WtNMPpQYgE6noWPpZmFv256+FqknjCKWil28MnPX32ypTUjZ+cznqjxD
ajGsul/m6QfrcpD62SooG/52a7zKt+kZ6d/b5mNv7yV9q4Ic+WpdmN5f1Q7guNR675KE4wiv/L8s
199d6LwdIX21mpAZRaUTk8KZLyq1l1E/C/zSL3SVHJok25EstNy/sauOlWlJvSntg1C32qdPsXmI
LS0w4PZ58uFc6x+IRQLnZXppRvAoEJsSv2C23fXw6vTrxw0y+HNIhXjXUDRxz7ZTWALkAyDjpSKS
22HtxArXcc0WVL3jMgnxTHHMXUhUPxuV6wCD6oouB5RrWi1NSoD8fz6o4KiLaMAimcBuHu0CZfTK
z6tOzzHaHFk/0AyclEHbppQQhgRLpdAtkYwCMBRc4NHeNSGlR483/vW5omvJHcqQ+Yf9qBk1Aa6v
4MmTqfCXOd2JPKE6mFmgYPQGQIphJ4SrmvQgJZpNsNq1bpE40J6cQ9aa0hknKvbXLMBVgR6DkHW/
zNUe7N9IedY+6XNrTvhebk7G1xOYj+hQeqr9tqHpdEUMUBFrvre+IaIyeHSajxksO3Q/i7e/685k
jWOAPzi1oFfrSVaIZFyBGA/ITGvYpgUKLjulmk58+p5suL+MGHS78Z+8MHN0mRuZse2IlQ/lze5G
LlHDqPzvWcemXs53s0FC7yKnMI9ygRqytlzGkvd2qriEGdcL5CbP6PIH3p9FFCTJXdqC9PGKsGZ5
o4UahO0rKVT9tbWgsbA6NX9zAy6KGsbCTEpwaEBNg+7ptY4P2YCUfq7eJA3904dTdU6vgLfFakjd
Aee0ukSCad2zPw/VlH6dSKEsn2rbEGUorpzZ/4ZCuuwleM1dkPz8sa55O48A/ZR+jLqU/ZGhMGdH
4MZHh9/+FGPQ7wXzB74bG4qKDAXceZzHPUNsc+lnDxuStvTNbyuPMCHDHJ9LTnGqV/Xtm1kGSM/3
g8MFNsQh+LGZBoMyr5PFSlpTeb0/ZqoxY+ObiTkCqtOAZEvE8aSxcO5PEq2/5MfpqJKEibZqSwf5
v9gVZwbo1xkZA2oiClUzKd2qMo65JzuIzJalqTzrgheI30EhjXPPp/V+aHQNWZQvtuk/85v6VszO
F+AP8QmNhljjO32VbhYYt/cxbBTsOKA6N1MR/2FsfUpCvK9zZ2yd7Vjj84qSkh6n+UV4x1IvYczj
VFnAS695flTWSDkN/fS1MCCKOHUqiDCFCZLvsfYp4k32W0B2pYDsPLL2EF+jUE+A4JTg+Sau6vsq
VIDRT0+FZdcti1w97S/vhiVe2N7OMWRAaBMXH3mITb5pSBRIs9FYJwZEA5leZnfdadbyjnCzSN/y
qpaA2HzftKC5NVyKFIsrPgTmb0jGD8i5Gj48sD7gUtO1bTDapehTkeRbxQOIUCt7K2R89yie6fyV
aMlHSSdBhsuSmjQF4XUUFHLfMPR6WUf059Drg3xs/+xFkS/7huLWbH8orxfVk4nbDYGN3lXfzs29
ths3GqAr6uXJvtBv+KaFHNAxf0PMktUlbPGlg1whHXKfm3mEWYkzCuaQ6MFeyhNsQjtiI/e5FFkp
Cha2C0qYoDnQm5r8kUS0GOhy3YMv8R48apb2k2zJKiGlkc2ImC7bDuAdWb9lWURfEkzFx3K8J8Fo
eS6V/QVm29iGLE5KGry553TOY9yaHyufB9FyXKgpeThC9Es7uwFwUrXbpEJF+MjrJRclVg7KoVPV
403/snHmT/K4U26q0q75BpXZSMxTnPXQyl1dg1MEPnP+S9fHSB9rQXFBpE/YpGAcqriH2XT/LMnK
bWuGfDkOoPPgQCixpnQyIs5Key03v8hhY0FdBr3emPxGlxH7P00CgcKHF5HVhxOYwMnf2xLPtDXa
Ej+sLDbGhCebOTrT/0uzuj7TDV9BvTkkenJoWQ3ZpEjGhMlf+tUU2hYDXrg7R2CdT+L8WOQhaBA9
nBJVNmkp7hdu9rEJX3C6D+xf+S43j0P8VXvcu38V8AixUg/TNrDuP/MyCpGQUM+4evz1Wr4TqSSV
w0u6pwdJQuYM6qltMfBVJLME6mZiweX0GE4A1Cv4VowfpPcK9gJQPEDpPgSlvW39EUk4grbK/jf7
t1nPRj751xVeYc7TtBABV1pGJaHrAU8tmi0PLQE7mms3KV5Xh6QjIlxMvv+HzLijvev58+OPS7U4
0jgYJK8r3DBTXGEoi87bJbdAmcJCuF8atjcVyuuAYkRbOlKNXZGzKUebgahaHUlgfL5o5LsJ0+P4
yuzgOumd6XqVq4ByPaO4PTBLB2jnp5RMtdJmQtaPN6ftJE4dwIlHLGIptrbNxVjyElQ24c2XToWU
pP/PFkp8HdgU+1vvxRLrPhiqttOoAFD69BgPh6tevNyzzNdCYTZcmbR49ovuFDg94Gz33R+avNyN
fMY+6xQULSgT2ePeEa+qHZrvIjZWodWI/V37jZFhCEP+zXmEeP7aJE+s1/7x92W/zBVSeQbo9XYI
/jbdute9OKRGrtPs3LLniWNSyJe2rhwSGBLdfsfJ9Bqls2NO1crcorp8NMeUHtN6P8nNeryELqQz
7NnyS5hBXqWJWW4+Wtb0xhfjcRTTI2YVujzAmrqE0m6MIxYC/sf56DeR5zfUDRHPCS8TqVrRHZN1
QdMMz13kBViwJu3g9IAY/CAqD2/V9trzFjgiI6RJ8XEfPEVqX/wHGeJhP+vt0vP3kc/MhSGgXB2S
cRCImpJPxFEVL5PriVS7OShIo3dazRhpvoRkotS0SK7rtIgJjDDT1KzauocFrCeO0zscNHj3R9PS
SzubQLkUsvBeUgF29bj0eQOyy1eJ1d/3eDNketf2GDFQyC15Yiq3spCNdZg/555Jmov8BjikDt/9
wIxEnp6AJsAfsqnPjCrZOI7OyNn9ksFma8cE4FooQF7XkfUDk0Y2FeoZEl1eKowkqtsJzEwHNB1O
B6qy87VGek2EoOOADjvgSEetcKK/mDAf/dqA2GwiZsm4QRjx1TRvyDrNiGIClqtN70Rbbu29LSgx
SzNON0dazQ3+9ByKDE7/vDowjEuZ3niPLSHw0nfWPZRVdsrThxAjBx9A8vYsVLhE3ctQoNARIBqo
Jp8FsorXf56L6Lfi2uhNV22gVQ34FSSknr7OgR2gLWbhan0XhlDQRAT/99Pnvb6SiiHcbT8vLuo8
BSt9tidVrnK+36/WRKPq3lTU10cndQ/R5oLQrhdMXSMtkUorhnXksniDdHtMRLqIRv3QrP/W/IKD
LWhehK+Tg410YVROKkfcynRpcdnFGeZA5janZPptR1fk9IxI0eDb0z9/VjXld2In6JLSy3JcZmuU
6cHxdwBK9vEtU+RI3I92ikGgEGJ7QDjxuSU0uq5xwx2aQTnFaSdSIWVyaaNR5/zxku2tjoEUeru5
99/6fIjUSoJ46y4WWyc/di6QMdEgQ0KpX2p7/8gSn/7wwitG3yzDidHkndH8qPE8TpSvkf276Jsr
/Vgyrhd7LvU0AflowKTJhptCBkJeMugVNffMlcgoZjXA81gQc++vmxuSFWjeqm5OBBBGTbg7ee2V
LkNYk1yxg9ZNSMg8dBRGox6aty/uj1aWu0B0HzpK8zWBr521OODyX0yYd4RG160n55sj5Kz4L9vA
cj0qPG/KBjDPe7LmkShSE9kcpLzUGaiBf4Www+ml+4ByM14cb/GUKN+SmsOQ3bhHhzxCSxGE7vel
n/pqzHSyMktad1/8YXgZXWLA4T2cSjRr92A3HWgAQF6szld7IXiGBKsdJULJH6XJ+vqimq3SyK6W
+W6jbO1AjJbQrcCzuGpmayPwznXtVz+6h74/eNU6U7sDiU3uo67Q/LfOMRQH0xEQKoj922wsxpjM
9zch+dfegPz4uZQaE6lPQP7Kt+fZ3W5U41pK4dIuJnQqa9aNDdNdvrG/v0I2rCXE5R2X+Y3/ovG8
BmQTmjAxiw708/TRG5202OJfT/NDQkDrQOTnNQ6q88JeV+bVTxqRE3OxXDP+GM1SzX6uZ0qMrF/R
K6/cc7H+bULH48n0a4qmEbth9JfwX3JP7P458xxT3FI1VF6qDVpCaEMeezInWM2DnM3C0YjMDYgo
ZrAZS8Bo3vxN/KqEAOo3Ov4ceiz4rP+cimEVbt4ja5SUZaK756ysrOh1HMDTnBVs+aiLZ7FrLZaR
azrziPU78BdwGT6WLADlJ8IFxQR2syT+KNjrLb4F3U8yN8Ft3/V2bihNNc4OH/QeN9NsDWj4Qutl
YNh2Qqqw1Nvo7Fuiqgq1KTm69c9r9r1VHISc4KPqzS6IrYInaLQelJT3lrzPsV3jEWDyikm6/Non
ShQ2iDjIQlSDg5ttqMKcoOBEQiaQqQudHH4cNj0wRr0+nHdbF84eaUu6i/hWHHJZT/8k85y2Nh6m
kiK6YvlG4w2on0OinJrji6sAzUwtq1d288dKu6QddFID0VeSR1/ruOzWSkplcAEA3PNOMrMSPrOR
oiJJjUARiqNN/dvQSKVsQI/K+1ik6hR7DP5v7Sie7hhoXqE/rtJKJ9b95yaNqXDgc6d/b51bNG0y
nbnfFEsf+P6ClzmaMiA7S5JpTdXoL1ZT6rLQeZq6wnKb71/gWLYcIvFqKCiRfIPqIHTotUOSwZ6E
uPfH7i43pqD8mnq0JmNEJsnlRkwZo3MCVT1jmvhBF95fCBEPFXEqPx5pu7n/rlFZ8fikHH8Ul0a2
1mQqtPfxvj/qXh5NoQtwBBVbvgQQ5yBdB6TbMm4kn0oPtLTcAGOH9qVZSehILHYuw2dXHiFZsqPW
TIn86c/1OYaFFsjLILLFakeu/7S0JNJeZe03iFVZhVIGgAa460RKkdajafxtW/Zdqcopotx/fCH1
DN64igIZFxZFznsohqCUNtrOUwdgT2PKSZnsehlzRYC8+RRiSQycCshdXWFuXCkiTA+tBKczYk6s
drglG/FLBae8ZO57UozlNpbOexANV5L0TtUP7RQX8/97PXA1ZRyisPUHn/TxdNg3fFa58Vnvr+su
7KPD+cexuD5tIW4k7AO8Uuy2JN37pjvn7iRuAlZUfPpkJXPuh4mKe82Fzj0DSOJx9jwzfgthoAU/
EYgaMuzJd1vXmDylLi1LVxUTUZjX/xcpt1vgxGJQyD7PDQkJ9NRrvXxXfs7UeOM2HX4Qi5h+170t
QzAmv5YjcpUhJOqcJ9RUmiHVGFqt9GBO1jFNyDff+wfsnnBaU84f4i06P4l+STsqPdGdBf27z+CX
4ckU11q0SkfZCwlXFCnvqq7rA5Pz8dSXCkS5a4XPBPg+LpG+v2DFRIpvWu1JE7hy8Nsp6EEgfhVS
jo5DGGX5F1Fvp2uCMCJJaVbk6/1I4HKHdzcgPBnB6Jt3JU01ji/8fs32/TAFjOugHRR6Sl+bko44
WfDUTgjqblSOXcB4VqSal2J9ZxvWjbJYZJGztnZMe9muJ3KSW9QOsxboneRPdqI3u06YsmZJ8XH8
4yAT1g2CE1YlD6wt0awtwMfdRXfL1db45/JS7YL8GCBjM9gg6K/FrK8Oqjl8ddn/L4KtgxlSEO7Y
y20NzfW9maO2didHUvXXj2gMNhqqY/WLW3/8mNlxeF4tbFCIVwysfTM/l2I9H1u+EcK1Oi102AR8
PyZ6eGAkugjd+u2jb27YHIGdZuvQ8+S841f0xhkUm7xmK5AE1C50LxNh/spt2rwxErf6VSh2u5tj
uFkZ4joJw8uNdAKevGPMPRtJrbyf9ynXa56fvgUn/So3xJ8IlgiSBOKisHBPGdInAaQaZjJAZmct
W1vo3f9TEqwO/A+ybUvvJ08preG9+9KuOqNuYqxitCVVdn6rrYRUzUeLYqKFmuRNMS2sjflOKxzl
CHP7nCHIENyA74q0+yI2ITdliAk7zZqaB4r8WcbHMtil3cUpJb4VWICiP2SAcLvDt3kk7eaoas6/
ZdIqa/McI3pcbjl5jYGXK1YIlHoM/+4m2BlPfTb1eOtCcpTa4pKVil7szTArfrQLHOGB8ZH4H71D
FqIHhp2FCjJUazRObJM3DrKYDzbge36P9mFuyGskWQJFE4jWDrdarXt98UjT3Ay6+DbJUJmo8aj8
KNmtJRoWt/DXSxFXKjVYWgWrrUo8am743ICl4XQSC2N06+YekH/EOv+05vmdR/s1BZx8YmtJfkEQ
3OwRmLBfYXsD6nBTsxwnfIgUMvibJW2m84tIkZIJZKf0G3JlXL5eiibhPOSMRg+M33ThWBglKXVx
KKrUmOXX/vnWv+XEthtDl4OnTLPnvT8G5gKMjLuyo+TUb/m9oAWslHledUub1m54T+nvDzT3JYlk
lJKPolzbleQfnbxkvk5aggif9Lvmv+AsE/YboF+BzAZLgPqkQwDMvWH+Ob4lVoeiuuwIVHVxIJ/q
Kcm/VZkJ9ruM0nas+svk8hhclx77F9ETLnQWschnBOPMe8J1bCYKxGMQ1dwoJ8v2sCJ8THoyYQL+
ic2fcMed0NUvaafjQISNAjNvIxyLK3RdC/Soq8FPfbAK6aawvpa7whkXdNgIr9GNV05+5Q/pA4+w
yGUIKnJwmWOceY+jExQV8sKA75VJbVuydvvhoEOYEYs7BJk+9jSfy36+49DHS6I+QCtcYf+cBkWm
McGHglUoWgIaN3b9QzTKLJWF3WlzE77cXvibMiVthFP4oDnHGxq8j8FgtzOT3OR1n2xpfey6ZtD7
wRC4AEfc3cSptWbe7G3CiPxpm5g4sMxTXNI63bDZXysrsbISZMxR2KfnQYOL5AuBbWegs/F7gJNS
1s3uLfIjCQwO6lMO/YyHKcWtVqlvrpvSrVNSBUHYc4ZfIxgKXT4vWVaQPdCiZU4/qj8RBmElsn14
addV1VL4ZyuIdfgeT82V1wmZYBbOhhG9vUfrlyZLSkfXZW9nN7djXTSLTa06AlImPhzgHTsGk1Mn
8RVVD14syPixu/0RhfG5dFl7d1BRNe/R4ujidKFhjn8fjqPrvJElLlZ11U461BIk4Z0cVNLR5gGu
hOL7p2dHsXCVB3knEySC7if7hzs5e73zOP7KsOGRiKJOBX7b4IRDjbFZCGCNzajv3qKJzZDzuGJL
7el2haaJRKAlSLEW8kZOHKBOipKGWBoxuj7YYD6J8cBW0msYApJM5uAnyVUUlJL39Oq5we6t/L7s
EH0TS4HvEegJG7DXWi0wDHm7lqK5PGe60xJOLso6diG46AuZrNKlXDGXBoZpB04niNJajB8sYbgj
jM+/J99R+l7OcZ++mrTVvHrnCD2PynSNNeeAsTWTPC5wg8CmmfpGQav/WCvJ34XZxs9d2SJKarIs
yDjihFntrnd8LeRUZi7574aiF3Tlpdu/1rcfyNjv+8zoHDBT5lKxOxLcvzFGw/UY8HJ+e037U3zi
gYCjWNZNPhWbw48nuLSVFhjyA/fdkNnkaeYcfgF9lCjYwtb0WsefVZGuchQC9jP7EfoU2nihzGJT
X1T3eEgwTN5IO4sgsa2w13Mk12yIbvhqYRWTRWDO90cQ9f4765z6KoArxd/zjY8mgID/Ko8l0hME
XaDFSh6JK7+1VTTJ9jC0YglLutFA1PpZq8qVA8cAo9GhXHcafgEC1HX5Ym47NT3SDGcSsFJ/8ycv
XWImzrLuJeQx+PQyekirHrtOFI11hRqrtZbESJTxik5plaUK6y1zCjYsHdo8BT5dUj3qgwz2NFzg
8wYx2SkhS18qnkVvwyHbkGv9YnuBK9cHB+Wc/JbtGUQ74iuzGZoSiGb3UT+OXwC3MRBk7+aoZQ7P
LCNyZC4Ysle9LMhCRSKDCdbnBfYTAoO4WXnrOcTLuxRMlK1Z7KOVz/Vc11D8iiDUOxKl3Rp+bfx6
meuHz8cqcEmHobe1UjoEzz2WFw/rT7dGUkDNAateg6k2uyGTLPLIBxdQbANlEmGvc3hY+WAyuriJ
zj5IgBqMF+ptnUY9nQyDLdoLYcm3Ik3Xt0qvR6cu5L8oo47uBvZF/D9lCjnDUtSu2tVIBnu+HBWF
tCVarceYfy0zHhO7Ty130jxNoAik0CBHPIlYtcGbSWQpbjSfFutjj9pTbP59zX6a7oFq0ciNIf7M
q6Tyr3R4EYfxsVrzKe4JmyTnnzkNeHxJqMaBu0A2wjLuT+jvT5msghaWunBa9bJzWH3aVwaVKOs9
xCuMhtEV9r1jKRyCxq4BPw84NhvGQ9vaxNjui2ddNl/x+Mpkew5sMX7IQz6Mmb61Xqlrj8CWRQDT
O3lj7RicJ2fC3IbbokKNzBP5p7aZl0JAREL9z5HsJrCKUjCeWPREjodjEpH6M8T4omVdFnwDLL+Q
2l1qqeT4BqWCBbehiDCjCOKvvyKvZlIdQksg9qvQeqGtkBuhMXId+DLHWA7dUMR7MRddOWYclQ1P
mOgC7BtHCjnO6qt7NQMiatCkxKxvWjfDPd8RcLj7PLGo8npBpFaRgXMon/GL8p2T8JDbT+fgwksM
jVC9CnzFAnm9P0qlb6h2QNyoJ9PcY25uuCLtgIfFdmjBKxGi1gaVaG8cyShIOeoSOl6MWyBKfLfY
/ZTY5v3YAkcmx38z4LYcYs4ErvJVwihp3LUCZHyaavO84FU2GQp9flySou4AVvVXXuxaF1bTyCdA
IZD+lWV6fyEytea7IN+rdh/NXxzZC5+SB3UWLuNxCHjVuJGW8aPeAh+hoaXpiw+WjIu+cOt4XdgB
6ILeBxs4h9/AYsLMQfkAab16FoSla/UXFpnXH8+ADzJ0O/hidE9rbpuTkeJPkbF6iNRWmOALlwK8
p9ykzLzu75PuMi8Z9ye8NE/UsD11jxsJJZ7bBXWPGBTukb1U365oHETjlSBFAfFREN9QML4lzNor
tzrKi6FGPf+xCZJvbpAeZ4ve+SpxmGf4sdNBuToeGemkPuxPO+ez+Swatju7HKjgbKhxweSQQK6r
2KX8Q90+YlDN3NDl+FvxW8fot26nWsXRPTQnwaGtM//2MMfJNcCIIEyzaBE5Ng1iQWzAew2KatyC
FkrcTZhpp7yDdTqc3q9MQXOzH7qWb+GIMy15hLav+pYoVhtk/K9hpSij5fXynDwHddieSNBHzupN
nkpLgFbe6E1td2Z5OA1MI6wc4E5xnM5p3MtJs9E7i0QJ4k10bZqES5VyxP/aqrOj9LG/QrqfgAIH
ON9ZaJC1REzU4ttIo1GbS2B8ByUEgX5UP/bPQ3mRq/SB/ol6iWQurVHktvnsYY/N4Rhp2hT2U1/l
N+GcTVG4SczUdWVqrYh6JHFDNsIKs9nGD1vh20nAFpu2Hivy1VijgI0of87HrG/NhaYBBg1mzdyU
RIqzxqr8pqhLhRl+CbjHCHn838gM/A/GUzRHiFx0PREjLAXTgo2muNUPkxhwYN1/m6cemAHJXKb8
4MoOhI0GWkNAqqvy6qg3hT0WE8bjfZtx4ZvrT+noReFvLkB2ZYbllBgrdtwdlIqa3yuXHZtPWxSV
TL5gxjknOl8Ie+erupiazq+kK3CgYZKtxrW454i1QPPGol3ptw95fIF86lvkjZZRW8a6Qhu/7p46
FQ/5dkoIIFUWm5+jS9G6/KOoxh/aU1TWbIB+cCNRQ5ohnlOi9NYmGd2sLR2TSwNFOHx8RRvmrDO3
AoZVyj1u+CuseeGoiZs5+TAGBZhWVB9E2Fc7zZJx/9vS5DTLBLbAYe8sRRlqjqO0qMzilZSNDCuy
pFIOK7lrhMexnPp2kl3LrrMM6/en8LlGft5zmpfVD2YEmUZ92JXPAkZPu+HZB+zRk/M+/NXDAXBn
eNCo8FJIj3sHinYaxNONxVJDz+GadmxS4N4Zi/oozpV+msomRtiTuA5QJOUaihA8Rz1G41aiiLEJ
/NzqvRiHsOyKUUnoyk9oJvbplJSDAXLZlCjSHbbJW66Lehj9+fYwJjQp0gyop74omeJwbveOAZIb
/sXS/f7FxulTJNBwo06TjItFp6ZHcaO8J1rr6Xl2uAY40WiloCZztl8rYKTP5chVpOMILKyBnQFG
Wv6VIBfur4uDeTn+z8EzHv5v8cVR9n8JWYJVzwTbsItAF8BaM/uLqMHsXi8ztl8PDO/ISNTAELfb
HaBHMUP0wLDHbdSOJNOuK584hyhH5F9sJ5m1xifMp363ifeCgw3OFmAVGBYqRfXzHzY93Y+Taudu
Y/wfI1xcFAXEH40wBda0gQVOgSYbscjEUG7AcdmrOuj0zLcp4m2aCagv0YS/RcIxa8BbSnItjcz+
rNaJOSLUsRJkIhj/e/BYs4JkixwSsJWt7RVGPaFjOuaLH+1dnaYjWqvZr5KILuad1B1KlnRz7JxP
sdBgDDXrjdda/8bpVymrZ36xOpl2WGTcnbQ0LBkWuCotjYfb3Lh7GvtJ2TE9VeObEehWxl3Qhmb6
5XEysK89HbwEn4yMyeC0xyGV9afn3RKvQevRNXdJzM2UGuuB7co5hZNBfF5FIVxTjGuFM2+9X4tu
hV2d/fIhtPRI2PdkTIwvIrsRnERe4C6PxVwbzQT8EbJhKwR8siAiNr0vGH+wUpD7I8PSDY1NpP09
G+ctDWGp73ThEnqyJb42g8Islp8xDLw3GJvh92dJu0+eC+cetFgTZLugLRMTreMKNbrsR8grqF0i
bCnYn+kVN/QFQSglOk5IDjxK6DPQ+QEr6pBNi9ih6Ls9HRpeZDSDmQyOju303TeAsA59Jg9hgVy9
hcfUSo24xs0ROjXq9TdqYPVgLuzEac8UH12ngC0+6YDt8WDVH8JZUVzcfvIUmEy85xzFRG7d5FyK
GLDcokbBjv5VTY5GIy9MOjgBol7KrDltQPhaMs+RAV0lRX2Eg93jLGCWAMYwqXWyI8J3DWKQu+Td
92Gq6dqImd6aMBbE95eE251VZYREDh/zlyTL54KrZIBfaYXHhHv8m26UUbIMe8lnfttSZQ4zgshf
aNeEGG7/7QOkp9yw3xY+hSXA08lTnuaWxFkym+B+EFT0ZNQwhL3EzHxD87ZBsi2oRk4/msBAFIB3
KbXmpWCvUrXMjo/jyu+T3o5GNbNCAyxTwSR3wbPU3oVYozwPralkt+7lWR74wiHZ09+rzqpEabZQ
SyLA4zceP19jUIKpC8/viSp5VoW2JBS/0tHp+KpzeWWJOkgq3t6lfY5eqvP8CXinK9uKS4XPOpfw
jZ5oBYBEEQnaYQcjvHbE4ZogITApI94h+XStU6wQivAFGr2wtmKDrhEcasISSpPqo6GYWTuC2m7E
urNrSuUN6g/u7qk7d0BBqDah0sM9ayvw/Gom6rc/qJmwwQ8jS/6HUTtjgKoLreqrKnuDVPdQTLhD
Zlb3lvCPi0THC0zFLJ0KDXoVe7WRI21wpVDdyVasOy1kVMwdT6q0KzRFSnqZifqr4K6W82PlxwfN
wM8j1aWBM4+LIfZdAMdB3qf4pZ5o4YqAgBaiCk+pmjJIuE4lFlMh0nko6MquBlV+UDE4rGOCzJ16
1v0Iny1nWI6fY2+yWt5G9O235SnKd9+pBlrONST5KNFeCIj/9vV5w7IhiAYeU+r6HbEfM9GBxgb/
6t2W9o+UsiFNh2LseaKCthrtadhtK5uvJe8G5ZStayuTtKycw4eVAdC+06csxoXmh3TAHsXfNR6W
/JeybEogsZWA/j6RYksImlC9V0pDdmMTtgEUYM6Jj8Ev/FqTtioP8FwYt+mT6u0kvUQPOhRc3Z59
maUnb21ZC2beKY/Qvk0X/fjTrVw5rTMuhR7K0QksaMNC2kwjWfez9C4po8K8TrCcNAntGOEOmnIY
jCJhrUyz5rfObC8SErWYdV51/Hdc/ucKycb7y9EOsM2gU74EDFwGtIhr4x7ly+TJHCiGueTgBlpn
PlVLy/pFsgKLivQmXITJoykuQfeoUBECSUlDKiqR2qKREJ3u3CVdbNwWhGI6tby1afgI0BX2FiwZ
Rwin/T9bTpXQrJ4xIIC5iXfCNEfjMU2BNKfG/04AqGNV/j/jpQSpBXIHYQfiDrIkSwJvOYlHj6Cz
b5lz7MyIX7UsUKpfpFm16iBMf+KjxNyu38rmh5ZuDjzInc4+XzXrONKrC9INkAcXTRnon+DuOr1r
Lcap/Mhxzp3DRvOd74QoLOxE55MIOX/DHXGEeZ0gLVxZ7X8FuKSyXEUWog9pyBOQqUtUTKTVX2x3
cslxFKuomNsHRXx2lqzznOTFLdIjX+GKpV5fpu4KSVdVW+uwK339LQsbyzbNK892f90oZkdPxexO
z7RWcZuF44rYRbvAe8QTObLOpsXLQZzp2N2DiABqsngnAwC1WO0aGxdyuMga8qXLRccm8nztgkHF
X/TDVyjXBoLyfADA35HELUTFVuczrT7CaKAvzzBVk7icrHXsF+hM7kqRHpHicZGTiKPshWfxXBZq
7uepo0Y+bPbUYeUJrYZmEhCPU7pAkCWNVwwInSzq5dQ+Wpmb1hsfJr+24BUCW8/Er5J7ynK9rHWH
SmyuJWBFPbgBYupmxxmthvG6uuRm2RwMcZ2ZAuOfvYzsvcck5FG7DztXnBEtV7ApMQ4U/EhDP+EM
HfgB3mB78TbjShg20N/07Bdk0bqYMkMd/A3v5Qjm4j0EG5ZUNxpvO9XZKi1Bun+Ohu1f84ZUhiZ1
eNeor49b7kMuJaxaSoF4JMkv4wP7xXDrJW74rZT1a3Q2NGSOI623bXrM9hRWcGZ89Paj0IPNLe4C
PNcZ2ztymsLWzz+N6aJPTko9ni7Uvyb+rItEnBUDNeDF7A9YEQy6Ttp1Zhz8+206dB5RtxPjFAeT
KxJeS6nz2CbMNmOH+rtzT9neruLf1H5szD72vENlK7WxYhC3A+Ty7cK4k/4sfSSdI8V51eId5Kwu
tn0JoEz63nlWdqiOKDCzrbUnjrCv5wUWqv+VmkNrNpck6Fyg+cVlcJ1DL11BfNOWi2ilZ5EIqjCb
Gx7rgC913nMUu4pdRj5fSc8ERdKSvBoT2xiDf7FqvCQA2nIny1s7J61EIYNexVFbkwS+IoMCA7PZ
bYq6Cplg5Qdfl9Dnrnd6aiP83mkGGM3+ozWZSspFQNOIf0oXsAHxHd0mrrjxc9inp270yo0A5R6P
EkUmmwYJgcrt2Ax+gGQAUTm2J9eDnThdSGAVcQgqD0jqyohztLpQ+B63ouNYZ2yAU/zqlmLJJPzL
zGwl+3f9P6EavmrnbAlxcUf8DFKCMw6VqUMP4Bm+FxYsC5DPVNmReOhRiMYlPcPbrLgjXmFhlI1r
wogDXBNRBiqX4lkXoumeK3HFYz7ybAYWCQ3qcLyEzmLYPsrVW/Yzu4CxlZqQqc5ZyhV5cN6U343W
gCrF6sRo0sbnGdKGvjbvtvwP2MrExLDAinFqT3PCGeayipzkFUzF5Ex45ESjF7DE2u1+kW27O1f2
VPYtt0tpY/Gzj/tHRr8Wp3PQPMLlS9o9Pbu6Fwde/pfZcTJqiAejwvpwb95dyDA3q2j1coXhEj3k
8ruKsqGPqAzoQbYcxSnV/AZA8R5nlo7BuTMOpvys5DQhg/vLoCVCR2IdeY/qsGq5mvDpFcW5kvv9
muWUAvedCp0qsMkcXwavuZG8i43j7n/rLloAE5dI55InZc/FmXpbbeNsxNJgowETQ5+OsC0uu5T1
OFWw+AHIlP7fIlALZV8TCa0wRyz0KO8U1aNPlIo2mNp/n4mMqS7xenThf/gJReIh/dTBU8E/ccpn
YHca3aZxfLRcHzMOidDG12b6mu1SMH/AF+V5lLxcroQdlhmCt4RZBMEfsPz4kRrlSfz0Tg0a6DPx
WfqtWDuVPwhITVOOc7cTWL1XNfBcHs0MVjzqmNDuc+v0kUcRECI1XWPSU2a7E9PtdICIeUYwcH2Z
cFkQGyOnD42FI4qMuFXiD52dK7SxsvVYXpZt/gZ4fOgNZvsukp2lzDTP1YhkP21XZp5xA5giYYZn
+8K6tKtXvvM7vUkfVCKBLpmKm5o/A1zQwDihgSyj9M77lNDzVnuqnDfXoeykCkVXD+m3GWpDEEis
SZDpD6T/WJbgMHBm3EJhRh5gPljwOEf8xBMV5m+69HFXqxbPhUWWQ2uYhUmHJcx2aVr9opnbd0vY
2jTm4bCkRDoKnc2ftpuv+5eZo6jt2VK7f1eGSQC9WMDDOazuFV1mmm840mkjOCd6QpT4CjwWUlVC
3kCcHrpBY+9fm4RMIhO7Clq7inl6pTdNCnKwxnLw7rHVqEhRgkN1cXH2YWPFWujbxEPyAY7MAJc8
y/Zu2fA7hXor4eFKzBXrfRlNM/I79PiBZkiSvyspMUMEB/x2Zi0FUuO3jgtsCtvnby2pU3goawke
6ZuNuohp3NRP2Z50DL37a/p0xbYt3FkiTINNnsWGaQo6pOU6FlLEm6CyAZ78nUHgyDQBjZSsvPPY
gzw7FpCm14X85jMETbyfpce8cO67vzKLzHOkmmxS2JZ4C2BfS0mERot2mQXlWsPVU7Mg8Zsxxqi7
4zaCCQu2uaRDnBQwlFh7P7BGzAgENr9ysMqTZdNHWr1aB9n0v2PT4twCGzOxEl441bR0qdFhq6h7
kbLBmXN4XqffL/k2ksIMJR70TatBfkHcoaAWSRuQNuMBxKxkqu5hZwXws6zm1A4q4UA7vtU0XOmb
ShZLFEOhiUaL+XhJ8KQHh3tNnDFzkuecT4RaDVELbOvzp1gHsSFRgMJxVrpmwhCjQr1HmNtEYxOO
kIePrzBDG2Egrpy8mCjdBPcCIQbFw3GOcxomI1hRmctodW9FuDRoKZSRVJzdwwanQoSikAVpPvP1
loEjGrRUe3RaEEYpI5ypcqUMh88roA0zr6FkwieDAc8ud/6tSCHQxMgbVjhDeJQUL584wz4Ls9Ee
gt/WHzNh/L2kd9ThHtFMm+w/E0WVDpzluA/0FpEcBea4a2QXIHR1ImJrn2pjxem0vBLIPdgdc+Kg
52uA3gu6r7K99pCr7DA/kcLJxolRB9xv5Qi2OfITrpabzuYrbk5e9AUHCsWMdelk8+zFuvEMfPnY
ctBzfYzD8oW4z1wO8jsCYfaedeKK1fXTFVTHzMj026UPGyNnt7g0z3sOexd3kqdH8nj7RM+RjGr1
5/y3BV2BJGWW2fu7RymoZMO71sgBq6vPHonryQj4h3ye1NnF4y8oETcjLmEtJI0YKG4NzMxR8HuK
tpO3Z46Xlw7mgVQbS1iuG2l70aWJWhi5e1jtn1UB3teZDXujjuW3C6CYyTolvZcvlcj6T0qb+JY+
jCKxKtB00gLRKLx7CMs4mN8sJkCJkZRXr5VVcLwGc5zdWefaYzWdOwKHJEiI8XzJb3hQeMl9MuSs
ZWa4wQNaE05j+F7DeFI5ul6WpT9Ree+wbdELM4FiOdgAoDM9go82YvXJdZEq3I8NpBHdh2GT4hHm
wKZ2uGQRYPzeqMVU/FuZfdMHvIvdodZhQGsUzjJ+gAgKyJmDalO5o7fR5sP8iLF332vyCU33aXZ6
XzJp42jH0oJLqTBfqOqdNpsdQo4lUVizHRUfWaaV9aZ9G0TYAoa2qsGzctGkq9x/sNjCaUU66l7Z
7dIQ9B1yvBSOpT9u7xF2nAz0yeNRu3pJzGj4zaf7yr7Lbr29+Ej9rVLPvKChLEVZUQs0NEw3yzac
KsA+4uFlysF1Wf4wMp0oyj1c0npySNxUc6HGg2Uv1yY9k9LDVMfrBiuwg6IfJVQIBAq79lGxUrf6
94UchTNYCPmtKZxba13jJ5B73b9cGgeltEdd+wnEVTkQgtWJYLCGMQ5+8d1qgRvvQoSLzYy+2TBF
kSB0ldAhFE6zQCaksJKCt7zLnnQuQtHzz/AA8Ef+X96i1Sy5//am7nJg0kKiBUMdWKz8elNEcrf/
yN5lP9y91imTa2CHwsnBUfbXsydFeyEakhIo/UPbK7cQFHRtsmMScVUCwmT3VEI9xnkHAGj4js72
U7hGgMUtkvGMaToSTM3NsosJoZnoS5472SHd9wOgxtW1Z00cf/2kr8fEducVQFZOibpS931nuAak
1a0PbXhQI19DOVdPH/UBWFifDfU/QP5muQt/maikxrolARtQ/Z0+Ksd/vywSpFFZjPd6fuNIyCNV
k0hU0brO9t9e/Eh/mpMK8UdRrZV3lu/5B5vD2222CI72KIXWzcKn7gAnroRzOGZkifTe7KF9GSgA
dJwaYw5Tf4jmAkuqMiTfxgAYgNUVczLrZRtoXqVwj9x6ILimy/xrBYDcK+zPcuAdtfA913KtP9w2
Z/tY0RpeWm2uRczO/vfE4gf1f/hpzIbHLJyungJHxJrUq+n072wCDhbG1LWzq3aoT9Gxg3EO7xfr
ea+BrVb1UpLYRWuGQC4yt7bgJtWXxYaJ7hwNYCpqAte4QwFG1l0L6hBSr6sNuCOmpVtNPCXIylge
1v4/KzaoXjriCklXYV+OJvbm3vKOxF1bnSGJxtqeyiiUqh7joH1Gjp/KgFPzC0/+o/JhaYVKuSTx
nlQJfK+Or4bFU/hDAnESShj+meoTrNW7S0QhDIuE8Mj9mxXl3goOTk8Cac7HrQl/+cz/yxvh2MdQ
Yz//GiJxrDQNpQlXoCONahX3ekheN/n/s1Ou/YvCOYQcEQu+HyoVhdn2ikmHhj9cMqAB0pIT/Fm1
zFnJYHy/m9R90crYqtQc2WYNp0EQ4Sh6EueB7UbbzZE8UxZrPpR8kGFhV4EmTHU0QLCWHYkaDTl8
T5ny4xgnyRF/f7arhSQlgVfW9a/AIk8TzFR3bV8O/Z0mSoi9indzE+8KAZdC0AN8r3jRvm9RUj44
M9uFD1RSqfTLX6+s23z+kwTeUPHE7K7S/bIm+wY7IAUyGakXSbnqWuXEY/cgYT09Kr/uInoxVpHL
5IP3uZRkKYY1E+hNapDFjLsworiDZcPjzq2MFdKsTQIJHFSwew/F2zekddZsfwYnp3Pplg3plPmd
nwdZlGFE9MgTFovvqvqPCii+3VkOQDnuoGhqh5bK9zcUQPZqQZCnVHJYVa622UTy7ufsjvJeSEFC
SeWFd3120Cf9cMnKXqQGF/fLF15wKPIKf8Fr6cwHUGmQ2ZATDNISI8swnrjuYj2NmbUNYx+kImB1
Y15XFpyl5MzHNk6MKvNRqHKWNxwl8t2CE143lJi3qb7kRl7CgMItdXP1GsomGf9ardYYIOAgfslO
cY5o42YOnTzb4su9wkmCspCTdvxiLmDGro1j1QWMhO7c0hiS7L6M+Orpgf7LBIovGVw4NHznPSKQ
+TRgL6mBaKgiqm2n1IkIypLUn5RfP0JCF0qDbALTopxI6pcEmHsru4C1Q0VjbUAkDhkQEjM8jZrp
cjG36ODYmTqbstfh4V1NiTbjqUeXiNkP0JiqNPZ41tR11RwCQb/USahpe6+SuPsK7+2nJdYoMjOk
NIzAKGiSAJ5TvyM9J7vOoFxc5hp3XirmS4tENjV5pzmajpocWn5oij7HQoi2by8aoWDFm3zoR1WU
D1ECkBwVKzMq5Y9Thy46Ci8eoQdBoVaH3rJnblQOl+2t+YfyRxrMHsNCknWM6UWJ0EigQ6lOZyVj
zyyY0hH84n4WAsaCmBHl/EOdC1LienGNrizp7Q+/5u8PnMMglNllJA4V6E5FPRDO0OEwWrp/uwRJ
mXa2Ai16rif/AGxCHsFQ3DUS9IkMGAndXdaQEbhGAWO2jmYWgZlQOTtoBft2neC7DtpO6/1MHCTr
RvJrl17bg++VskbW+M9Z1b+L9bpvdxX6JaVr2zmGiYaZtzmBStaO3gfnVCG4UMxjOPigKwNc2GVd
sGsCZEWS722q724tUK5RV7EMsRCBDtoso6yFfF69l7DHifh7p2uJZTZFx3RgWq5okC5ffCTZOGwl
0S9GG1exkcyTIYv6utuTfzdSZUAVzJAbB05l0eLLcXY/s2KWdS2NoVSIAx6oAcomUDygWz+0/gKA
Wj/pwSU3ozzV1UDWiof54MvTQttEvagAb/TtNzTm6g1F6080Y6ngFh5fQVZwNtfDVDFl+2NB405E
PGjrKUeApg/wWeR6YDOc5savnWpchebThrVeewvk1B1WrEhe0RfiNWEn9OuEjl6cbCmenHLOShmF
tWsidcZqwGcc9tNJI/PTEHLz5R6xQ4ElYDOudH0F2xbk42P3lQcLJ7nTYld1BMSMtaLHf956X7RX
WdrQa36ouNoYbtD1Qm4vUZddq26ewH6H8PJE0TLlOia/kl5K9cW6L4QHww7hmPvaglqD/hQVyVUI
Eh67Vu89weqoqk/0G3rlHYI/t4L7NnKSpsZQ97CXytTQ/MlQzAMbAjISZOIsZLkeD+1hWUbP5vNv
4OrNA8OxttxU8uiC+N/lcZ25bFnir0sp2Y94VY5Aa9LFiiX2H0UC6g4I8gPlOFtPhHCJWopq7V6K
sxlYt0asjaMJORcZJaolErE4hLFTAudjNHks2HtQNyBFXGAEnNemP1Y4c28ElPaA4M/z8zP3sBMb
HvCzjd/UZEOZJR8cOAbPv4kVYb0g/jyVpkH/TZY8vgoPOtYeYyYRLQpvK985DKLjmBmiea+7TqX0
qjIyP6DauxpAJbWd+KVHVfhLACC/5Z+kULb7KUojD0rURSQv57HriywER1I3ywigsQYsELHs3fVs
fUaGlvSnVQFjm4ZxpmA/QwftKTkhsYctADvnfa0MzEERRrxif52IPYXLd2YpM+YKvM7fMgRUr10i
lDYcW+gUrhog6avQcfm4iAuIQ5OqcmTIO9VxGHR3kscFM7X4avj32M494Yk2OnE5HtAEhFOvc/qT
VDdtLdNvQxIGLWZLZvzmhddI2qcxp6QcjzOVL5rFTRZscyclaUwLrHdnUZ/mtsGAOimXg+1xQCUE
1euQ9IQydRkYJn6w8lrsfHanrMtzLpFHuCuzgAZSW0c7u735kWw4jolncpZfPxezrzlZhlG65HYP
uEOgLEkLCoRUUGdkRHt2MlEPEz62MqmdzDg0NIbsUPRr6W2YEuirbnKYLEz4XBUAMbpORGBwaLyH
MMiRzvTrGKMq8Avgur8wWbM6D5MI599yfRbUUEDQEXTO3cuZXbc4I4dNm3MDLAequA5RRynSsEB8
2IMtOJUieUrNpKPm8DKLuB6HAMPqJxS192X62lvD5AoXPfYJSfio2JDKJ2TUlqcqRWKRHn+VYeO4
Pp7cGeRZUlLsBn6rnaZQhDvoL49TNrytfDDUgcX+vPpo1qEpxRt3rRe4MNlIQ1f15y6NVxtSyGNg
hW8VQYozsyIPjA80zTL2LPS1+u/rQmlgHLn2bRypy3Jyx5v2lnpuHXqeO2W9kraSfG6qLSlT1G9L
SVhlduTz8QJ0rVruIpqh4NaqriXcJkA58uavZflTBb3b0fDwoNyApaUTo/K1DBTAIksL/ircnnUX
WUPQW0TdSwoZyMR5w8hqzm0lcwMSQa4hc0ABd24l6n7brQTq95GuIXUW2XQ5rZtL32cmh8fbS+nJ
6f2MDBzPBXoqebXK/ovBqeb8GV8lQMLvuO6IJIy45FPqC/I/utUNeZokV5JiL35URrF8J7n4gvbB
0sKl1YMuByrFdnAVq5nJWgEhh3CsWAzj20CKXWwhXgWIULjWeAR379rtcU9Q58CZgQ+8vKp9QGXa
DzGi15DCpeeNN+GUVw6tkj3132VRulNz2gfkaSR0cZMA8QQATR+I7nEEsknEueAjGuEe89HOs12G
WRr8LKaQBdutWaGmtcG5tGdaQ+UiWZokh0oU/nvHdGExTmOsMxpz8hHFKYaUPkNAYa8aXjXqluFy
Y9zqfpfWvFh/NvXSsQlctVRnQhuP82B2RGB6EZtfr2V86ijwxuoQDbhiLedGxDDy4Fcluaxt392j
it+W2l1ZKN171t5e9cl4NtmXw2NTaqylSq0iIK31AokritYRsUYlfLtwKQyuwCNmG52kcxnn0vxJ
TBYeF/Wo8AwDuzrXvNv+3I1XqrBQNbZdQ3Neuof1viPpTabHKOslITls3gD0lUSNdtasc954hUvU
Wuk5exGq6Y4vuq/vVQqrtjYF2OatV4unmmKcCM7hfHq/uotViuVpAng15i3uNwLRfuhgl03P3UIG
NsNH7V0e2q/qhKXZ1lpzWupsYhkJpMq3SAu02Ir74QiMbpXeEBbFj4yi5dqH8j+5kR714YPLmruS
4xiz1az0OaQWusEu8QaOM3Qgkkp2nfXwvzrlboXMLlV6AHNUJcj/QvAvbURbjzE2iDV7koC7RZes
m0Itn3fIZ/e6jkfq5KBxG+U8mckfc3x2Uxe0cM99ZMEpQMdzLfC/FUDb4+kwsTk9/7PD70rHwK7b
AQRiHyIKiaBoNHgsWp0bszDDbPnd7vYvlOCwADVWnUTCKln6ZMv49IDxTxK8uMg5udJBDikShOdX
tDI7UtTwRdSDjqWApqRNaWufnb9ldAj6w0xhvP/AuzcGi+RiX5Y1lFmptHaOknMQ6oYtt2SAhma5
k/zdnvzjGlgY91M//nXg2GMzK8Gvz0YDPeOwVqqkYetol7d0F+R9quNkkZVMeJ2Bs5T67lPNu4XE
0nl298LXB6hWIhBCFzXmmWg8IpLlcJph24iPy3AhSuyaFD2LCrUdw345cpKNBA2aIgA7fVO5DEuY
MVOLwj9xcZr7uCUluCRcfT6jYpg8/G+AuEpz3WjwZyC+Yb92wRUISc7NAn2zNSWeCoFz+c7suBdF
4NHieyTsCo2uU2vdXCO9BKfw9IX5RpHVV/Dbq0zN9/i87m+82PirpdWGOLWzYVIzPhHQC52cISHm
xkmZMRAVYfBUtjDqw2aZft8fUgZBpBYplPR4OOj5YqHEK673sVb69MzoBB5lO74KLDZj0WBndrUb
zT4BqP6AXq7dlA7WONoq9ofO4z4J2XExV1/R1xk6fdCz9F1Bh/QSsk4LOM2m07T3QEY+yOEX2XpD
uFYgdtW7ARwrHKIR+gRwc1aqvCX0kKggdLo779RZHDZP/FFImXYsSsJ+9sNyj8bhwx2mkJ8HoLfW
mkpSL5jCNaRe0teVcBpvEhXUvb/cI6uwiQUMtQSGxcZdlqnyYqblrwT93mbXgAxKoe50oJN0q7Vz
86YuiuG5Y30KM3JxTSKKV3tQSpCMuTToPFog2Gmdnr8W0CE5CfEZskChK2awmYD0BkJbRoqkOvze
NPzcrBPbNOW5F1af58KUEcuJeTW1kGcX3PqxkS8FBYdr4O4NNFk7NLs4cG5jJBcLmCRPt1c3llxF
JMYlFh6ntpZJo41HpCeFK4QzgZ3xDwqyydHzbyxhClZFra1zX89PPfNkyi1gbNsqdFhb9QE3gl/x
pn3FdqiSMX8L8LWn2wZhiqsJ+FyxaZDRL8fB6gvABnP5VfSlfbtg7qIxNCcMsir4Z4d5uN6P4I5g
6Eedf3WSGR7QgbYpOxt1sf53zSXc1pCEBEsqSTwdmn3TQQIaFW979PQilTyoHa9upoY5Q+y2St+U
lezyxXXyZtaFkKQNsoNYQC8K3rWdC/ij2YyoehxDGf7BxjhL9zzt1GWoob6VZIP1EGmX4AQkQ7vU
IfB2fuj9IVrvsq95xLQa8DGe5yI6Svdd6Z4Ju14fVUX1wx/z0Jqz9JH63H0IGtgiNjW17/E1lh87
s+ccxg1obOls1qgNRK4Rt3ZfT1wX3+7sk51P2ETm9z/0ClPXoeKnZlvVTU9y9PxlO8qPe4Cl57B7
SnC4Z2me7kOjNRex5Ocd6N2lFdFfBp9CL2fOUiYjrlrJlQgbCiFVsXaAFWxzABmUhw4+LjhE2UwM
/+t2+s5LxKWVnh7Kk6F7o7FEj4eTG7D9xeITujTK2m/UMbYO+9pF6gbbmFQRp58TxTk7m+u0PP1a
S4V0URVd/OmMd5EJxs/1Ck4A/B4TsB8414BaN1f6X7Uv5zGWxYHpV/t34aw2T6UUJfw4ISLYy9sK
dQHFaIDJ78KWL5TmubCCAEpMstLcFuecrj9DlnFq6FH8NnkU6CVrTYjVAFfYQgnQxL+A5Q1hnIop
atbBgNp112UE+GJpv1aU57E/qeX64wqgRN119MdpWMYWwgLqVj0R1uWuHyvZODGqdF190RCNpHdl
O7JlfWpH5a3fzrvtjqNs9kq4rXVSReRmtxozGodnKRnRYZOX/8Dnq2xSuonuzQeEOZZwV1UfTB6v
qQkZF4yuGJ9pEOYjoRLkKFHo8oDr7R711w/1X9jJJ0/HRZ8BeLyBQ9MaNt4ErSauSgXk+XBGG5Wq
O0KY5O13LOQJ7gK+hyj5gkxJ/P+GHUuqgibhIkZAgL+KDxSrqaDbpMtiiTJvv9fgqRqrUSThYeI7
q2wnK8fQjlpvvXKIyt2W1hkx1N6xDA+lr1b+R+Y9xaxfaGrQKNPPuFQ1JKjouc9UPJOCDwuD1nyk
kMX+bL90/vlGLvJs3g8bgZsX74/4iKXW+uuIuvF0C8j2WBG1h7Vs1132H7CFeZ59ccaiJQYnD17t
tl0JgSgOkoadWYQt4JztpgNCJGMcTN5io4ovh0YWPC6Mn022tHmibSe1p67uL0GDdq+8kr8geiqq
uLZSxWAj8CFn3aCo6vpZHXLdFJPCLMUYFfrV+Q9qku0+Gckch1dMS77BkbMnVOPaMOGIWFczKHSn
a08e1ZugnTFZGye6EKMAAd429tISA6XJG9iruw/aBje0mnFjX189XNRqVZJQfaApJ1sC7CsHv5fd
dG/IiWcHpoj4Y/zvVHLVWWfvhN5bPWHtmonCSRMznnBoP3cLA3VBncEXOIuvVT3QmPBF8nVvm2QU
Z/lZeEb4NoEabM4krUYBuc4X2fkFcaK4cfmvsEzqLypYZwudRRh7rERyBTHkGfFErmZmE2EUYKSd
Do0ZJTV0yk8oDeBkRZv+pLHxbzIoT0b8Xv7m65pU1xylqpr2WvfUtb+CrRPAxQogrsB1d0bxGHYX
CC+HbI0MVAEcUZ+YMzLlcvJYdsJAWP4pL8cr47mqwx1/r1O4eowMHBqruCg3Q8fcm9zDZT24G4a7
wvCFupeEBNvvfDW2EqDgnnSAOAmxnEo+rj2I67ugEEn5tYYvOaVS2h20NdPQx1ujCVF3QP52ENJY
E43yZEE0A7CoWMiT54oR3CpF/epAYys1UjhKmq123gU5rrr28Vb96uePW2Pfajo4LFFsCrfHp4ip
ieiB4kjmf03xuEDEwiLSp2JmnfSKcwXD0BXh05gk9KfNKTGVWxBObN9SVtCifacdTqtO7bUWYNEO
xnAFBcVP/Rze1r4Ju6SUGznJiSzGVyRpi9zvJoc5KdnIo4tsJ8spYQJxgJEE5dt0mLUXvXsyNKIP
aj3z//2o0ESw1XHZBZtyjBzAGGYoIFweRlwL9mGwzySqYzrOqENoSVL8DESRB0aRg9rnmTy/cKI5
5RHUNeAq/NfaT/n8OvuMh4ko1K02kFFx8HM2YGyFzH4W2FFcQwvTRWBRlc72Z381u1NPjFfr76RS
tKx0dCtF1IC0TO080Vnp3wAqA27+w2l41NaG1hU+3oSWtRQxWlSp0frGJDYNVioqoLA5/5jb+Amw
lFMTWuhUn0cZ60Jl7Raf6yiVHtFzfhd0/tm0I3VESRB/9CkgZlMJszrtcw+/WTGNMHUYt2SjQZUD
7k9MSaZ7uwCAn/Qe57gnkXiN1hnwEgbF/FxQH1r+HlIU0tL08A1VMIWqLyE67yfVFRDBSM7KEe0W
zV9/raOkdjw1+6ekc4dQoQKkrctvyOhmidcza3QKoxvejAvqffmPc3+YWDzeD5Irep6qdbJEdTY+
R9VBdScB2SNQs5dIdz6PSmmnEdILPOgsicJEZqC18pcuinkZWb9pc5ZIsPEsNFtl8YiGUGM4tyiY
i/2ICG57Q2rfLYzLjAg8ylGo/VyVHsPx+PVUdHqACagu/nB/q0eN886qMxsiv+aVmfFlHl/qMuDK
jl5ieBAx/bfqc7S0E1WOkGzcjOhb8f9WJPC/SfbEu01t7vZSgB9RKnQ2PPdA2Yu6PoM/39jGDfgw
nJ3sDkPXWAUCzRBodggbcQfPB6/PxnZWdkaf7/UcaL9axH20C8oTQEWNzO0fNW3Rj/O9Hvqp7ixz
E5/xx1MgcER/viKDsy2m+7eIomfGR4thmwC4sjjSU/N83DRLsu/2a3HJovbhgebi/ZdwjBI36KL7
Iw7RD+Fi1guT+nA3nvCpb8PUID+fiEKJAYd4rbaGe8vZVUi3O1grLYvJy1tcZ5e4Cgx7a80YYMON
H+VBmwKeLNd6lMQb4lEGuqG1y4hdhADtNoP4h+qnPmAAyXxTpCAsoklhvWkq07x1Vri40J652ypH
T++/DXxNP/1jEjyXXEtjLbP6dUSwV6U/Jany4s57Pn/46a0Qe0xZkbN/TJNzUbwXTXlmrtMeExTr
lSk7Ent39+Cxp3Z6urZrJMqpK48jmeGFx79lHDLVzeN+v6iGKKrU/f4oDpm1sBoA/XCRY94SkIPP
8rP6ttW/qaQ7/yM55w95LLFNU0qL3BRnvEDh6Vy+AApn1jCiNZHShdaY/Op4twnaJNWZ0uzXPI+H
iUcEeAgYZzAZs1AMPjuzaMEhPBo0VKeZq94S/+hP4kphxctrxB4xXWDTX9+K9h/sncFhInc54hiD
CGSifFIhuBblVILvSWDkh8JxTHyu0Bre755Q9pShZKQnEdFTsVrvIV3jSv3fZLLzKjb3hOFtmfu3
JHUvGu7FmNw6KyctcDNAAovS/B7+gI/zDirsal0h08SffHETyxT5NP3v8Pnt20HxPAN2TDIbQ+5+
DORB6cQCxskZvMOcuXdIpBfUs/gmKGc3yOonlXUyP7q7Jx3kmGd4g5M9xZUp1Sl7uWNYFgTO3EIQ
vwwYptd1dmtetJrpiUF6QDnSoTxGrQlyLQvlEGMj9QCDPMPyasQkc4RJMj9gqISLCdfTG03iL47E
dZkUqnd5Gu4KzsXmtEU9o8E2zRjWxsDL8OFLKZVCOzeLIXylbaZM6xtsHNYt0k1XIXckGaOeOJwT
9qKepMg0YUKccutCqkqFQTCqhVxcWONrh9suyO/fp6sFRZDJ7/yxh6te4dZlU3CZvJTz6kdGT+1+
kMuzLURXLmrKUUT65YRrnFjDmiI+x5cegheMDFHfXaon/m0+ymkyxfh+HnKSzMMFSPRMW+hnQl7d
wRd86x96C4mE0TEVkDH3BOd2o706dLwzlQ6RkbZnbLw9JtW+NJkqA4fPyq4BmGdt9baED68a5r/f
N0RnmCJctCch83w+rCSsHEDORpvCHqF3cAphwN3o3GYz9aUYJhsYX9xuZh2cKSGKDjXMgdAweTW5
bBo7rn0an9DT3BbpOWLYuL7TQgT8h6WH4DaCpIe2XXVtPphioNceq9kxE67nGR4tgmaYP3pKfNd6
C3+aO057/5XE2WL72L4p5lP1meASC/BgAvaEOiaKmcEaS70bl4z3BwW6YTk6zXMKKrc5Xs9ErCig
cGd5nWo5OjV9yw/nWbq0ZeI/Mowh9/eRy82IwvdmkP7IKdSbq7+YsiRxxx5BiUmlZH/+K2abtTiM
TyBDpG9hxWo3D24QYAf+A4PfbHfAYypB9yKuOuRy74CAYo+PKURmWdVJqPPbIH2Pyt5pwijD6Tl5
PKjkVaEX1Jtj3XBc8tGzrnNcaAnx4MuHu95Hj0h4Z0NP182hX7s9A+vki+fslcFbzf/nU1Uj8Y63
6xi56EL03AJTkNQnAfty6lNomrpZPK0Kpc3cQCpKEaUgiQywUv9TonYBPWwtBYO2uUq3IIt8uvCN
iaELyxXZAxQobJI2GA2/P1OY/2RgDlaMWX2/jisYVoqlfljSRAKKiXL/VrAp+HZflAHWVWH2w5j+
Qv3QJGIPox/q5b7e0szFpqiLME0CiBpGReJChLIKLBod+L1zzE5W2qICVZBnIWxWW8Hg2cElD8yI
wLGANHyu0PIxZX19syyVIgSNL6Ao3QDdZyWqQGWlk48CX/sBQI1Jkc2DatfxkJ3G6kCkmlyu3mxX
4DHAoYDzm6+Sc647drF4qTCKn9yBJMNPJe+tCvRy/QZp8uhW0mDyLxlJNebtDJkmtKrPYFn0G1zp
i6Ccg2hxltGX97wGJx8inpBMW+7xstB+xJZgZCSj3dDpPvTXuoE9z8jxUo05xV0adzISbgQo/24C
jUPG7bDdfkuuHEVDM+u7SfhAcpovLtPOjtjo3f/IHnroX7N8jdaFshN+jnogBDFFoki5PhDjrath
xjSJRd3DuwHKO5UVJmT7zM1GtPstB1nkeMEdJMReOpTtArOW6Lz7Smj3aHR29IM/tImpuFTwtuV6
t2Lxg2mlWXGx+2/Sl2giJIyJYbjBG9jEkDRDB1k5L6y+cqYIkTNNEKxyjncOvTCwbnsOUpNV9kV/
Y3Bdx6t8VTtaqB+FaC1NpuJDuq6lX/kD2J/4sym2DuGgNUx1aeCoBFagGWqWZdaR3wLN6YyGYsHG
3vrOBSQ/wzzEJZpo+ESMCyKRUmUuInvdZoMLvw6fzfk3Uiqjs9dEz7NSot0cuxmqm5wNd3fQLWw7
BV0vKRC1W5CHJorzEVihDz4UL0eU5gK5nW/qi1ledmIfDklWMEFnOVJQ78ZyGT3SqePT/1gb8JMd
hIiFKgREj91pt5r7tLL8pJIq9tAIcfHSIK7eDIdEepNdIejI0VjXOtj+RWeZqVE7WC9U30aWm9r1
qotMbO+zaW5o3LveuLKCpM4DxxorVQ7ppgvGU8LOsK8AGY3/p21ZibXSPQDHgvpyZBjGaYVe7Oyb
N88L5rYoG7GqclCDn6CMFngH7E11cBRQY3er581jQie/grTesHpCjrCTaiazWnYGewZI/w1JKFuD
ASQAFEDA+leNsHQGL5OYF1Y71INdis7LK2z+8GmyiJx/kZ0/Gm+XjOu6NxiRvHqJBrh1Cz0BsV6B
LC4+DtoWyr/kmI3orbLth8XOndicCSTwFu9483FD09qzPijOovJwwRXSjrzddXbZM12Kpal8JgRm
1CawOEKdM5e2h4mnQkiQ2FMjEZE8/cRAw6h0FDXaHST4kWhwqJgyIdVIk1lB6MiGJLipnvfdKXgx
ZuLEFJx7liae9w5tWbnVkGBZB5dKJS/1oa/aJ/A5TXM7iIV5qNcClIRFf/PmhnZN/HgiVzLNoWMz
NygSHE5QROOfr5IAPgLFNnbniuLzfOG00SjN0OV7w05sRsNSVSpgx0nMh0AmakD7UTAQ7kNfX5xu
dckGtxvifca40NxiFFgSS63rrlOTh/2AIZsQHNeRNEtmDWLdTzEWbObMlSq6+bWOGyzHscfkywHr
farQSHIjQIgCBTxKX3PzEjVj6NVRDZm0zYJglNzhz10dZJuhDwrvLRx5CxPJiEgExltO5DISz0Rc
sHzVLRCOnJh8kpm4FMD0gMRtXE/Dm0EPnQANgKeqHypwXIf0/ZEvx3VOaP+mlAGEFNL/e0tLlPnN
61p5PoPJSH9Z53gHWrOFw3eVeGow6TNGO+6NZNgT33VvyHKeD1kPTRI1LdPQY7BvQlwQBd6PYaIW
H6F7L7EEfr/oB8PbdRPxEKfSOzQFZf9y15ilbtIZ21l/VqWGTAcrzec+PrBwVV4BPSMjNWxkp0D/
88eGef9fZy2HnuwzZ0m/Y1w/3JOMDajcnTUvhpv9m5OrwVmJ8JagsXmqcrHZpW7XgZ4c5I2XAI+W
9dksVokeeRmE4inP2hONgmscY+CcP5/zWv0jX9P9aAuKOvWQwv3qT6MRacaEkJFbLXqHEXaydwCt
yWTOO+1/vSJqAEaij/9WCTibadl25O/vii+3JVHj64xLIW03TbQKev8HS7n9zhG6YK3kCcKAPPwV
4XXFA6peU66G2HVe9v4SMotWDPGY3/m75V2Xs6dZVZnmwwqE5eJMbfgs91w2pmWlW9yvbJ6icQRU
B/ruR1oWwYhjsU6fXvFRJBhqlWg4qH41Kamvw4Lo2HwbzZuIQQg9R+3EdJsvsE/7ZnBu0/njGoh8
ov+tiWKzS6dOsIZ98NscJQNAViB6V50w/gOHBu0ci/3TiDHbWluatG/vBwK9x16aAabTQ6Zqr9uO
Iy507BlflgNXLQ/NNuyFOkBfZRMAU5vyU/4z6odgXha8li9tMNSTe3CAXr9GP8IQ6ZDAGkbEBKH7
ISVfa29575TGyEUhVhSbShpDJZF3YU/jrUia6FRv3OkSomGi72b1JWiXf9vLd8Y7to+ha9hQ2571
+MYCnwB7g3bYJnyZ6ChzZ7F2TkuT5lWmD7AoInBiUrCz/PE3+oPtHwIvwh/vGn8V30TKLu5gmNbr
Whh6mzf4XMnpJbjHTc3hNAWVWAu7ugxOMhzDvTMWIgFRKJuTarQpBZAmhJOqWzUVAJql7xaKjjhY
BTE/+YrCejqJDqhqKnkJf5eBzEcnYi7zG33peu0jqTdLm23TvzXulJZZTdj0929PKUCxkozkmUc2
BhWUp0CYaDMglkxTNAzsBvm8uER9QRB2NijqNFZ+CuUlqUA6KuEqnMN4vZqeHPm4Cca1upJ1EMRs
glQu9jjX1X00VYRCD1hEifclf0Co8LMRtgQd75ippIG/4MwftVIW0U9URRUR3341K3sW/2Horhed
g363iGfadjPEsNt5YAJqrBTH+ftFLoKht8XSPX4qdLC4io/6oUpOoa1kK6D+529+TcWyXMFqvOwC
L5fA7u1f2Qjhnkjhjf1EgU/KDMZwTkGouTH5x0WOjbGvCIFTgCRicNLYiijvs8S4hJDKVOLhLk3M
KK9QiDdhvkj3nVeoj9nqkahjTs9tY4hx3IrANRfFry9D7CiRjHY3Tk4PQ3ENV7kLqrO42QkpAhP6
2oq5+nReDu9+L84UuuW6AAS+b/ugGQv1Ya1QDnmlzO+Qg5qSiyTDqyB+wAmMAjiH9Nomsw1dEdoa
T3c2zNOAxMu8p8RVlBJ/qqxyIgTndiEinQoHeVPNvOEDOy/py1T4K5q91SMUKsweVD4QmrBzGVB2
4QwiOPw7+2TYoAsP7S6Zdzcu4YMdu1CTW3uRpGGeedSbyo+JjCYaDngwihwrwis+m2izZdGU1WAa
aUk38PwFhtXFLiH0gSAKFv14MdPQJnG5lYDl8939LGv37YAKZaKJK5cHhZBR3eljaapdBusadhCd
bGCNqdg2FvrtpxDF6sAi7KJy9n/fMuv4/R/UbZQQEWrTEX3YuOhlzpHl8/yYd4ZoPOC1S4eKzHKH
MsPJYApdWVRvRFOk5KyMSUz97CXSCGtOZftXgsVmuonoQM5p3vO9G1VAoUwMFcDTXjZGV6sIApqM
VZ4BYuq0TNx9f5KuK9udWrS9V47QVKa11qn3wHMhu/U6kjTaODhyPVZhlLlrBe/R3gNIXtrR3wqq
iscly4SDUlu5xX1woPK0rFMUZlahmd1NVpkJU0OAfgYXiUGDf0c6Q9pcnPjFXQqmeielDEGJVO+h
lOoRMXvgbLz2VsUwz7xkP3f9eUQYQinDSNspoMqh6zn6ohw2de+qBZ9l2n/6kc1yeddxexrKU7CN
2eGSQv2DBikLDtvucvY7CTpGUCaIZXXv1z1dC1skpFZHBULWGK1tCsDm/b+QpM2zApqAhXTJPAyd
ouF+0XprBLFxDVDv/+Vb6JYrvp1OVhAIgOYfj/C7K8BqKUiTtwEfId07g7Mj83pzQjLkGhSsSIaJ
DgZ28jVD/wfq2t8wEtCHLG4U/7OZWnueCjOIALpDwFj9FtZPU5FtjDbcFLUpr+4eP7GPTsQhEg7W
91QgLYWIV4GUErFZGxOVBfCqeq7MhbAsoi8pNoTUyAZI49Lw/o5bjH9zGwgu2xu2UVco+3ZlABdh
TXPCuaGfoeabE3a8+9/NijUDp+s0aCsfnIwZAdazsax+W6l4ndkG/MEYYZ1YNoFCZNZLaE1VZVuQ
dl/UaEH4IycshQ/yEIG+ISjN9tTCIEDDAiGa2fIpfEfKYNURVkm79uu08HQkJ/DsrnLte84al0k1
0TKOMcktiSVXO5UJtnMU0DVbu3dYCSes3aozNKTcpg8futOEToHRm9Ybl7XlN0+lTXtM4yr2ZQwf
uYlfTec4PnfCqRGr6+wNhfHqP/xa3poVVlb7u/bsLqivuF3etv4Zlh3UYYPEuW2c2LaoYeXZAzAU
PRvIF7yCeL51Watqj/k5CDQCgpUbc3hOeXSi9pGEF72gNjbbdQVriuY6nIf7Y0jAsuovMrDDe0jF
Uv3VWEhRDHgHpwm0VqSkcXwy/IqbdJhYigitELAmRRPbfj8+oWFPi/adtqKAjq4K72qK20Id3dJi
qHUCQNNs8ggDs5O6nn5QzmZh6mxGjysB3tGK9AgZg2PDfH+WtNGDbpC+HtUKRtNm9+Vz6GAu3tZG
lWXR+CG+46DiRhz3K+TbceqxyHx5ldoczcpLIh4lR5JyW4+wsFhPbp6pXBdx5HjZcIAHFk/cwIUA
GZ278U4tGK06ia+NWIhmxC6ZTVU7FJlfOClcxcmenhDcxt8MnbK+5xk/tYwfj0uVx4H99SwB50KX
5wO8VhlqilMIrZsHZDaT5KYc05fHkbMZOAaKOHL0x3iUnPhAEWNsGFOBCDH++IpiFZrh4MnRZvQP
i5DjyLUGO5aAcayT44gmF+tDAaSELB0qbbWUb7sSsaloG8t7nhuL/r4+65PYmR9dNOUJlZKXkXZP
xoXwYNhqp4TqUUPtgv6fR1uA+NKFfS0MerroaRj7p2s+rpMvgWI9PjzKP78arIkbHM5w7cVKMi+9
kWuOlsYudqFZTfYjvmlJiGPQ/PEC+CjBKHYzx7VaCDWuFwnypGT0hT0AWvokDC6lkX2xBV6K/M5o
wfxzn2qmBBCojo9L4EbWum1K46C7j0FV4QWSwwWPYZ49AtUFf2NduzOjDi0tHhLxNFA6mLRjEON8
KvRtiT1Y4i/omAVeLUhNLqNMV9fZEMXCq7674WyBHoMZJHa/mF0nyZAtvEq6TJdLDsbYqgyoQpUo
735elBh95btzSkCywZ4CIuTuN6R8fx7BDnaNgnCLB5ELyn+2y+mqxpw8je+RJAtR3Ql2eN5M5VCH
FtQbYuR8hM7Dv9w3HRytsxCzsE3eJ+VW+wPVOfpUZPT2mKVp8fzbbQU2UkB6wSy/vfax4jFMvIeN
F5XHZASoNR18P7M0uiwImFtjqEINgeDDZO14vRI+snRZisi9OprvZMxBpdwdlZN3nsc2Zuj6rBrW
g+JEROIbdtcatZTkIl4Kh7yG1W5HgRHk87fD4nn1bKBmmguRezxl3hJXGOgIqN9GeGdZ9ypdbkIV
NsobycjpObviaDK+iCgjLKIJRdt9Lzx5cyJNBrhirxIEdpMCnd65nfzrkbB95J2yQ+qBaRSpfzry
797kb6O1dcfFy2oYXjkeK6Pa5XH1yn6Nu45kBmpflSf8Gyr2bjDt6uZiC6upq9WYpa6QahSvLGmm
LLMCZvDP8uBeDRrAMv5r4DD/M7qMVjnTosAThLG4l6J+fY7N1gKtCyve33r3466j7ved15a5F1dJ
iIl1uS7UylP3N6IMyJV9AF2QfOWO4Wq0porvFHjea2jSFVp+jXBqxZg/iQ4/ewE4mVo/yY27Yaak
LW6ABpJXXyvQWe+spAdxFFa4kPCrKEitHgZR4sXQFZbEoQ9/Opz206UJcGWHS8Tvl9Fl15ottNE7
hnjhHPvOeYmHOxrmBOEzAAmBgGYVAytC1pjuOPSY/RprsoN4O/C5ntGzvr/wVUfoUXiJKpcL6Ykw
XRi6pOua2y+lW7c27wSHywqWWuOLtza9f0zmdZo+aCB7UbLMBwEX86P9UfJo4JuoY1gfx/ItjYvm
LPCOJONVkc4UG2LWtLstPvnuKXi427xue9LJh63ON9PbnB+2BKLizQv+zVFJlgCkSZHCJrYUwtJD
/G619f3n+w9KAz/8OxtGoI+k6p2fHjJZ6Fj1iz4ts8ZXBc8lrNrxzvRZwC1LoFCeIEQOgb+u6jDI
p7s4+zo7MCPR9ksGCBxmcuMruzV/N1tOkqnCpOpzfxIJkCP0CBXEQf2bLU3LsR0Ei1BH6n1o+xwt
cJq9GrOAhdrHC5C5CXncoJSpYD9AZZ03LtYEyNkxBoCmpuwDotXPV9rVyJooYH6Ii+5lH+icN1H6
zsO+1Vv6CzkoQ5vlWusyE5Sm81sHnmNMbnccVlGCc6e6qj81mZGRkFZauzdcJd3Pvl2wKEPhXCWy
4Zjm9RBZSHpWKXVj4TxNDfxfuo+hjO1enNgrGNBvhIYdBTfJf2Nu80XuuerWGCa3JxwJK5MNUkD4
fCc/pK1UT0w0z2plSHJ/rNul9nyneHk0SxShn26x0CurLJXiXEaW1bxUPdtHSRyHIOK7SFUrlWIX
4jrrl2sJlLW46TVaKxleeruQxU0WXgoD443Rluvl1wtPJIl8Ojd+6ZgNewWuwpZh7s0lzuK6jeI3
iTa72mMokGBjZG2kTyIkSkVqC0DqOqhh2qWxwZgae2+Zc3AStJ2nU85r0LpI30Bad3/teVP9s5o7
vu09uUaY22Y16Q54UQvRcd2t6zuuxebx/+S7/yyyQtbQg8hOrqQ7OhvstmWCv4kXvdpn+Ouzvijq
qhoEY9wXkCVNMbT2AYGUDeeOau4V3HG652m7pv1TAx/IEI6afRo3gYV1fWHf72UJkNfr/kBJmLOB
1J6/NsLlLgGEBIVrGVup4kVnHCqXLFUbimX/rtrdiDT7TZYcxmoNafoVvcOSt9Vg7s+Kse51Kl0w
AB9MZHnfbsqL8W0KD7Y/L+GaRcl/UmXw6G0NnSkivtw4kaTwfgEv0kkBu9thMMC+wIfCay/6HndN
41O3e0e3JWuY3cQVCfc7HcoZe5FEbOZQpJQYv50FFYIJEhE1EuC9+fZkw36BXMQfwsAktG3gljaJ
PuVTwqDWDOI9nMRMqe13Fn5uw8etIUEInm7PVFBsjI3S9HKqt0SJSFcspSAO6Yh1wjCnQ2kcRPi5
Qwr4NwZzeRhFvPhmyuHcTZD9r4W9vWpRdRuK4fWDlg4eW1x+WKj0tNMgtvArOSNuVe2Ut1kjaFZg
b3K5d/X70hWCsmnU2ONxcokMz32PkWjTkz6j5ksSn6dgddx4RpmmHdSPSqBqImy1MMIJLjyaXeiF
PAPyIvFpK+viIF+6yMQQ+QqbiD/SqrIIr/tof0iqqJiIQvnjmjXTJKdiSuVC3d91xEz5QZsnvOxZ
7vDWp0W6wl32FWLAUJrc3R/ADlX9PmkX95FEgeaG6xX4ZlC+Y2eakEs2hV5dr6WOJBZ1PxFeelIu
vKwMDUcQTQK173HDCTTF0VXX1c5/Hp7ePObY1kc3n3gQj27e/RKPb34y/0WvJv6zLoF6M9EDfAtZ
xMgaTmhjN/SUHvxQW9xgadMPBPwvczqOymcrygXT1t4EPg0N2lnbYTzabhlHdW2RLnuM0OXf5pDH
7bAqLxS+9ikAduYOczM6ReWf4fur2e1bEWiBF8dVwzJP4vI8R+TOhVBr6TH2Dtz/Z5U8+I1iltnB
GrlLtmQdFJz+ijK2uLJOBOt/6V7fHezdw7//RnzJNMM2J59iCxtMU74iN8EK94NRMaPFElK22GiS
KBzurblc4/PEW9Rv+LXb+dLJcruvdd9VuB1l4wm9RJxUdziLqLd//KTO3NIcZl37DI6cqdKxvE35
43zIO3FHaOzjLdZN5IzFGcDeyklMpCXi+EMbRn+YiJ2whExGkSOdavf5aVPnQzUgJS1VGEKXWfmO
Ia3Gaci/1wJaz/ehSqoOKbazO3jFnC6SUCPl0N7T7uVA/WiLZClxZfthPrMCiGVt7IcQCp6PSs1A
rwrMpUg9Ly3NAHgVs76S5ZY5FJi2wPNSR71/+w48ZVLgf2e98Q0RD7mNBUejk5xo9RoioQNPyVoa
8kYcUKw0F4qarktvC9QFZthFmxyHAX71Sw+g+DIWucIyO4NjgkcgNO5cA8/EMSJfy13kTIScbMy7
slFK6eKyA6IjsqiRzSYgeJ2kNwXEK872YssWMddgdn+CFcCUVX6ZpDFXOamrBvGG1MPV8MsWeSgC
qkPSvd2L3MhxAf4T0ChpF0wqOvi1QRMID6x1Dmt4coBf4Z5lWIloiunruU8Bq0a0E9d6QsIEcwJj
QsX756Herp8KI6vgR/DdRAPxl0fL7/IgXMSxwm6DKkFoFQmYOMoDf1WjrgacAJmS+iwVlipQcSgR
G8fIf5DHSNLA+O62lnTjQ9yCGOVoER8LG9w4PJNnspX9Ma/p9lXA0nUk0xZC5GS2JP/D6jGQ80zP
Wg2zLWVdPHA0i1tIoun+bSmrRxqqwrxmx9njoIZwLWjUZMRb3Q6O6q/O6oUbQswwutkqeS4e+Kdp
nanDoHs53F6dwUZpmfnmLM8+VPVwGLlfgE3gaUcVtWA8YAG7ok4kKOyXahDX7sMpEhl2461Sus9f
tLQCOCthA8VZ9MFK0iEbHUuWRVy2oxkcFJojOZid40EXkvSf89guPqa9Txgmu79tiXy+F1TWYLai
vjKS48b3rN6Q0EqHkpI2QhbsH62jD+QaLLMxHzBhvESFkwmDE3yWyrdBMLHSD5ufYpn/isFsdElv
P97xWCFhK5yW0POgM8AmUn5/5ZWbp0HKbDjEonLDMTApvzWleYyvvRfX0X0RcXMMrXTgsFUSd94+
N6PgMyRlkeu1W8c6xKx1lkb4BzREOzKPVncNebgYuJ8fimO48Mqdjj3CFfLgk7X0W0A3gYD85dAj
loZb7TgedVqWWNEMqhX3MvX5Ztfro5Kd0HVpDMXSnVaP2b/9Dx9CWJ/rWaKuY4PYOaKF3yhm9Vg1
P6Hm5440u/YMFzmWJwKchq6OdQe5t+4QhjsAqkD+HfqM98uX2EtpzwdbFy+xdW7GY4374hnx5YoV
DtTqxArmr47sHrSHzittrUtZ7q1UkUVKCYBI4fXQ71p0kqo4hekgcemjKtdFQZwHyW+zqZSL1ccY
9RVcFheVBMUMgQea4+x+3z4jJ6v3YRxUSIcrwACf5Hpj98BMa+B+xo+yDb+gjR9oheis6lSHiTUv
cxj2bUM9FTKatggU7gn8Yta+30Vi/0nZ5Src6nSOy4Sp4h1MOtP4sJrIgkWI6ySncD5e66PV/MuQ
WS0FOYaxabQCO5y1YwDDeZ7WrDTeL6AdLl3a+a8mSdoWfzGBAd+U6LYJTso58i3H/H6G8abgAfyN
gtGGlW+lZM1iAwSNegKR+mv91Af44OkPT0hsal/yIEa3k+aGXNX15uLBh+jqeX2G1wTy/RCKNQy8
yI6DpG4Seerk8rU+WDg+Qvb/WShvdJx4o2q9fDgGrccnPvP9sa+KySQflHBMpPR/+g5LVNZZahnV
7tHawG0cGukBhAJKMGjSFd+VqMLTzSiShtMbI2KO0CL1+gkSbgpFHL7OI+PHYRXAiD9gl2E2+RZv
nlYUwFyE+zbQQSSi+gEn0VtAbV3+qlQKd4rSj7jqPh/Wa6K8ytXetlfGlagRN4fzWBHpmXek0kf8
IZnn3/Yfwg1JroJTcEgvVjzrgAdrWvc0X1kY5CLvgVLetSYJQGHk3+vbJICEykWofq7pApMauKYq
E8y3WKvTHc7WEzfEFR1Pf26xS3NRevuAuM0zy6Gst99X9ZvCwb3uHPSbpT2sRXTHtoHT5kFJ6DKT
82TUmXpbC+j8EfXxOEBvGarIFhBtesuG8wT9YDiEIfjDeFEpieZ+NC39XuSNCAinY7CiliPrixCY
GEUaEZ0lA4i5BQD7BzlVN/1bhvuqYaPlLOt/wRPcjfPGuHjEhL1Objw+TiZp3m4a1uaRBGFbPJzv
gR50tQVgv+vWhh8F8CstsruhmJJ0dvixT7Jon+cSlKyrNPFnq4SseI0O8fN7Z2CzLKfjKg65J1bj
YDqnR2N+LMqz+2V2mLxueKh2139UpeTCNlzVRyj1y28ogc9EvOAdai4fMInuPm9+tW4Vw4g200bS
6MF0YRk6aPI9OC2IBGvF57kn3cXMzBVPh3W5JctsvRLuA2HnQJbvLYuFMAq8B++87Fp2R20VV8uS
fAAUDPu8KWhGjQ9qCNldcj/v8KUEXyf2btMsD2fzcDYRsGyxADLLMqfOxD+Hu9QqdVpB7G6oHny2
gC0+jfbtVbxtqxv4gr/OsTMui/rLYGrVpL+7+uGpNSX1NxJD/AIVALK4XzhC7YzCqCva2GY8cvh5
u0qVvIglgBiBUI/UvBmhW7mRCG/Es0NZjANjOW84IuLf0L95a9mNpGEoFQANhByGpuD24VYIcXfk
xZ9wUYHRXckmY1hR/IWExvuQuEOuzrmBJhXI0dHZTlyZb7dZvxUY3ZQq2LTYGmXTC6+O69nJZMGs
j9fn1vRW1bdRT9A7MlfYmARi6CE4oQsCsp1Nntvf6I0MwaanGDQjUyM+ygXnTOPROkE942qMAX+p
PZnTK60UmGcYcQo5Mt0FzsTzYzkgZcxNe+NGwvbKpkEjQpQeQXtjtqfs4aWk8eeuYUenC0VQDRKs
Cf6DoTEsM9WSGRAF+d1cOP5on7nd5GhvRjeYUlvcwSLglKXUisNRs2i/OE56tL5mRwM3/bgl0qyn
vDa7M8N10e4Xk1ZZlCSxtBIe1gTBkoz8LmuEpVKHNW0+Y1lICjkGM7j4myEGroE1mIo0vZtW29DY
X/3yswotZIY9rDuZvfeEIYUxH7h6+E/aypcHmHB+O/u565r4nCsPwLGVni52bg8NhUp+MFydESoj
rB6Y18+JWn85Kn/tMK4dxDo0Wbi9tI/puxPmnrDHinMA5tvfzmOO4ey961anCFNIttDN8oiWNJnc
IAcUesoF8tYY2gBpJu/Ymr0T21xg6k88XEI3rAgXYEcX1mS0qVkgwkgz4ZwWW/Ul5C08QNi6YaQb
1bNOc9sdhbqOtet6VbLmxNEn35bVgfHFT3GY8tZsckq0pEOfIMbvF9cvsheu9IDwK/2wipVj+XEh
TiGm81qgILCrbO3oLcjMgvWHyFxRuweC3htQUxXT8J76PODJty2KkrdgXOn+jRoYPUKdr7U6hNcF
/xkzT4e08K7SUjwXdi5Ofk7YiKGoUuR4Q5Sx8WkIzdQHopmv/EIKoxjsIIrAh7sNTbQB1b1Yvdr2
Emn1cRW8u2xxT/EJuOifoU32TUeP2cbY8DkrcDGb7WDPWNKP4RedlgDoePczQ011TckqIifNv43B
ZA6Gxd+Y4SIeUD4acaZutL4lfnDeOx4Fq3uMA5Pa4GAa8IC6VnFCSoNG6KAQ6LuAqcjtKCRpF/gG
kvA1ET1/prd7im4mLt35WiDNLWq8ofCqa6FoFgfgEeE0AMBOKAhlSO8Cl/7DEowNgnIZKtAbIT7G
nSDcvc3cCNlw0nLur689HzVR7Uax1n3taUvRLUwwso4ejfHHhyBBdYEKIk6j/swi9wktpZ1vcOxZ
CTRu+byhK0nMo8D6davfDxQPDXoRALwRjdAe2qh4ecAcb8++KJxBVRG5M2fm/JJgUItVDGljVuNo
OzjISGcwGlBcKDNAivQ0U1Cj8KMxdMLLVbiZrzandyJaddv2Rfd63/rY+plgPl8fqyzUriDJrgWq
v+3D3PRSSdChU/86UYlpIPcnzxgWa+xYRNnjY/9LqtTzTQhotVLivAQdx40d9tntjwrw+sXS4UpH
ILK2zdikb6pGIs0HbDs9g0gVCFbgELTz3m18F0YJZQ1j1/xF1gRM+HPggZhOTWmK5Dae27e/xcjL
VWN8rC0DBODYonCbnrtPlk6ymzGWFXz5x6i4hv79Yfzl2vk9as0y9inbub9fLGqa8F3DfUL0t8B1
g0ZsndZQ4xniScxHG4+H9C6bu/87+Ak1t77EPZ0U/AUiHq4EGRv/iVIsV2Gy4W0K2QQGUw39g3zC
F3NxvMVLnNtxsrPfdy0ay/D9RRuyeYNGOchL2kYN7aDj3PQVsPomemXneWZ1s+jzVHvbEfvGfHiE
RZTks2brWsWtPBgTZQKQd30aYNxLBdPdmWRasOdkox6Kc3Zg1kHW9tXQqvqltxVmRQkOkF8uNTQG
k4iSY8zznBv8WjF8rUeCmhc6ArwoF99jEGSDVpqQLLscCyuXyR6D3JQXxY6r9JMXbI57s+XrPGRO
pnUbn1IlpondfNmKfTKOZcf/ZG+4dYDArbLvCsZ0BOeG8qke4L9jsQ7ASJmLOsenkixFbFaSsAHg
b546EWbzYr7CytMOck4bq43E5xwe71g5svBiMVW+cmUaLsFpsFPISCK2cdSfHpoBpsf8j5kQfF8a
V6BsTXiIsKBu66ukIQZl9FU2eYRKcjE47XGbUz1hZyWzJ0R92zEoLVJF3z0SSQQ2Bkl8uT1Df5Sy
MhTt5bT+oQ9/8hlWbU0jSAqakdg8oCBGZgWjz4L/4E8zfi7GIvCDEOctpY8VCKM5nHVPRrJeLhnC
EF+fIaNDtDKCsMm+u+9JR4VpqVQrrYXd+LDjXsLIbCCU2kNHDIjpkaOad8Im4Ss8xhohjqxqcExP
DRzu3h1r3usqfSwjl68xuiK7CWZOZMp+oyKEaTPQ2MCrINdadMDu+TnoF+fnDno7g4ejsr3TcPL7
R+c6svVyci1UTX3bNIvFBx9bGX1VlTaxUrpqKiLIY582jHaAU0kF9fmSN6g/GjHIWYdCSco+Unbc
gEx1E1bZkJMTLxQQP07EGNl1KzLCR/cm/A5wR/x0YMbv/jinRwy8Pe2vWB++0Sx9Ci+QFL3TMSXw
dDLuGmuG4hPN8kj8sApkfaChwWbDE+nVWxHh/QnOc7KLRVPzg2MK31ewVACpS7C/3xoBY794g507
ASOJ/bvkn++Y1DFhEOUgqAaOqtYxHj8nwfe7cbhVNRQoQ9tqbfsWulMo7egDt4HR2KNPRrztHtB6
fjxZ7NocuFXdV0DBThjVkj2ld20LuRgz0o4oUpU51/2ikyvnREU8/y6YM2uqD4neCUyAUcJnsssp
5PX0XpEAPZEb/W48JdI9IfMX9xdEh/YmJ/tACAQPtd8gZyberii6DoZcfb/6swseH5bpI4rjwrwO
vmd179bN5UHYOt7KV3GU84lzuVr+5B9cFt+hScTrMkxmfLA/Smvdpmom1fN7kWFSMSaUdsATIDIc
T+yToxD1hLWFkz+nzwt7eSJ7u48bQ1wpk7cPh/xJQJ1en14f2V27JmqLLsZ/q8JUBwSIjOetivUa
UepiEO5gOs55gycoHlsJputU6+Frr1QV0s/072bMV/sH5hHe6+LxJd2BwNt4YUowJZd9WnKgaDqI
hT711/vsrJSweeuuMHNsjPxQUxN7oxIB4xwDbFxv0/fLVPHqAEtp490/lNTfEEcAa7y51AdJnshI
J+jwWUn/w/er91C94ewlXkyV9v+PnCHVtx9B/2bZ8JHp6puTC4rnBC1b/UrQvOTbNrMvr/STA5q+
wC8IvaEJg2VuFKDjJ5r9avQ6pcVO0cDFfNOFm3ZiR0TcZnMcVxgDpN20BUpa7SQBjBOUbrRcNXeo
o09OyH7CYK9wZP9/284FUJY4V3oILxmIxcS1TYfgPVNYp68L7zuskHqIgGtE6bdhTIC+Cx8uUyRO
OBLv20hzFg6uUSZrVqub/DFkC7WSAanDu1E2ylrUWgyUkLIoxChwtxMAM/nEb5A/9sRaLxJpR1PU
/sOZ0ckZlI70nA2x52dLXo1i8eH7k7hDk+YFjzLOjUw2YqtstbIMCtjJuwpxKOWqlo3e3+NVYwm/
Ga8EBNy7hDOtUm1KWJcgaOiI5UZnm4pLuVXv2o8FBz4MfxRoI5ajo6BbxALQWn1dVbmI7AunjOBy
OfDpiKMhkeZQK41ve5cKh4YRXWAoZ5tE1zvDbw6vEN7O71idboWpTvq4MjykXt+55bL4MItFmIAd
+vrZ5OY5L7jYI5w383hDewPE9dzUfyRE8vdktEX8tn01qr2TmHQ7ldrHs/Wsz3FGvqVhzYJIEdmb
h+ikWUTlYFwHgouSPP911mn9BJ33Vs6/VfrbNztAe7dws1nFt2HBEIlRXyJz5ls0XSYJb308KiDT
cD9fG92eqdS6pVjspwwrgth5SLul6sa6ayd/vxur0dYCT9mj5dZma+EtLLDNs91BMv4DZdDD/Ti1
Vm8FdmwHKFLPFA6I+tulfrE0z608BHotTYsE18vyiDsIxspfk9G4jaiUeatZpWNU7KUrOcr0DUSm
R0CRQpKRyS/AJ57CvG5XaithbgFAR8NkME1l4awaYToF6OxOqH6IUf+ztHc1LVxcOeFSKFxgEPlU
9Uf6gKVyo4jPn9azU5cqXTkYA79UdNVnf+CoLJ1kTJMWPg7vDiFBSyCO2HJAtSShddygcj0pq2LA
TmWa0bxzCiiSD1XglRk2oho7L3yuzXugglNjbERlc/Jc96YAwFGfYCuffa/mOev1c4pYzQLYkq2o
120sOV0ExXs2rzLBXLRSob/oRZ6WSvXHqN3UP6s/ZPaQugej1vL+Ckmt0LRv4AFQWj3YmCeZ5lDM
bshLU8ORETRISqd8SVYVAE+I8sBr65p3YCW7DAviWwE5C1eM2LD/zaCE6ZS4k0DV4iobnzvjtuX6
751FW98JmZ/EdIzYo7WwX0U+Oi0FVKE2BHcTUlMtD2EsWiGo6BtEmiQD0J2NgJsl1L1Ac58vq7Z6
/62wGYP6RaWjDW6tFLCAp03BB+qlmQsuHm/jxa89SiT9xV++bRHUByPvnabPoD4LXfvHGa+AOuwx
g0R+6smXyR/PFQeqXpj2bnbRVZfXMwhLwyNf3+gGHe/8IhNGWGBnFvU+6jr0T/sQdcTij+u+lWpt
7Ct92WfyHR5GK1hZ2Cz17vkWXKM0cHnZDKFWcQfRElx4zMVks1eaKk562RoiExogNUSx4paZ0Zs0
EjtV0HyUi1rN0ksDMrkuiPhORTdugiFUZDI43ag4sSIadlqvRer31ih1Va9P45MPpDjyzHIVVv7K
ZeOYHAjIvqulVqy9NFEMpyB71Lvu3n/8H2bX12KPKAT1Fa2RIRZO27p7S6/cOHUBvqtUbPwTpP2X
N0cgDB1L4UEzZvSl8xcs9iZqp7sIP+Ye6iaYfpjhhT6IM1ztbbni3U2OlT8xQaKd0Lk0hI8ZH+ZS
JTVoh5O7syKmco/xIcqF7vryfnERz1ONMlOAFCrfvKu9jQjXHK82YVg1P3k4vYtgUBp0WJG2YZ2S
XG3o1Fy9ohzXxBZrWXc/yIubob/iLTJBezuhVM0fGRNl/z7aS3auE5QqyUVswnbDp9stk3WvyHqy
ucZ7agT3m79PjUXmVDCKjz1Gq0zqo1EUkchMKfrlJxuo6d2vB6IQBR7A3BLbPMR8VNi1PpRA2AT3
wMVjPWCEa9ZvkLN4/kb1FQEgvvq+GTL1KyBgU6yiyi9HBm0lMZfRcV7J1/MkL+q5EeZI8ldhe4Fe
a7lcr2718JB+KtfZx3yXNzLNBNPDIx5vP2ENLh54YIDgw+Q+YxGmWM2PgoVMs3mJ1pl9m1LZ3aFn
ui9fCU3QZCjID3kS5UXGU5q/838Ane9BoR8A0K6T5+d6tc/E7mf4RY78HG5nueMk/j3MUClOc3d3
i69Jc+JaVzL3fG+bLrTy7D3XPyO/lc9y4x/zpkdOQ77V0i8IaYpE5RmDBc5z62cyJKy6j+Dl9TUt
8UA4KMgTEVnehdMbUOLMCnxFQbE0oyZrQqOourMoh8xS9Zn9+/xKM90MSdWs5XECEAYpZWJEZ346
7AwTy+oPLJHh83Fw5/Z/sgiZpzROvL7vobyMresc5HLzpTMyHIFbA/+N+nxC/Zrnm9vmsorfekSj
OEJ0z+Swu3T+WmBYFnnYZjj4DSAPM/8SYrcwf0FeEXiEruvo7s+uVi5EfsJ09weSfq9qdlGTzADK
J6Efh7jR9696GFIqRyIGbfqXXIzGDFMHVvyGJQrMa4/N1uKhH+IrE5Bv70HGjjifLulM8voTmkjr
8BNwuU3empZ23v9OAguLt8q+IFTb1S6NIszUjlRydmGK1JwdQ5XR54STpzcQ2gdGhw0VsDLXFpY4
eujFBk+TSzsB6hVpe75zPGoaCakmZkaxEaHbGJ1pElhossNknjd1Yd1xGAp4diCH6u4eEZOaT+xV
yXeVzvZC0wCdlPaS86adB6uTUw9Gi/vW1x3+cU/IFGpXOFnjLbeo0P7mAJsmCOXEwUIQaZ3qI8h/
8VBWpAkR439NrqIN8PZb/Rwg9l2zOKmnoWcwNXKKBaqM64XHi9t7Cxs2Qsa3+TI6yN6Ltmd3M/rD
U14vEJ2JNFmXm1qKjaINxsq3iu3AILlpbqyKsCblULYU1ba9eopSY/quQDKRCKyEFT8XZdhEN1JE
kQIVp9yhPE/pj4z9ovr/yTpM0g6mxU4Jt5wIoSlD8tjuWVasNgYQ9Lac9AcyEp1ArNxNvn4SYlOe
ITvZCMzdj6IKQAn5h79LUmax5g6Hc2uHkkzwV33qEasvfup/kv+KcyyXuIWLk+uf37N6pfB5ZetZ
7j0s8LWsT8KH9dNDehcXvc3MA26PQcjr+fyR83Bq65VniHtuZIbVKCOq1BLM00a3G6YmrS5Btes/
p9q+vlj8YCBJFbTI9YgU1ttKL9JMlZjBqZYSytWOZ5gmpFxsH9GPUIPjWc+Cg7wTkSTegGxExa6o
JYH9vljL45Z/7JT7jn6gFQSmSqftR5AEaaxcG+BE8PeblxThP/ZMDLoIVonus+Kj4mIIMk31nqii
Sjd8psFfGVM/DqZ4H6s/kZKxSivoUQ6xlqhTSuxI3i/Vaw6GrFa8E98nua6jgD07fghmc1fyIimX
DQbmHJcIt4zIzN1092XP+lKTsKlTVnjwRbhAobgAqINnMRorNy5v4lrLRgII2d0nepSmF6i5aBOT
6R7ciWMwDjBYWwcDNjCwHQbUC4+/mJfxagE5WXa6pnHKxQRTsbTDJXcZWCkgai5EJtxZum0DPKuc
Jntjy8guJ6zI6d8EQfvpIC/y7RN7F4jCw2CQVld3w4lTTbU0sbtD5KlnOR/7xcIP58WPe0o5gG2m
nO3seYOQc1Bn4q8Wd26yLxf/jbCjZ9MVvAfKtYUsHdyRuSGV8rrwdpvNPOuUTHm3cj9GSWkHm1AL
RFZ4PDJ/4obG0vNWGrqieAv/MlvBQl+TM/UlQKtLUd1T6Yq2aT/Eg6jcSotzmUpHmQ60ww2M9MUx
kxEcvSJ1gRRAp3S3yuuJU3ZrLOIfIy2PThiqmAZHM62C8MEupcz2FWgxbRI9buHyNSnC9PtGVphl
Fb8jwmeEOp46xVlY4kfJQ9TtvtQ5M91zst5WyNS5oOP65mOFQ4mtclBOpTMhjBIoNKlN33/L1wkx
wFcxeCrbmQR9lyANiq9/M6ScJFmERfbU1E8XDfSosdIlWz/tmpB9BznbysJ7C6gltQqRlR9Hrbqg
bAmR+DLj6rimDar+MlKARvaINGemZ8kZZJxfCbulXx4R+nbKpBxC6ar24eLDiN2gC9j6KmSS75GJ
5aQUwfH4HuoH9VC4Vk9k2NTl1KRN3zQ23xry+TQoMtp87cDVxcqciOni0Bhkp9zcNbFfiiSsjuDv
Lg2ies2HArVcpsGTreqAp8zXh8Bd9YwAG4iyB6Kjg9gp+yTu66vooR7uCtEn7/KnVIZNr5AToFOG
v2M3Bi7F+7zWSwpuHWqHovTFMPPd/9/FyPcS4pLGJM3FC/NUF2CGYLqSUwhq7lxZAugN54nF7+Bg
HPFodw96ozkUXBe9NWhMW8RrM263C2hHHnb8lKr8bQR8ArXku8v901IOsUvbfgXLnRe+L8+LS+3x
U/JUQS3PWrtOVL+ktNbifrmcBUMfJVLZ04dKS7UcMcwtLHwzal91Yxzv8CJyLNzNnU5fnDMNnoWS
F3sLISo2uw2e4KiTllITApwnNFJLruf21KGc7c60BwS1OZH+gZyZiMECW2vJ88Dvf/DLQcr1p1bt
C26gCdyHSK6PRSeTq36PGYMZpFXTFREWoVZCW6zwCJ4V7QiB0CTSqzVFZ+UNVIUbZqQ9dGPuORGS
x4rq0hHHRynasSVoqSyl31p893TWRBg0agcng+T2W0A1dR2yxcg4fJSSo3NYol8u4EY8Ymv0GO7q
wQRrouoc9+9Fg+shceNpYjuBXc5rKjY4Ju5gygNoUDOPp1HUskxRlVG505CNQwyr3bD8yKFrHqPj
24qTrGLfoATLRU7qksryyIQz1cr/dJz+Cp9vrPt1CxvSX5Rz6ToFx9nwFp0E0B1mMlk45wd33iTm
604YyJGenaA96zduosvP4QpluK9IZqNPSpiRximbH1cIUzTLTcgkGnBZqPXYKaRl0zO4qpf7OaJd
gl3GlLga1qidqNVwXriIfOs+LevdxincKqK8UBcgxu+Blm2dVqjGxTYLyLsaOF6oh1gsNRXQwf/U
wDlEYdXwyS812WTLANHvW7ZBsahKi2ni8IKQCH82PRLSwjjsuDrhiPiUdMbT1RoG1POYEviu0DKM
I7pP3bI/6YFJSNVW4pK9VuMO6nwpxfWEGEAMYFUKcJm1bzHAm4X+5Esxvi84Fb+ABPwswoi1FY/1
t0827LXEr92ldNhzuc0T/lDCNKBMBMOQlMMOJiD6gCW1/SbSY0jppHTE+tGOp7HKMzsbO+fIEp1x
Q2+9Bc3fnAamUO2w2SBU7I4v9jar/FbO6UEgPjBr5htxBK9PngM7fse8xBYsN1WdssaHLf3+ZEcb
R6wDdynnXIeQJ6XHUEA6UfytpBUfoDBFCCKrQ/l6F/pMXfGGhZFRfT72y6PAlXG306h/M4xP3Oat
x8Tp2yN/vcW4+gaq3Hspb7s4zHJIKV+Pese1Qt1Bt223CeNTYYh2diSFx7vQVbCHZiaWbkLDjV57
CStAlFNRXYZKtxkrr9AG/zR/1LnKg3+Tz0ECzJsHg5gLxh3vHuKWX+WJBnzR/0AveFJeRGFXXmJz
YvHtzuCHCIXUsKD3IZUmSW8x8pQuiRyKB7Rp5pZm5j5w+EtSdxWCzM2bdV0Cu1e0RHDpE2EkpIPO
zOAwOcPJH+hleQp/0xN+4XIrzP+5EyNHV9puBxiCTGMveSGzeSMEx3vZGzJgEnpHerGQk2XrP3Ow
QNLO5t6QafpFo91nOOmwKTWD+vgcm26Ey11XfKYTxquk2SdXHnvezUCKTZ9HgwygWE3R2frm2+LV
K3DwprfDcjHxbOTNNaJh31YBtXJoR+GHLE/N1k2IPTxDpvXRerkJn2KiGLBAYL4EhR8aBw70O8eD
dcYw+clyMnm6NCBdiZW3KHlKlm8Vic1rsbmYfQYYThh8xP18Vb+iYCjPaKHtnWsIyehYtn7r4cb3
BFn6FNPGjfMDDejJBJHPBc28r30vKle3SlKAk+yupWP7bbkIp729Qa2suGdFxoqe+9DgtW+8eDAi
JlLg8cFA+Z58vZKM5RCTjHSzfwN7oGP3sUfVaIExpk2RTItUwoV5WAyUORSX5YLHIJ0EUss66m+m
JvjbdcHK7DEZFpXrWbHFjTuN47NODwIRymGFFZRRt9HM7rH3dlUuFYxlxnTlFYSOnLfsSY3JLdR2
fq1Y9c5LB9XRbHT136nKuLXqfBJhvh/Fcc8TCg2WHDoKNl2U/9rDdoH5uoC09/6dSXHLm1h96G9U
+gF9uu332RSbkNDqrGw5S7lGePEV/kTGeT/bZ4EMmJA1X8/r08KDzj4XMv/soMzk5el+0em1gYYz
LuG2NEKxT7tDwJBruno6ihc6w2BBX1E63w4ly0Q0rTkXx2TPcfjC5Lvtad9sQK+Ys079Pnme7k9Z
6EyCQrg5djHPwIZJsFbYsI2qfSNBIX/8h3bxNkIdiN/AJjyz/c0mz7Z4XScQEIyeSU7B97HAjUzW
yIUF8+4fWzy7Hq8v+ChQ1SQURIjGmGK6Jj8cFVVHZU1zPqlu7TR2cOOtiV+FcF5jvVnpf3HGyqFD
B2yaDia4tVpRSyxEOPgRDG9/27tJ8J8oON2m7e31pqp8Ahm9hwgrrKVgO5rJjZckfBBHEo+K068o
XNyzIbTP4ipnCR5wn0ZGCUnR7gU37n2zmIyDnWDyrvKyNhrVwRZ2Nro6nk94kf2pIPe2l9xtYq1p
8pJWh0RN014rCeDQ9DmGn/VHkpstfPKKwnn6kJN4/OQUH+obOHmkUxjWP+6ANmfXSKUvOblPcsOY
aTiAGu6L3z/Ep7bCcKR47TMTqdT0AlBCgzflmLjU3IpgLnQk3FZChtwG0d0yzStzOpr45bsEaEeB
N2it7+v+kdu4P6WMYmUjRquTs/GPtJp5Zpys+6MhxbrwBqtbFaX4x6a9GQYNUE0xK0aJv04QL9Y9
b+wGpvRslSMeeeSgu19UZLNUYhxzecACaZ2M2PjXB/8GrJaFPMvQitTcA5nhuSMA8dDNru/xD2n1
blbN383YfK1OQloAaeG2NVTO1tWErJWoOPpYKBSebUXMO/X1W8qeyeQADknQjqBAqelbxeNiIket
b1i9t5hhtKBKFGxm0SNdJY4r9FpsVFU4ZBQHzR3EuDl6Dj5OgEheqUcuxii4ngrDko5pNt1k7vS2
TAv4xE/eBeIP9XxYHKMKsrsum83s59AnsYhvrmWMbP2ryO7lHxe6MikmyV5Y+5cxZ7pFAwnYWT+E
utMDtMDTD5NEsSIAbe8lhUUW6/MOkKEKgs/k0bfuArhbVaHUvNmunlMFsMh9kdQzzA5gQtKEraoq
wXErerJM5I+6V8oowYma7uxfGqNpnBtLlMCCougtw/igwxWj4nLNVnyeXiIPanUhGwmXphxV9XcX
on9/3DWuHTWMUdWbwhUVxspmNwmdpiWsGiJzomtBHN6+s2ygkakVc6QMHa4RWosPX/R5VNR79a5G
egGEAaC2rCaqaLoTjnc5l7UoXSxPsFv4iXV2VmIwdhpASO24MQYDs0otUQqJyGvIzUoBaxeS4mcv
CufViv4jKu4f+5nWHHxSdWKPkoCzblPqWVqEw/QEi5MpbA/8CwsRuWs6vjFt2hmeOl+ajnFV6zrB
Q7Y/D9BJthJyuuLHYfCxsdnxMHWDh2XDhK2ZCvVjRs07AL5nn/uMhpWxaFt+LGKRGUtu2PgsEtfI
s3rSLrilIu+gl3Jpb7mxKLe9+uEZt6ajKtpVQSy4oaD8eXhH8lERKWaQoZjoUVTDpdIwCtaRsUDt
0s75MLdlNgojAuX1G/vh6xVHRTvCPewHKGnLKg71uB8/yS8dRdkE68VuBK1vOrMMqJEL9nyHwgT1
JQskVBNjpPvx8Q9kuk1CCtJtuLsCQHxHzX05rHggqevkPw5Ih+REGjz7QzJOd3GUBWnZpKktqSvu
FRezz5OaHYC54hHfTisSkjdUSzP7/fldhB0RhmjV8UFh13fSuqPR59B8MqDu/SAVgfNFP4UGjfUn
s1m4cC1iCaaqS5SEw1lxvOtum+w4XoWm+4m27S8d+WMlVyEJ3iF8t8xpUEQcfY8wwO4wf2koKSjA
q4ByXQq7RH1QtdMiL+3yClCPXmXc0hVxdY9YA3qQ5Pkno1k6t2TseUPW/RQQTGmUgpQERR8R6W4M
7l/B/Vcg2lQrpVnRwlMl7gBd7dFg8TGa0H8LydeVce/1I234H8y2p6mKmHGL6tkqla1tP2UL3Kw/
XTj0hGD6Z9NIU9z/WpC6qryReMtyRMzMre0I3PuNDRoY181J6lFu1OFIGm/VczwA2O5Sz7RduLn/
l6DTE6MWSSf83pZfbLx1vV3YiB06AXfImLiVRsT7Eee78J/KFfoDwFrqxXdq/TiGQD7C/liaqYYa
qfPXy7B8wiTGmOhbbSq+Roqe2hxQqQ1vF3AGQkSdomKwO3t8d1Ne9ZUpjfoIH1HpVP/1K+2zEY7y
Q7k3z73+i7L01glWeyn7IbccOAL76nuB8XSn7ml6NIksQa+ZnPu5OGUh4M3xC7F2Sqdyiq7qtTF9
piLoFbZxrarqSoVQTOn9gxQ4+gV/wPBmAeBZHq64KbnRKDkpwzrUsC64eg2yPsZXTMjONhV4G17S
sVLPpqu90xU8X5Nvow4i3xUCxUHfqXnTQl1O1pA3KY5o0H8WBowa3u9xvG5qTMP4d7yzp0YcyMEP
GglT/obhenWUT1qJY/iPJzVEMhWbsnB8Xlgaf1hPZ3evz0J2K2Bv4od59xPLbVY5Ko2gCYaMZQlZ
4MJzX0ElrozOHJzMwCHS4ikjxjf2Lwj7dIkY29jhfhAa+SL0mhegkBbZ4gcK3G1vBZV0DHmvWy+L
1bbN//Qh19srNrlsRZNQa7vWoleziAED+YA6w7ifNbyYUXf3gHfnFoqPctsIeP5NLvrCqHMiVVS8
E+O6QrGe/Clp1PUA4dqkLEzOhW/i48vqefFoUQDhT/voy+84ygHvhzwyVtAwhJ7xCkktncR0/N+6
b8a4/43KfsMCrsP24lOlVf6mYDAOSHE3c8yP04SfcKd1JZ2bbeAHyztzmNJ3qyjqu2Gx/+FvvG1X
RnEpBnv0qH86vSw5I/f5Mn7TwimBDZZM8DqozbW0U/T3sq9IpgoYIO9k9e6/rU81MgnliBNBTpnK
rBWXD1uT5u5V++ZnujzAPit/nuZFHbvG5Gd4OuZCajk9LcxwJXircvTjLc+RN9wsqUpQi4x5JHWr
bGs9l+KlOhLVTi8ZMiIIhq4YRaigF2yQBY5XpzWXpOL1/Qx4QTkyyh+LxVCB8w/7ZNf1K7VclQQ0
DW05+lR9y4cXIjFaX1EpS5TAlqcrNUj2YuQeSzZZ6/drk41iV0jrsZiA/H+0cxNanIjfX2wV87SU
pwMOVZrBgBujn3cPs2gFaia1HBFdnGRPDY85eSEhdPJbPZGFHu4+04qIpX4v0INs59lPqIKs6Ipo
fbKWSudO/LDB6vF2OAFkJum5nHB9qPCUEhVwF3Z5SsFpx1jtpgKuM3KG6z2gBD0jLNl6NHIWGu/A
WEI2N2UbMFwns+nZR9+xzlYqBxqpYKNMoOo6ew34ZK1DbsP0beXTZSHvI2H7KYV0HBowpUuxo0e4
pT0qBg4rU+xKNcOdi8akc49zkx6dxq9geefplukeKezXfS5KlwSLDptBnYwgHS2iHkVYeB0GD/XJ
dGnQJbFzR1JnlhsDnZwDVm0zdvQqEIQs96mry0iUSZOzW/goUHJgMAqtuvhPU7a9LMeWVWC31kD3
XG+IxFKM9J4SQG4rWbGyt2rncxYlZsNxcWihzGRl6JNJZoasXutBPkBh6CihTIZ/DcPQmFKm0G0E
cDgtNwK2i/MAeyz42PU3NK+9EiwzZiTgzWw7RPKod6GeV+DXpDtd5XN/qZ0f9rJWDdIYEwD4cQRT
0wJHY+G7/MnzqnIUI1fY7ICMUCcMwLAwNkcmGBH2WgDn0JgdXahY1MVOolxJSH7l28hRIUy8e1gL
U2nhyUkdYi/uQJJycWKXcxsHaVL3rdh5PR8ZhFXqwc/QH38DNMor18rhSJYwd41e6bg7PaOfyYBo
uD7j3QDpqdh6cDd0BTzUBv/5CE3X0i0RYEgKpi5O8QCWFzdTPEv7t7pEFAahZc2lPESx7Rql7GAS
IRCd02VwB6EWdC4iL/uNyJ7Zpt3QSlq7r+B4DF05igjuBKzuxjIyJGw6+05Ek9J1HbkCLgbYW3jM
NksdqHf4uPtg1dhFWPnjHWR84EE857tK5gIyDPUlhI3ATjQNvYXg8wb6jkz2GPXS/HCXtTCKtwyJ
IztOtmNMuYHtv1sGTYWcyYATvuAUPGC9xXggGcNFYEMNgvagyf/JoR4e0R+eYfPxUTlQuMvqLcwt
7SHrCkhJ2FvCOD/SyAVzEyLPOTXS4Tj4wpnSoVDOixji9PWTr1U7bSC9sExcKZrwD3E8lNPSM97+
aM7o0RJgmZGqrVXg3hORqprj9cuV1cKcvAM66XZ1ntZEIJEgYsZ5RQyFEqTBA65LIKjhHQtpkRCe
WpLY+Ut83K+CVV9yg6nT2TYus3DAk6wh0MHeTokoc1sMukJJB3/lDBi7Omxv/B5dYCcxjqUnpqWz
mV4ip6NK3rIBiw3uLlEITNds4VnqzU5CSFTWHp3xemC+R+7yntTW3s4FOlRvi3Hz9fQ45jOZwb/P
0fI79BjV4VozVCovrAWccyqomekBUSr2LArkgMVr86WBFTI+3OZab7NjdbQLo5XcuJmLTIiSIycJ
I3QI2YJKreWPzuXegNBz2euxYuCKvPOj6RUdGyjBVo3v7SkGfXamWGVsCR7n2wILVK6lHhwDm8IL
3B63Nd7C6id4VkxVnoMolrv3Tsybi3OR/rVKAmfTLmHAl10D4Ipf0q9p0mkVqu9r/fCzeLDoGVEj
3hi5gIjYPOyETSNQ3kCnoFO5xX6sWu9iCLbTBJ2MrfI7yDpFwU80HweTLHVKbCjy4G/QmjNHV5pV
BSp4DeSOIfY8kdAIA2UujeehfcY4agKwgWSsxq93+Yzfz3D7imTRXcdcRZOc7nHiPzzpglMI7BqH
c+y2jbRZj7D10ZElb2aQfun4ascVGVqSusRAvy2gaju1BWqhaWXIOHZD/CXdHxQAbZYJe7uubG+3
0XcYf3xe7JvHvolHp1Vgh4xNk/1iMLb4AsNJJpsnlIbRcAMSW4GFkido2mLS5u8IH3VqRYlMHY4S
vlR554TI7srNwQvmHGWeytkwRN7NJ7nJqjTUqO9c6bvuwpLQqO3b2KZy8GQkFdXk28pZ8U0I0suY
CIRlJs8lk1LsdN/1ge8Cr/bTbYac6c/XoFVRqqQfWibvYOppzN0geyvb3TjI5ZiqQIo2hyiWHbdZ
LAtFSrLotXcpII81zmY4mHFzsVK1d9xm25V/V4IPK8t35VAfZoRN5sB+3jVrssrGtuhdNlRBTCEK
KuLXA76HZ+r9At2DNcrOt8Qa/ZsFLgE30GnKzqzaJ+bJmmsRUhVTF5gxR4P1AjmyP+M7uVI0mts/
J6PKTMjPJBnf4IN4t1zq+kXvgoZXInjfwLMX6J//rKiJ6IkTIuDK+cpTm/gwQ2PWiMekU0VvDJ/k
/p+DnkG4fOhb0lP07pdJ8H/gbhwqNE3owX7M4IW8/udjplvAt1t5wV+nGLp11VhQMeFJ5fvEcLqY
oPN2T5qfR6bj8hllD1BnYyMmWJmvW0GoL9jhnauwnYV9W9qxm8HYoNiGwfCj/OWl5RdYmbtH2l3O
I7jPjHftINaherSFypHiE0fvGsIfvR4h/gCXmjzKEwY7NUnD1Rb7t/8gxqoxYWlMk5BuU7WuXM2N
Bg7NFioLb1c+nJ3l14yCQxC/ebUNIgVK9TzUKlSnhGn3ebi9mqbHGgqGv/HVzh3V1hF0WAJFle/n
46+CJ+ByBl+8GLBOVApyDgI25Oe1n3Rwt8OdTPHr7dgs0QFIxB3isiIltBGnuuXssEOhZN8sqCOr
71Mc9hMs8GoQkUeXfeY7MP0AekYNmd25ldpQAt7M/zOyd57U51QzWtT+5+ZyCy6A+fTdjk1kdqAV
i+vIZyDfiilgC39LAAvjWdUqTBhiGtGl0FBiZyqMqLvYmsf9uia4XXZvFmw8TZk4DezyPQ6YJKyl
wFyUkSlvN4bd0LlagXddEjd6zML8XvfZ+zkIoApE3h/HQgnmPS5hHaj1ttIthWVvRqmV1B752ivS
GK9n6zHCnSEnatVU5OuLEKdFO9JkmDcmW6usrWh0zurmNRAnL9EGAZ/lD2kbsndyddB/a2CPvi0r
y4PK9dnzg1Q9FjLWOsjEtgj8i+5lmzEufrbt035l//Rh+e6claMqjV0aIXABOXy5F2kCVxphQzn+
TeLNE3J2eftqE9IqK1/ZIdxVjCyC3g5EfbdAoIoplpEEy7YKZkRH4pLTGnWkRwTCWUnDJsHm/tqM
F2L+ujpYX6ZJp164WYUpZbsjLjTq7MzWMbqDlLkYDF0bE17bJVvKfD5u5djiHCV/GKGFQ2zKukh7
q2C2A1E3/Ei45FnHmUf5th0BUq+UeHDdgdMEIuCk+lk7950tgWAPY/GUV0tedGOdZIm5qTcOyj9q
QBqip2OZpehlnKugROAPJZnzIJt0QrPY5KtDjeG+qkoNzIAeQ555O/TWPfKqGyDO4MjruF5vN9sy
jVSrRiOCpKML9LEg8WKJWrLELx1bDkCouesdiVU/xCz8kUZ6zHmHJ3DxQk09W5t4j8GMmmxuccUi
LPW/4EdU/Eq2qMtDwz3TI/wLZaMfwXj0J5g/5+JTsM1uuHLnU/PuccJLaYaqKK5pFuloHbVJH9EL
nAqfj56J6o0eiwC+cYJWLuDt6P9CE36W+XEwUvtu6YbDuzCy0rdo0VTi+x0eYWBiLbJ/CCNGGM7B
tBlTuK63/4p+8Kz8eHGoQOJDrL27RTGsnfNEfgHRFRyEKwVAgk6YJ5rJaNImhFm/F4+3QlZfPjEQ
3Os4vztUXx7Otq01VfF0dwiybRGjl+i+tyRwm3+z228OV/OFQXFcgK1/YAAlJ/ma7i3ztIxZ7IJA
NVHKN3ZANwb/9MI+9DRJQoDbSNbNXFtgpjJj+I9HV3QUzbtUmUsmP+fnEX+jGI18b36PSn+eIx0Y
9ohBSTgDXbczZ7aXxmN4i4G+J9zT3NycHMXtYrswIqudJ5yDgkVIP9b17h063wrpLJ5vsPeLqANm
HcluwiH7b9/66Lq3Cmduv95tLQo6SBy5gg3ClALE2pwh8EeopAzwyzrVAwfsSaVaVBsl4TLxn6FH
cj7994aRk8Vr5V8dQaBuPmx/2aDrWUOWTK13cGt2oGJTZby2R4FQdXmwwE5+KL21AdEae0L1yXvh
89kanGN2mY0fy0tB12TLt/s4DTjoGjNW0SBD2jpk5DX10CPhopErfuThbeKBCY1OmZYiU5EdwMHk
OV9L1iGsbmn2nV21kG+S8Z0PRp+thc256CZag/TbGqpdAiJ45a/TiF1VTaPHg0mUbxY3NL99kP6e
wotrZbplHOWeipw5UwXVGVltd6RVf4VjmPBqJfL9ad+AR5uQzYKozuPAhqGmUQtjtBwLhjUpCwL/
tPp3sCQ90wVvHDY/sVUPACDEWnL0Kdp1C4KgfzZey2obFYxP9MKN6bYzbn8gZt21YMRDSMOeVW+H
kzHwu02GnEOpAmGrMJ++qZy/sYHdW02Dj4fI4MVDTPXHmbKXCYGivofy4PgSIGaO9nVnu8QIoX3a
uzQsC4kteJ5lzXJvkRLEgEUETgpEd6ia+X1KWuDVl+oQMOz37boAyiF6BZNJy1gxHZDMidfgIhJP
MZxfrgee1KGCXrRGvxps2sxuFwTgiWXmo0nmsj5wW1exEgJ8RaCHEDvVTgrurwl69DJtJJ1o15t2
PNouJmbQZx5+krseEwKRnxSuLjLE6gHOZmDMInH0YYnwF7q7op2NWhPebobVd26vyR7PHtseXA27
ykQKpNeH4S0UfR37tTEMl42yNrM8644cJUgCuJmiNGK90ptbiJh2H+JtZYi7CUUbb538Svv9K58f
Pxgp1btvU89zNC8tuZooZrqK+V4z9lPdSqmEUA++1frGnMvY9aHabZi5p0ZE3E1DEHUujIxqCXHn
JMOh9xMISHBxtnLkCsnPf2pTCCj0TdxxXvF8QmD4uxhjo7hL9v2C6IaxDhE0yYcMDB51fG2FYQec
zUBF4uEueZmsVgCb8mef3g950TwworRhyHuIzRDXrK0JAsBtyVl9VfCeRfiwxHU9GjYa9yFEA6td
G+PAvFQnRO8+A98A0Bu8TxMQp4je76GF5Ad7LhwRFFT2IlnGB1EtnElmUjdSjwKHO0ciFio5yTFI
h98l4wtW7obnRklDs1GCvbx4eVWyCJ+dt+hyrJjrUQCaNNHGnh8ETbPA1YS4gedf3r/oc3rYIHlg
dM4tMTqGkM8VN/ssKnxwGgeqxvgNM9z7blQFYyPdW3ThC/+VPWCz+e3SdTYjflwR5F//HzbMhy6i
SEUeIl96w07+KwsHQvhvEbjTS2NsGejo6esRfLXebEQNmXabpaKo5NoFZu30CNKfVwIe4quBV3gL
qGxac9ZzrBCk3WimntChA32IHHk/2Hwb5r55ehmuID+mklwcDR687dUU7a++bg05KKuYsCczGfQg
EopLtKqQn7tOb/pN0tYBEWFoee7cT5YHOlMvSiGRu2oe/u9DTbPJZDvu8XEs+g6ppwhIDzXjJJx6
QiyvqynPS18cGtBjYA/1gHZdZPgRq2DO1b9SrX3N234baQxcHXKPA8cxF2jrPLWGbbAuL0+/x2Bb
KRqeG9mIdZRdEiEvLVxs72rIzQdrIWloMmUrblZ9Uy9G0dmrkuf/76AM9PSn1oCp6ocNh6ODW+01
wCqVot689vKRgysNjXW/rnkrxQRRSVgFWOO4eDFVwZWSTA+6JPx0KKwsQDJc21XHIW9oy2ygHddC
1itMb7khvXS6TnNST06REs+8sIe0UCzrQDfREspXwbyoFZbFUWfUb7E2G5ZO2ua/5Qzr4THsMSNW
KZUvyC11cWs56oN/gIpsJXL8w4HkMGIcsJL8/QM9gWb/oDMUNgGy2EG5cZkzvRHMq1Iu7Mg2SMHs
0DaHOxIt95PztYYRJ+5flnNSZZGVGXowFqibtokhXm/stdM6pAXb3TBG7FkxcK+D4XVQGHUX0put
Ussdq50kQ5Bh4DDGI8w18FkgyXBBMvA5Z7XeabfVrXk4f/O8dslRyoVrodSvg9uXEAGJ4Ok0s/gQ
pvCHgVYtcHvRiwTEAB9ZRTe/MZL2GaxaImPXxuyxqqmyc+bvBvxEkm8+DGS8FjLNmaUK/8a648p8
cpxArK3pX60NSSSYOTN6xOs0hGYMKvwpGnwXbT2EOLiPk6eb2DnzOuf/pHeiCpdT21BR4H7MlyhU
WXHAY/8VvJ0tD0CBrbhzg355CQm0UwMdbjn/12XxhUwTh1W1stSz5IzkUE+IFTqrt5Dx5QMD8Pw9
AL8dmx7yC5JZ5XsgJEzCGFstdmFp1+0IeCQTFGohkzO9ypI4cj3RWl59i/molV5VxN3wmgvwm/Rc
I9r9BqNpTJIZGS7JKDm6O9vfumlcd5aZtDD5LC8NwmzV4aCU509T7Fh7bVBPGOTSRCF86td1T3+j
VPjIWX1ePu9a4PffTjN4jMP2sA0vsGdPS7aiDTyej1g5T608ghmGOmSdnbjr87aoAj//iuV71Vzb
TBkm3QjgDLHktQwSJq7YGeZR5OsSHQyXs3fbUyh4H6sw6u8jD2ZgcYUp7/uNu4jVvdcxcbx0Ob5h
60+cZQI1jkVsSYdUlG2O682z6Twr53N14ftLhea4cqSfgr8JU3KK2OyLqtqctia8PgK/Aj1+bz79
Nz56Qbrq6wHN/bDVEgKHG0IRrYeHh1j0h6dUGbybIRz92hc0DflA2RxfXG14Pc7k4YEe4sv+ECXJ
MTDmSDPAlTrrSX0f0INlzTjBhgIVkiju7iSYSzBk4d7IPaqv0Una7wYSZs2Z8sbDL4K3ilUCOJC8
RWdQ46ifqVW197hfXPvD0ZtMQOremNDWJibxhmV2I7cuICkjCL38caFUoNrEB/eIql/KHF0DZTga
0eJvTg1R/fpR83QKjRdqNtJwhPJiZ2DXLt5o6H5BgRYLcfE+2uLOJ9IPXEHpeuude3CEiYxxvxpM
4Cj7w8hBXx/MQliSYv5AtVxPN/KE3PETDt81QJXyUv6GTYFxv0zBHs0U3y6IEXfkX9BTWD3AMNUl
I8fw4kRfA2ETMJtu+17+lUSza0WQfbPCuQ4lY1WbkLHhYRU/ZFHoj3uQ/YHAiTJkU7eYLImu4H0E
n/vp5Ak1DrPlGgXYtWO0uQTeMjcOfEC5T5WjC7neynkw2IXGXDGMQmO08PHwj5xRPzmNLeZ2Wpm5
3BHIcj26pRbB0MixUFSsPSDvUiPT97qbWFAEbnAdROEscki45GngkYYmPUtxw1qaNMGNG98sGGO1
BnQ1mexIOa1AY9Sj7WY1WYrmEcpr5M3ZT6ldgGnYGwUGeYdKvzvdPa00INjJ770x19L80uZM4Alz
6cvqrkDDM+n7xNKnwWySg3b/+l9KSwd9UnJ6Paq/Za8mQCS0hYwXUbgpRrqHFNjA5bRVZc+HC6xU
6VKIKXPHEmXPqH6x1qrSXOtDnCKowLDSeZ2iSXPuYkwMmMadBsscAN2xQUQfklmTMVIycwodoj3m
4TXyqElyB+y3CtSrUrkDjkyHz/zTgWBCB5Q7PguKQrFDbX8xtFOSO5loFqBPmbmMdckYrh+irHF+
RPr3gwq2gaFw50eAmK1EJ+9h7xYqhMdcUu45DZH9JcryoRDWOzr0ILWUva4r4+xIHIHfa12Jp/Nq
5C6wz0e4aDSjQELfBBG7fvblXI+tXVlsKEtOH1O7n36VhfSP8EzSoeigwFtFPsWnZK1NpQGICrGD
SdI9yUgDRGEDdQ2CoYM42Z/kq72rMGnQJAu/JdEfb8v8nGjUg8bLE/c0gym4kK53AS673yND8fSH
sMNykQ23s51ME77QGU0JZ1pQENMazX2Bz305jlQX0iNUnslZVt9rFnCeVPW7aC74PPPqLX1Sj5yr
klX1oUVJDnFQUqweY5S/aY3RuAYF4r+mqFoDQtmwP7xXcuAfcAfhCEe2XwN72cpeLU+iG+NXYCZf
yJ+i2/L4rDTa+VMiR+gWtott+/Q5jQ6Sy6WcF0seEilREAuh1fIhphXYQPprJYrf9gqka9oWBUQ9
a+QoeMw1YSCuFY3Qrtqj/J/SjCqLcBxs2PQDBGg/Qg2cYNgUtDHROFpPjUNKqX664eTrg9rgfgdN
e+cFn9ZVexnVjm2Y7wZeRb5ZARAYho+G7cho67PViZSZSYlCl0CzN6VHC5oX9NrnSPtWxmMMUsC8
AGbgvCQS9TPGUy2FXwHyP/CTweZraRdJT8O95o5WSaEA5DvHzO9ceOg1aPWkOKlSdK/QV4n5EZG3
sld8KcjE3YjTbSXsMUKZrY6mBn69fk/E1HLJp+90XxvuNCEpt7rHIdHKGmhEO/6Xyiol/ShftVsa
idmbw4JU5zKb3q6qUYxHnAUGae8Mv+Z8eBBckfWgqYYs7hetmaLqiX8sz/hVGckS2vbqim5L3hOp
rPe8yioo3Ul9qGz5XFXrEhnhNJ3Yno2dw+/Fydcx19Xohp9KtX/2dRzEvxK6DBjMqMvY55t0GyNK
982ESzkAC/lCRIz9dm5uoMfpyo0xxE9vhKw1XszxwefpVDbc40VQtSHua6QMx1V8Xg7gHegP4gEd
rqA0xjIgHommRhHo0s/KAczQkUo7GnlEAl+bl2Wby8mzcvEejJkXhkFqTvbO39BhnkUJy0rC+rfl
qubdmH3KbWD2D2KUl6yXgIAKB7OKcjPhnV/JXIhJzTujA2vPj2SrIOiFZ7JBinqvyOXMTLT7jzM3
9laIRJPFXjj5RmslhKe9CRY24OsxB8W+pb7XFCzshNdjFZ96sZQ5iX9AX1UDA4Qvn8zwA6IuYodL
AfxdHKHpbD7uFjkyvcBiW+jwdcabRWH6trBdLBsZv4rfd/5PHBfA3a9pNu6TbdbfIf9n2Rw1VGlr
0Q8uqU1rQpzMBRDV1SVPMVmb3oyhnEncXXGi+QdAdKAOpWtlzX58SQexJQpkVZLkoZ0jjCXebJRb
w8g8UkKVehfgDzwoesm8qUj9KRrrF0i4fkZ641ml1EdkoO6lTpl5wgpBoPWIRZQhUmB7KIyUFXFP
Mu6j2btnPe5KXB2MCED7ZPbJ3NzHxjELCfngiMmwwvG7MGG19+JlZjZv1GiwOE+AxBzT882Bs7Of
bfKEFY+843EVWsXUEB2ifPQMeAtZFatpEBxLmGcjOT5XxaDTXjqotONt+DAkTnZovGyXK1fTd0Vj
YNP38hj88eGxeSbgrboagFjnpPKgnZnl2gedYk4AirvqQdgb0iwpMNv4zRSafXrpJtIeyfZQ5vym
8k96RANzMu+khkKQrIPYyeHlHk8n0qkyOajrxBa5CvzBY9skCknDn8YykJrU2ixtJxst5YSiPxtH
nmkFsExHxX9DwVeKmBO4lCt3ENkPeo7NgQfYrlCJIp5+FM2iVNFKPwQ41qSSFvAmRGoyxondFa9y
ZXQXFILXGisbMNUHEFJJRNHd1EwbKQDtg5RLPa6chLGe2GtkAuwo7k7aQUd95DM0wMqQobIN9oYV
A5ew0H5dzwSdkp8Ns4SZD2/qjxjIfn1DE9R1yZPjLhN2qbBRKiQ+1vxTjmMB/WAXMaHBPFGO4ZIS
it2WJOR42frdUjfZcjOFA++frTUZnQYKzRTaZLu6Q8SqVwqpWm665NlVtYX32ADyifWSM2+v0yG4
w0/pcWihNZ2Yk66JOs3Fq86a//6+ajMCnQtEgj8ILKDCmTljMwQGmqpVMSGAVB/YeoNMZQwthAyk
pC1lVdBlDbEfkHsk6OpYzopMvDL+GB71/Os2ct9ZG/OeXdXlhAa2zOKi4Erofo6eoFsp4QlVikXk
vmVERxKwOLD/79DXpWr8XhLQcz6iR6aYn/2e0yNzZNpeb0/axtJvlXWPI3NLYSi4gaifKYz4G5BV
bmw81HtzI1vphFI5+k6GMmFgincs3c+uHcJ32ifBigtQSxUvVSnWHcEPmuDTW/ddyjuwx3T9NdFQ
v2kZbgfEb5q4ok19QXPv/ov/ggJ3TpmGw3bapMxyjf5z6BNZHs+9rpBos2vTFTucG427+Dbgo3aF
TSRZhPcncikvHiqyS01HTbkn92O4m76OPor9MPnU12dzLzouDkeU7RciMPRRrcRfjNbyMmXaHAcd
4EIEfdBKbLB7LssWiJzUzFYtFgehVQrclrjFuWVTSzA3XPsQWgXJ1smAifSZdsIl65LDktCrKFcT
0S8Vc918TNMJeNIqe7P2B0BAgF68NIH1HFEHxGjYfoLVSOsFEp+vlElTRTdY4HBnvY58C5AjOqwN
42Pxg+wu05hgorUy0nPjgnoEbqioCh8BGX1OR2cKmPd+3RIsP+rVhIYop2WAZ9JcdYI4JPJQYnKw
GKZQMvegO6MZz5zQ7TFEG6XdAIyPTreSqwtptjTe2Y01fRKFIqSJzUrRk5F2UvNXb13krU3X7/P2
XDytgFW/ukddKjEBKznZXgXDDZQK8NRb0PFDUHvyYln9pAfY+F2TpuM0FQUq6SMu81Bab/ax9C0J
whiJvYm1pbKzgzcFND4PsY6Ap/hLY+aRoMr6HFc2khJq0HMyhcNJVARLepmdKTTe+kW99mpfLN+L
eOoGgscDLY+9bb9jat8wny9MTNOWrbK+my4HV36U4GmB4Y8YqfWA/7BzKcgdXUHmci8F/tvs2iRo
qN35ovzpTHuVK7+3lGv0SXs5IdZHQCYBmxeC8Liu2OIOvxwG0Xqxu3eSwHeeoxFG3zPKXW6XEvT4
y6HkxKS7j93M4bnwjbrTWaptD5pJaoir0DNeuFdHAbR1uRsQNqpIiArfArIWLytv8fWQlwEuwHbh
YyqOVRAYAmDfRKGlDISnVWHVpzFC+ZEOgqXyCud3vxxNuKxIdmedLGq3LohCKyW9qvA4AZQ2r5GB
H2EsDvUJnXcqfYd90g/J2vdsKzFE/6ZM84bRGZORRWTzAUZGQ/ONjG4HZI2wNZy2a/CtrWkxU33A
QLypUHhMBrqHOrZK4qp4mCE3Fv2V3ge53hSlf4c+f50wsQHjE1LFdYcD37wkeey4Cyn9uLCKIrVG
+ZUC54YngeSbVwjDe1nTnJWcbfWq0+PsZLWOwl/aeMfs++ybbYFwCemhOYWI9UyHD/j6YNW+SF3Y
BGvfUpnSg5B/FUXFMbNzCk619vghu01E0bDna91XbBCse2HtPWLIf1LWlWuEXyxySsWLk0RfvIDW
tk6vhhc0MvdeZSsS0l3O+zs+4YdwCGAIdAk3u12W6O+BnhqzgejfMOKd0BYpe9hnL/eFzwzhH2tY
cgN1seSiOLl2wPTN6lsrMEKD+U4MVNplVd3PFIhJ7gnPiUHhT1RpQrnfng9ZNa0JsCBbidHyZ7Hq
iWlYy7xp/Mq6/pe08g6r6GeZklWg6iTHBA6XdlaBeDTXWHp+zuLijPFJTZhetpkp0VqT9FHYIyXt
CPKlqDY6SANFBXhIRRsJj2l7CesfeZHg4iK8DeCkVOY20XDUuYXJjjmNlQEGvrDwM/4rUR236kzh
N4eo0VVQ0DDD2lR5Yq0d/hQOk70P4tzENf6Nvl6xEh5Bi7nip0V9Vjvv1c3suMpGTeHRGbsENk06
MPjcvrtBDR6Jzrir1+oZ348pmh0DaMCOSGm+BnKYUo+mdPbQ2BPNU1F7zDOSp+wUqIrtd+iejk5I
wvqbeNTCgvFwgyPtR8sB7lY0zbAlGWmpu5xsDAnFnJFC4+XBaY5VNTqxca56HyFpg1QSwqwefX+f
mdGXLxA+Of+aYwFK9ioAOjeIgnE9bJbUgcfBvXCltb1kjxsc4UneDnugYfpjSf5HqpWP0C3qyi2D
cJ/l1A7RKl7ExCSnf4TSM2HAmtbjxA4YWHFXQ6YySiBExkRgGeogXHAYqHl/tyItH0c7re9Tv6/c
0F1BrCtg60jmX3NE3YKk3uP6aWaKwBOFdoq97u5W2txPuyKIJLiOopkgD2QX18z3LmS9UkmVz8J/
GV1IuveWxO+NgHBoFzhFGU+n6NDbm7HwslrKwla5oq5xNpI0Aco0P9310co0K0WgBxlwOu7duhJr
GyMxtIJd3DM0i6ivGqnDDyaj4ORRI0WbPelIT36zbgOeQM+u4NLoSOh7HHqkEGnHjHqnoFcYrWHc
shERtAsih462zWBBItRJqm+NTTUemBG/Ina6RQhA0SaEs6uTseTD2d0AzF4KxLIwznScodJ4uHsa
QIeuKOreK6ZKBQYP8+30lxmffgyz1mw7DJqFlrN+DUy3i+Pss8k8lx8cckgVY2e7XCI7QY0nfC8Y
2fVYDPtQuE8KQu/QssgSMih7hsLCxeriPcQevhEcMPy6fX98nRaZtksJtV2HpVqkElPqiRrKK9j4
I05kQtUEwM5fGLIshNwxQd4TIb3DjVBGWg6HlsVmCudpWW8+enIA6maylNrTPzgwrP6wZGsheJsM
hfcYlN7JueUyPeAANLgpaufWuNXVw7Au1fL7mbU1npYG+Ab7DVbuGsivTmJlD4UKPYDNdBK4uESj
t6z12STq65aZBK+sxpdzm5kKilhN7wTZ3MWV8bykNCVXFt+5lwyaVCcpflW3g5kk1jeRARk00az6
lj3/7uuLIeOxn9dPNG7Lsd/6THOVvs2uZGX/QqHhMwX2WNcr4yy9n1JR5vOxP+Hty8fCODVzidgn
NiaVOQlKTmVdLcUgnxBCN7dRW3o+yxHXuMjVtLMSljk3MKLSS1wJPJg9GA2LRNHFyc7KhN7HBnrZ
B6F4NIg0TD7VWkUDEfHvKrjLZ8/We270+fCTBMkojWy08EHbFFjVxVprLoDqetGnLog3n7S8uFXI
vLbkW5TJ7v88ao1IFDGbVz1Q9RSFfnGC9n1XSm02tGVpelGlu8Ddutz4Nj+yRhAGTqGPNWaNjCC6
quWDAvesI6Y8jsAHRcHIyR7DKnx+j/MAo6Mt8ahtBIBGbRVSFtZAm67sJGhWl+A7177mC6WrIRK3
a5VCAem3XuSlBouMCFl6lzdbyj+L7mCE+xygfuyNAFwoDL4vuEjIyk0bFpgikpSmSeQziPaK3YH4
PNsIupPcrqdhfP/KZKIHr21D7sRUQsLHon6hNPPalc2FRReyovgEptRuWEkNrenn6lryp0addHfu
ZVIaXR5t4b4lcv9OgN7imN8/Rs6xxXJZzadaIEu/DetORB8r9TSpZfcmcb+dQXR/BruaY43m2F+M
vZ+JtVNQpOFEaGXwaGQeuwKHrt13UOMxYbZlkRrC0Rdpb3J9msrlZMgYOxzCBpg5a4JMNtKFU7qP
4dVq0yIPitPuz0qi+s+O2JDHyUL4voBSyu3LLlglAtH8qDeSTQRvsxwmgcctV3t0g0btaa1hzxYe
wQDr7SexUMP7CU55RhSuihGf/vRmOP6Qtd+EMMiv+fUX6Q4K4OdM+k2V7dmTcyG5SKMlZx2Tk7e+
ZiqmqlgemSoJIb+OaI8G5WTPGU2l6bErEVURD4kdgRq5sZPooYlMB76yjXajJQ+oMhWPIzsGnypV
RPYLf/mo3HDA8oLLAl6I2Z6dosuBTZEEWY67XkN4WNJYI5FssIPNnv3Epe0sMmiT3mDxyyK8Uq8l
DzX6jpWI/CKd1+IbSUNXG1rlTIh/xv9bHeUQLFNwKaVMo1OXZ9bacOZb9clk9SUrRhL1JG1+gx13
KSf813liql1yfV1eh5iaoKiSQTNzvy+yOfIiNLEpHR9zwTpYTTB+zA/u1/TyUiMq7PtPqu8tHvcP
bGv+dymHpYMXSIaBOBXhBlvmbM/IhS7DRGMqywyk59fKFtLPWmxGYe4Sbkh+jsMKeG3G0tqShrLh
DOeVqQ4XeMcxqYGIHyscpysi0Bt9ijPx9wHbzbnF2fCX3Mkx+8d/4X1pXiwoirLPaM/kuHPv/Rjq
xQWmz72LxIWpHtGkjyrYS7OgfoB3WTj10bCDId4VkuaohIgy6w9CZPejTiTYAfTJEX33vBHSzNXg
9MlavDYMt37STKBKv79BkRfmDQqgJ9mYpAWnft8rlBClnat0tFX0CgCWhX9sSvxseam5Z6MMLMkD
VanGgqDyxTSwNOm+6UjqWlUA6IVx0kYxLQwS+fC/LV/GfDvTXFXE7fMT9Fqh69MoocXuS8dRy5Mw
8zYwOVwUGVZq2GQhTVR93//jW2HxNGqYJF7OP38V1sou5zsf+n94CRB8ke/9krzl641QMH3mSRzY
dm5gWsA0ix2L3ynMoOinNTTIGvqFmXzvsY6XxdDv0N8Au9jB1FXAW7oMkgLXFNP/G49+64hL/uLC
JihVnko200XL2rM1vZencQGsrDEbaTK2y32aKoRuv1rme2ow+wykFhPHFssdn7pI8nfE9AMVP6Wx
s9qDJsfYhiPTppdnqSud4ET52k24a6mczdpjnxjXBEAISM4+IQ7MGEbJJN3Ulya75YIWgN1RP+C0
z+k7OEuVOK/WTuOpeWZFpobI9TjLd4WPp8Apw173LNbJYlo1qu0Z++hCvbgz7JyUN0UDd616Qa1s
c7AMM0dnvNjw2qSkO88/g5kgUhaFpq3JKgVGgCeUlJ14lTp/DbPZOjTMuzZM18uto5tN6v+0gZVE
zIXxYDszx8fVdduuXaFV2YxEGovGpPLAp7TpUEtYRYVPAtzTiW6JJpkd9BAR1BkKzZ5BG6i3Tox4
6BrRTb7Tca6wr8dQYy+E2RIYHKXoFBjHIpeHJnYwKtj/Cmy+w971DcpCuVGHB0clJiMPAGN57YaS
OWYBu2Cslk2JoinVoCM3Z6M3nrr1qCQ5GZOSZcDMVNC32Y/L66DjH2rl2uzSmSVc4s49yqhZ2zFD
BzOo1bYYma6wxgsWtn7J1isSgqpmhxmpXfGN5t+B81H6RVdpNJNsxxfPI6S3ZTiXJhtaE+2NcRdJ
dOFsLVCPUfUM3FMLTWy82vLQAagRZ7zRjIZgUF7pxPLMRMvJEHkYCnGD9vcFZlzmJ1PP/y0zK8Mc
1Lw0vpTiK+YdXyFDU0M/yW4x+qMFTHZ6HDP35Dd1cpOOu7fy13QEFaWoMhqGTaaaavnAiiF184eG
VZXHM9dz3c1324Un1C0VHKQ3uE9sHWs2DjRa4Q4cBDFEhPioQ2bxzD8nJOPkxWGfS/JtcHC5U40n
axvPFGr6NzkBHkrNK4bFXPjYEEagfhtXbPqqSzqFLxFZ6wLytRQUazVofi6ir3wO6+wPYg/+P0EJ
/FEIh/gDZ4xnjvMDKN4O4tSmzAGTsPp/HBd7N7zKhQ9k28TftwWZ5utJVmyB2wdJUIC939kAWJM6
+AnHkBqSK8G4Ao/7ZoKyHOTA4PmRurDKDi2T86Xmx/uUQCCsYcO37eY1yCA83cL7O4cogeIdrMUp
QxV3HauTxU8kqTvGAPBZN4JGLO9M0xxJKkJzgM0wee8uRfCCHTVhNEAx4es9m3wsw6PoHZf0iRrj
LWR1tw3qxDs7SvL8zCfhFj8tB5mLgc0q2HTcjajkPMWH8adYreS7JBqG/WngHn+rYWEK/StRyueq
cwzQwy+UwRZe6smTrNuPIgxq9IM3txuMmU0sW61eshekSRXoMnzpDRPy+tbNna7z5gbEJIEPErop
j7cvyHSQDZhkvdUPqnGsSs3R79RgY3sv/n20Q8BdLscHkc3RnmVDDm7XBNqlWCWSClCkt57vbjoT
Bc+gt4ayYoJohdVKCdqfJlzomEY1HkBATi1HseXL1WmbZIaVN9s7pS7bJSNbDYRmDsyh0yxT1XTM
zIrxGRtKdesdwpw1QT3TVBsOXhwNUDBjbEWUcmesFyUI+T69ziN9IKspM6a4CdUGZ34X/niSSmPg
xYGU6W+R9klAHx4hZCMj2a4paVoz6PUJf+lhE/qplHaSNFHRDGdjRxmFRwJeDX2M3yymDt8OjsVc
0YdwDB+Kra5WROcyKA4ruZe1tBE1kBxIa+pA6U6Chen4sX3XCvjL+fxR+GWoEhSlNKHizOXE/oR/
BL3dr4OXOHOnQYJv+SRo1oczbaH5ffeJpqEfIJ7gFLCLkibed/V4LrWwWPrSpOyRorTFLAenDn/Y
ewQVdkyIIlbwZ/IQvwp4DTLkLjPrsqkoCCRr0HdM+AgUvmFrDHWtOP1LTBtMT9nyjjQlwXsha1XB
g3/IQsFPOK3GfRbuvbz1Gw65E6s385IFWI5K+Wki2bJlTCpbrJTPLibdgMm3wGc+0Dn1OITpOfhr
XDpBaP9CAkhMeXFnd9la397OU1aRkFJlt9XxsBZEZN0lICv2i/K6iTS/PLDA89i7Y4Q09m2HyObF
vj/YSywGDPg3oJ16biv4XNh9kmo77/3Gf5a97hpMvhTKwncK+WgLoJZHs3l/XKfT4uDfiIXkxHi6
ikq7GNw5kIHIfhkebEX3uQnUVx7IgN1LmQT0dsTqZuEcfHtqElIVTXCmPgR/bUz19gkh8LbiK4u/
5bY+6oNotPcNnACJU9RwEeObL095NtKRNu1ujNs4xU6gPU6isqBi8WpLyNdpL+V2LUHCGsmSdhSh
LVHsBNnsALTlEfZZSKBQnOwih1B6GlPXgtaBtbd78pWq5d4EV2xbLnzOQ9gZwqCD6a8XPXdJ3NoQ
9cBqJwZDqbdqpMGo/BLIcFWVY17BqbPlrJYAPFdmVeBIA6KvM+vG/uf6gBYbisGL+wh2b3bXkC08
wI75Bt+jswcgYR1XjlfgG5cxLK8vbkET+qgHBE+91jfvOaWpuSYcfIRCDICCSI7pfyisfDcNy0Rx
Owgl7EwGMapJreEwAlW4ansto7EbFipDR2DyaE/FE094A1oBX3KX6REKqsrbD7gFj+6GBAGVJ4dI
jcupVed47JC6feEplPPzT7HsY6umzSdQT47j5Cg0aDOSiMOlb1PoowQa/AugN24MqzDuOmTr3Sbb
R0vS0M4hG++ktzp9jdrEfB91n/vU+sA5kz17HtY9QXfkwvYWWEH14OZ5A1U+pT8D9X5TsizJCE29
Zr0yXvCfF8z2ToHFI3SZ5fUGb86gY96F4pGu2SUgUiaEuFIBjTUfrITonUXBMaeMzDkSN6BAcRRD
kg/fGr3j3ucNq7SGWBc+rgsLwf6XLGEsk32hd9FVVglgkPuZu1JCrCqP9rbb2c5lHuu8jxjj+zx0
++520pfcrnckYVcKqNECjiMgAdPN+A/JwZX9wgJqN5Omig0QfFvr6jqODkC0OU6RyFfhxxcd5Fja
s46dneUtv4RYHtEhx0VjOICqzqAUncVQS9H2B8oy3d5xYeaiiFgTR0zUc0tRoKP2sDIZVHCcjbou
g0uPABOYLH5sNt4+vIqXGAVYd0vH/u2cQR1/cxySzLDY3/sKc3MFqVlLZ8Id8uyOZLTOeDUrSKvz
9FFohTydzoY1xjUQ/I0GdW5hbSNifInyutkFRvS1PEptprBv6vfT1FC6RdTxIFCsV7j03xdkAIG4
nx4ESx0gOGkGjVPSg6kBeLGca3QToFlthY6zWjBfOk5sLioIoKDAaJ3SSFP1OcZPoySzJUmNAkic
Wt0tgtdsG/5/2u/JtuaN+uxbn7vQQRE/qWhgk5405xm+AXUQB2AUhij1yTdRFEXkeDsRCychUn0F
96G8JHpkhIx0TykA0tp6787d1xrCJEbJSyY/Qc3Vyaf4wgDt40NtjljOaBBM7pMXMNTQ3BkQYV77
6HLYEf8SteBqO/JeKO7h5yykFWE46MkqsZ/221WWIOIwPTmZcOMCKQb2wF7GIiRDQlghakcW1gzD
2Ftd8wPG4kXGm9OtZ+QZZ3458/GtkLZ4Bldc09hv7bSKtuX+rrIyoZMtoillv3oFDsb70ebO4hUz
+cyhkv1TzNRXSjx+smz+OCeA/XTZUR/56+RWlqxb6KRYtQv380i1Fb9Hk5zuq9Hx4J/FhRin4ac3
VjNuytJ5R91/wzjoPi1DM6r/HOljdlhsbxc4Me0Pk4vh/rDLkAEijU/XyewEiIXhy31Y1NOKI2q4
AYF6qmpFj/vitej6V3ZfmomzRyKjnD/BC8ILGQ+9TVSHnfjhaZ+GRcoawl2vPcRi8D0DrA4vXHDQ
CbNKGZgTjSkQZLfO3QltbtNnwf0pyhTrGEJEMgOFTDGES93qes/K6gK/sIxOL2HDHM9pn03X269a
bcuJsFU4chkgXBwLsBp3jaYtgdTxW+CcTUvY+JSlnSdVTb+Z04PdvaQPTPidv7wIfPrLHtRl0JsT
/0S6sPKOKS74Ta7nNAQnSBzal14SrbvXFbTr84tRNuygZIjCBUz4noEndB8MO3Cw+DagmDd3/kHQ
FH2ghuDQo3RtFmj2B9fPWRiD5w67AV95dKh46o4Y2T9+EObrgTQB5c2TlotiCyYCWX2o9ueBmD4R
9LdV/HEGBUt1iivS6VETrn82rLAcvYb4cF0la8USATsqAkk1f4HwAomcXL3tPKkyEq5S7JqDin2Y
v55mbAfJ95fnVzz/yZfGV8pKUVCMQV7XJ4YXlVwNdGkFj02l25fidIihhdEqT3wAg+Zx5fp1A01l
NgOyrFcQl0GhDHEVH25vehqdXnCZaSt52jE3TZnffFvjDTYtiR1KYJd7I2QpYHG6aEQh1Phoik21
fboNTH4wO5ZCemKtE18NNaYZXNZsnlFhJCmPkOTOasG4AWPCX6Q8kYw4tuwT2nx/+9tczQDDmOl5
ebImQ0Z+ItXcvXUdiwUQQQX6jQP+pmpEB5iGEJYYmjXaBTCviz8veR8HCm+6z0FgZ39ajTubHQq+
oFFzwcoJOadYH1UxxNHZjuJx22GTE7MJqBbbgi5yIdIqjploQkl9fpeVjk2l4KK6Ph25Qnp/D036
e+UkjfokEvcNierOGhHVnuvmPsIDiRNfjU8glBdB/XGoIDzfjbtG8phawlPBA9rqzo3Rsbbfx6de
C0f/cv2gscneN4q2evxhL3kYSmYgpMXnT2LkOd0jHMVgd5TK3Q2gtherjY2ulgbCr7iQHvdclN+o
pF7YQsTkE/tEwBUvpdDuP1Por1Ad9vQSIivD/TOPN38LNygFTv9ukAi1SAegyLE6PpkxFO70HUc8
mXB4B8qntHc7IVTHGmjMTJ01/r18gcAvySA/Vh/zlLgphrrYHUHVxXSuwEnKIrN8VlIL+PU9J9Re
WUOCEBOBtz+hfrOE77UJSosbHlSzirAivEBMOf+X8n+6eFK8QABB8/Dc5+jm8BSV7OQMj+PnQh1+
6hIZG5ir0eyjX/dmV/F0U9YdBNG4mO27xyvbonoKvHtx3XIVtr9GOa3Nm79XEXiPj8WYvpguUCaK
Wxk2Geghv3kenSBGOGMv4sKc7O4LzhAIKa3WqHihZoBlqCLpcenzRsMSg++HVFOxvQixAaWdktUd
fZVJ38p9sQVHtJSEnvPK837qNPcnTB73rpycbfxeyfP1nb87C4nr5RW17u/SIDDTY+9/I0dHatCy
PfeBWYvJlOgcfMPLH3EOY8yEVvK2N66NX7hTN4iK1zlnMHL1JO7K48IwAN40BpvTHT+V48QYMJG2
dbIqSeLt1oDxdcg7C8Z8zRlzWMAdZn3YJgoVbMiIxdfz8QJ5znr1SQOVKv5VvX+E/NfkpitmmIAW
YxohlQdkczGtRD8uutUx42o2kdfqqfUPOxKXA45ksRPd77pO3D155uvColc0a6xUZNWn/tHDwSCL
TXP5klMByOCPVrN2RNPnh6RphWf38s0W62bw9djkL3ECn20EUAJKx2stT9nTmUtDLqJnJ0LPRIQP
UJY0FL0dE5tX6Crl0z97zKzVnC1/Sh0ZsmExSMWQ+JUCkLmHWzUEO+slpPlQ8OqHI9w22ZBXTIJV
oXrze5+NtlOhhqOwS7EkdZa6h956hOlgloKIJvj3SDtB1v+un9imXzGBzcrdMycLQelogpOWfRcI
9Rbo6UsCGhT1kR1+KR2sm0YEA0JKefBSlkO+h3kn7Am04ZXWzyGe0yTmIDefJPnl1GWeouA26yEm
rQImDuj62KeJGTUQRXJ9z9BaKbphMD0gwVFl0o8BV4HV87TQIh4a3vdPjqi+wPfF4SYSld7hIzfr
5/GeyyXb8T3brBGF8aiVfAbSDadKuAiJ00Hmg0E7JcJKuD9zOY9O3m2PRsufd1rmg3hn2D7VxTXK
FDANvsHVyc1cdzEfTzdWIBMOLZKKOluwHoc1pmaQwz08htqp0Xnme8/1jYJyYJTl5auVCO11oci2
wsp1H1V62pZd8TTCgCecY2aAzK1FQHqI9Eqi2lP7s6wc8lmBJXakdBbmoGPWzFxXXu/UijVXotLv
7aV4BZMFgnn2UDAoIgSmd35rJ3EPwCEj5sgbeqJeFmg//Ln8HD1CjtQpq5XdXN1MnMgSuVZniF5Y
vYqM2PQun1wJOt/HsGgVuaPLRgjv8txsiQe2sLBTdY5vyvHoBBGZ5U9SFmDKvMQ0NwnT5cYChy8M
hyF1PEVj5cIrzgAggr9TL6j9HW674UMp/7BGs0hAm+NWAj5k+qblyNOoEQScBHmkP+4MFguI56kZ
55s3nHDR5oCdZaVNg9ViGmmHp7vOgvsm9sZEj7MofHfM9/WV0bF2VfyOIxZXsA7QnZuRJtPy5bk1
41obWNMPxoWuG/CPsZBtE3SctxIB1Gn6PXYzBeob/MbWbnfhTdyJcfHHR+G4fgRB7UhDKkUiie+s
vwo7OH5C303U/r0LY6UjjObWTkPDTsuaq3NtzrGXPaxET7vZ/09d0oC5ElzTLvWWWNgPX55k4r1d
ACiW7Dzoth5l+39fAeXC5umXeIAgPwvprMKe7e4bUZsAvKMqJ2BxJBvlyKxRwmPZ/uXdQmSWAA3d
GiLO3/8v9rijLp1WtGXOWgo+5PkFgW4RALYxDF1WEmA4GiYYtWsOnc1Bo9FTRX2eb58QLBKn8RNz
vG83/Athd2i8AXma2FFtPm19AqNnbIVtla+NlkIkPfaMtzoOUPWDF2qGICrs4wwgVz6fmykm8zT3
Vt2sxSHyGG5nEDmMIPSbaLxDIkI0KbSn15FSnBmO4kmsJQ6umnuZTg+5o5Vw6N3K6bt5HF04oVy8
XA1wCF2XuYkOvf7DII4+nMnAP6jObMSL+iC4k2vU293rJjBX7p2yCmtmeIzWkS/9zYyMWWWMsRGN
0YSLhaDy8w9UXImuKMlhxyzABcR2W9euPsdW0C9R/gsIn0be+qgayGqyVa+c3PRF2b8n2FBwiGxq
7wt23xu/75jLLN2Q40Q9J3HcjwH51tGah3YX4SGbKIHmkrxbEdb9AqiomlaychwS3Niw5zkOzDC5
/PZql0Cd+wL+7Y/CF2CGVytTuksggyHtexGkrRgXWH9AWs1lgM7dTSt7qNg32+0wlmApasTs73FW
noYTL+xWmgMP8E4x5BZ6dTf53m9lhwI7ttqKG4Vdv16WB5imF+9eAhfVHqvOXuq1tbdLuz8c+b27
SVnydkiOebsiXH0EleGqMElmPJ0bAAycJhSYRfYIDLw66F6RXcyUPxxueb5VH2aWME+j4PFnyTEZ
K/kAoWzZ90UUNCW+MXNc0WSl+J0yFt40DDfZ0+JujowbfoPJcmuoXf/0OTD9obpinZpPTKmw6rve
OLwK74c+484aHFJEWojcdgHkJZtSZ2MDV7wN8Z+cTtHHAKl68lRovSq7riaWF5gl7BocQI+Rpkec
geAcgYv0W53n3lQQIV3jfVdMicQaRvrKW0VzRobhHRn9PW9NkVXdM7ncy6uSpyWnHsNJni92fdeW
ougrNa7z4q1QnVb3nrX/BXlwDDJ4e9Qoxc4GNSeTw/3oM6x35k+m5fZMlNoy5FNwTy4EVw/91gkT
FCEWWiR2Fxv4vsHuOyFcdl8SjhOI1wBTHhCzCD5lJpKjH6sFaKUfSul9AWKGr8oVe/ecAAO7jiFk
As+2QdJtWc+aPEekp6ob+tSZqm11VaNJe68oHV0Agi1IzomqGozkzT5CD40b1fQCYDQoy9dHdSbW
2fmC6q6W/l/gMunJgdQyn6Eoi/y5D8cQPeHEu2d+t6sT9UKMm3gVqA9zm6Bjtsk+8/4cY2aFs3Wv
wjk1+cR9QxKtCVuJbjlNbkVCCe/awdDXDFcEBQo8pg+5DnsDfN4VJoxgSg6cUIzNFqz0sUsFXvW9
JhB9Pe2sK2h+zs1g4VBFV3t5GdAfuOfkmEjRR/Wv4eHtBeIObVYjp+BaPlhQeKRgaIZnK8CdrMob
CdXdbd8vScmzrMI1HFP1LW1+VbDbrqjUE6VrhLMEd0XOCTs9YtfHU/Jdy0+jokbTk4U72ZTAk5i7
t2UrAh3Y2N69F0TK/usIzXRuIwPCL9qd9rzuwgiPrV4ioPaGili1AsrcNiX7FY32IetmBcl4Sb58
NW4NobUBp2MEpoLC8aDVvOofJgg+3qLJuz2iYy5fe3+fG/J0zjJNV0pYlQ+14VvunwvEcz8n6T8D
6fBkyahK13mI4Ipv7hhXc4Ade67qYTmnSV6F50hSurhTQuTrTIeMh5ef6nBSEVRv/UYxcgNBHr9Q
nywRBZnF3xAZwpKT5OE8QKw0tQpPHtOJD0HMy7H5kV6Xzl4QHUKq52jUY1G7SIjI2ulrta6ayaDo
Dt7WSeVrrv/fJikJSvpEoVWbe7v2YONHs71EczKbYAom7sJW7P23PUfNjTHFM4cqdjh8dTU9gA99
sKd3TCzC8QNvh0FSik7ujhobhCaaOPTcwCuZSMPaUdTVQgAU/SWu/kX9mYc5qZzb2sq4DPzgyOLD
7ID0rDFQx2BC55K9LmYUd+wIX5O5D3PfCEvxnQKL7kUCkNYJPQnZsuQLy1NJDZZy9Qo+ocnUha56
PU7os/x7Us51vskpBNBJf+WARTefHDHi9gyX9hlwahd8iL3xsEc9gRbqGFtPl4PsTdbsMU0zUwz1
y4zM/B4ucFVzEOoJehjvmXo77DsVXfah4CDKmucNw2xfUtbujaLv4nYkr4x7xfNV+YIEJTlunMnC
h+E6k2D4JdpQfDIryXoj6Fd09dLAjJkjJmwmlWCIHVW9j7y2dBoZWQqUsAHdPAJUyJFj3CGt6ugZ
kqSkjVOGgaK5Y6tu4gt8ByXru4PVZJMa667NCHed+BQKsoIisHkJfNd8i+Fw6BErKRK+3NNjPROP
cByBo76b5Jocu8VnycypQxMEnfh2a0/mF49swi5JXG+gfY+Bm4oVLTDB9Js439stvgL/DgvpuLEW
m97xGEmSA7zXpSRKF5QvEJcsye21alE5FlV5XXd+gQ/sE/4LGMK6ZcHEsqpWXyfECq3n9x1vJVtS
RMcPzY4XqjKEAr4ETsLVyQMKBjUoHJ8t4risyLiIhirTqE9lg6sll4ALHHPzSeAiZLN3eyQlf4DB
d0O7gfMBxjB/xIMGJj+HD8ng6zBv7V+DEGiMTa3XAqYgYiYrW/jQ2uBmfFg1x87u4bo7esTrbCid
cww/zWrhgLVIXNrGohPBINDxXW9k0W1s6f8Qh/Qx8KMtDLLcTE9kVgAKJsevymIpu1oYbf4BS6dF
ObA6iUX8Mw6xfMFSmWi1baXTDc0V+ZelBYYIQ/mv35cSAUGyWEZzrNnRzbnH/K00FI54tI5fdht9
ziEwMisbn/s/iTVQ8TxqN+jZdjaGphXU7bVWWveB36wLHyZ4oStSSREUuYJknxZUrKbXn697iHOU
J7FpvpERiEbkxkYwIgkRUnqSSoel5Z0ONxN0jsiDO8P+uX+nR9toe4xHmSxwyxRkDUOXs4u5IVBg
BH2kybqlaGnE/+UyRf+qa99W2XkEJVDUvRNOFVr+KJjc4f1wvnMpZ0vXnYwCkDn2xMZPyuO1a1zY
pSOcDOeIvTzlJp7xhfzNn5hS1pIMffnfRVlhfb5K7D9bppxsZctAGk3IsPymehm7vvod7B05xpB9
PwD/lewZy/Hvo65ynztt3ijaq13h1yBXbz+430d9qSs2xNosFFJugNMEOupRV/4TLDk0TOjYp1qc
YZkxM37jnYOBPbhMGrvZd6fcnRDh6pHslaV8sQxjtVWj6d80yJnCvlGM3+dELd76mttbI7mHmXNm
J4Cv1BulD+rcLd+NYtDpPrt4m5fnecCJonJGPR1XKDWgZxYQeEXYUBNZipwGRYbT1qTsPmZ1oBis
OexFtejro8mXe3A8WJVajkWC02r66KMsQUXkLhy5SEfnKtOJ691wuqKBYsr5LF/esRiVt8iIS8xc
YZxP+k8qomyCkG+3qNymq8MCYYHZ5/X+Nlh41gme07xmVG/T5vmfcFjUW0mIJwtgL1kgVIYQp94g
fKJoleDYQEfIs8OvkkfNJICCNsxyfca2aOhTgge8Gx8k/XXNzdKe9rQN8kHIjw2+8RLnYxeEziYN
AJeODZpjI2DcTUu6qz9HtOqCUD5BXhEUwmTfBwm5JFE6bZi09HcRRgGIdpfK2oMLJLcjQjizxPeZ
7jlhRFPfODQqLLVpP7ydlx86fhfKHvDn+BEql662kyXb3Lit0kY/sS7lLC38S1Noenfq026p7J7R
6XRzeEMMaD97gXiG+/GrRfgiR2TJAzcVpACPCzH/g2XzQy1DNBGxRjea284w+2sPGyLDJ4vwRqVe
hOqKGlEHeX4O1mg0XpVmgSQn2weyn/g7iDNIodHiJ2njTV1eDeZbtiCxnB51opDPEVb+UKg81ab7
DKnRJao6BbZBHS0yuqISy5Rywqbl8XW52AdWAj+dzTHLViiad3SVEVE4NJzt7G6Vbl5gwp73sn72
LyLkO7MI73B7dL00GIA+sVZuqX9SlIazFuqaQgKd1988PZDV2s3B9ZJv7DYm1Un/gUxU8JcGtyC3
FFHkPoO0jFXzZd9sveg3zwvnTo0mH0wDzaSzeAl3JftA/oq3aadQnhu0jv/sIu+o2O+NAoLRySIz
YbDHlMld7AqOq9N3xVh0PwCAZ1NJh9Lm2BH2qpVh5cjBDPrMubXg9QOEpxsEk6sI8aTy2LsHGojH
X/iLdIWEBxNwrEgG/3P+TjENcn0OmOxBP1zaQw4DyJ/x50eqyKRVqGJJOGVlzeItCylZo4yEFYfs
SjD5EAJNElRic8u1NU5KfIstB0ibvsDFmHCE8tPuTgbYWngLs9hQetm3ei2JT+/vxvJo7nkRstJK
RfBtvxWi2lCUJNer4nzDQISQw00qhCWqUSZ0ywh/BKM1uTTfnxNx9pbuEHPJl0qO5V2BxbLhjJgP
Nh/sUdannPdhj/9i5aBRLFn+Wi2JQGbT+9+YFWNyQIZz00yGZvRE4jo8Vv8+NicTMqBmhG6u2xfY
7rOeKVptXMxUNs1O0QhQySiy8WRtHEcVJ4HMWb+YEYiLAslekI2cKNsYRWQbwl/pPsHRwU+IpJGO
0OQRBhUU7TYq2h/+UE72Q6xdxuCTShbhufQQm9S0i+KdMMoHI0h/bl62EE6wY0luro6F+qhSC1Qb
ulPhlG1MGksyTxy/7BI2spyD+EYZmXnq0/jdtLvNOjvYzgKGffVQkKOL4/aaSEUkMSaY2wp8IeHA
XHr3AbbSUHmaWznAa9Db1RQcn/ZwBbc+91Xa/ZqSTsX/bW9vZ62yHoz4/XMictWomnU2c/gGlLDi
Py2eGNIxV7kH0u0cseqteM6K3cKpcmudr1ADWZy3A2dKRtRROuPw2J9JRDZOJ/laCEu5zw3YG03m
Ln0AQzCK+B2ckG4xZeDiDg5ekM1zzvoKMIBZTY8XlwFG4MzlKSg90jZ1YpTFONwJ+vueqbL32n2K
yLhQSuVgeBz7DL4PjGQqgDKa1Gtp1VfwuAInmS7YNLGbCwp7+aKZZxH3Vqf9Mx1wgajSQsqnRsRy
s3r8iE+NeshU7JU+o3rkbvCS+aIPsyBF73tgNfVmd8elhdcFs/mtx7EtzL4rq+mPx5bCHW7tZL/l
xxF1rkJsSnJxbCKfH8IsirhuMOe/RKJPe5OrvlBFFp4aSJ//R3/JOfG2p9lJbzVXGWzW03K0J+fi
VcNFnVnNhafvPXkF+vs3hxHa+WUrzVpIek3FALBJJ6lJnVUUiAVWxEsTTe3/N53g2ES11C/KPaI1
H8AOndPmEJFutJcvG3Om+9YlfiX+4tz7Oc3i58AEePVDJk2QE2XqmpE0KCfZ0sZAMg5+W3vzkMQo
Yjd8hvVoNdpFA5hbH4OZ+8+0uz2Iz2CuRhnW9eHPST/unKoo3Ob0asXCOeVCGm7CFh5NWVmlFAbQ
IguXTGae9yTPLITEG3R1/HQfoTm2KIOhZjBdc6KszMbg9JsO18ajzu98QeRz57o+Hz4qJpvQLQI1
zTvCdpkxntLDiTLQqNY3OfaEro2AN1wDDoKeBtG+tj7qdjPl03kcD26l5VxvQuUVVCsM9LeTHV+c
gYI+Rquh5ejL/A5BQgL4XPwTvdtEqIWCoVVAViCzipc7rr8oKFm5m65zAbK5VXHZgGv6EIgBQoSb
n8WcSmZ5z4ltDN/wqHlKI/YRyhG43+E0wdOzAC+rvRPnO3SAcML9/1pU89XC6MXdpsYKEGKWtmth
FKJoUReZ186P/CUDdxDU6gDDLbfZLY6rZJHxFujuc8LVOUmuvcKzx0UqLl2fWz0zZFbxYGPOYDOB
HUX73p26lR0NjZsKS6YJVVkHHNPfLhC0MweNihJnUdQDmXVjba6es8EcMD3APbhmp+T/Ep23s018
x9fBz7iG2o8jldnEpgO0r2lfhYOzT5frHipy7NAdeIdueS5xalTkMiLxijm5pkOW0LLFCeUVAA3r
n7qfwdJjR/qxBsyDq0+TuTWfazTl64709B46zRWnB7tvllGwMQaXl+hxllg+pZ0+4PpqAWTOWfHs
osoAMVUQxZbXWqEYZsLEhjmEE/I2YCXg/Si3ZJbW1qqmhKwFFCQSsy+uUZxlI/vPFbmAUvLZAcGO
5uSejGP4CDux3fzBWBsJTtqzhnqU2dDhYECcCbaFp6jy2a8o12Gep7iHghwRVl41f5qF9aoMcxMH
rBvHSmMA/mOV9kQpHDNIB9fxYhjO2JxuGHkA6P/bPz0CUxlgSWPvo/p9M76JJDyhj8RH4UaSHxey
PjyVlrL1ph3FW7PFFtb1+7GO2I/fVJwo3K0a2aMz6bFlw98NDcVHLXEa8/oTCfGrW+mNeAa2sqmn
iajyr9L1opmIbXz71AQKbKR4Z16Tl6D0Cxtjxizw7Nbnmz72JNV/Kf7HSajrvhxmE6BeMVyuJGCZ
KZjmlujy9rHle6JxGKBwy8oiEWcP75UCMoqDlDuQS7iE7Sagz6kzHoqsaBo4J8UCgTjDbVF5zyNN
D/gmiDhQPBrUR+i+Vnls/VnHj4Ppe9DW3GNFMUyVGFhlKg4mryeMkwFBzCLpx9rOaQwRd7Zviel4
qw+lf/zIpQ1V82CRzQ7hnd0vSW3U4jbDEtHaK1HHhAUQ2i7PWnknQ9PEw9KdBhdBagqP8Tjb43cD
5WMz8ZxRDaHPPO0tL85oC4trSRAC/hEfql5RQstQr6X47nvyUyVbfT61EymBCTCsBy2pwdgwLyiQ
QhVLeuIegXc82mG2hHyVK3dMMY+0MDdleM+87T46uM5jgZv216qNAf4KQ5B657cabS67qOMv9aVc
FZuYA+rNuGpOphiETTxVkj5F5YOWI6InRZUJqDGSWg0s95xe+N7buu33NZXuKS78ZqR3/b11xSiE
MOBJt70ach3A9Tw6ZwocCIhQlRDPcX5s0sOGwbWv44LY34NlEN1fY1AEhgyrsEQei1OloPiZjAHZ
ZCkTBMooz+21YUC7LV0Tg+AcS/WX/pFU4QB3aQtP9ez6ywZjcfcKP/+uZg2L8GZSdadUv1kjTYdq
CMZMOGnfzRjOOz1ML2kfQCN+ZStgiBSTuOx6kpR3n4xUuLh/qYLsp0G0tHFHuzEIArlwY+yVgt/r
6aUPFoGJ8KT26lrhbJxCH72K3wXXFJi/uA5vhaSd7xetoOIJ+zdoy3oWk2ghx5vnwa9l9GQnzlwT
TuPTC1NeEx0ITqZ7qTjt7Ij3n8Y3hmx66Kr8SD6T45jVKI8QgZDBzF7XijSXwuGNWZn+98KmUSGT
Dn9oxcBokHPTeFaCV1mYOsCjr/nOd6uZRNKf/h1ov5lvSmrQqThMqEm57xZS2nOgkhVyq8pgArld
1rEyoxTQo0uDw7bCbbMegXHJ8Em4rwVaxnHpZjkYDaCQlxsBO8X/3P/z3RMk8aVlcLz4JRpqaSed
+L5+vB/vaz8whiPA3AtF4xcHUM9priziITRylDT8Y1VQGuaBxlCpx/tdcwWDpTx/0Z0H/1brFhaV
K0OgbA3P2w1KYGgTOBD33WA3pu8vjOasERs+CC3Vb4oqtdgpxF5IxhMXjBEgoL3p71hCmVYvMpm5
yBlcdoQvDTB+MWsMjyY+Yq4NRAzRwf8JonTG8r9nEpoGkyozVky1uwtVQ2v3UOVQ5eLmju2QuAhK
DwHVSkoVWWLMFymjnWEIoWNw7Qj2g8POgqj5RS7cySFjxmKbG4CYDCz/5ejFVBG58HhrWbqo1cVI
Pt1kp3jVI9IPIckM32Ha0ak7R9K3+B3S4m8hdvP4UE/YuO7XOCYB/dxrvh0gqwJ/PCmzmMzna8T+
3yigvNi1bPpeAq9MwOzelLDUEFwRvA8UGPJS0TFGy0H/B7NK6uhvlfmfH1znJloTpAojKZRUqeT0
KZsEc+mHoD+rm4X6AJMw4z0wzysPRcLshMGPTQIK6uJ0M/t3KQ8QmJTksdzikmTSZHKxaBZEH1Z6
tDNRzIKBLZ2kqvOQUqCf29a1RCTsS8uWg8C/Ax+FDtK408m4PeiTlhse91SA+pWVAA1qgYYFx7yu
bqV/Eli8WUO27AKAv7sghU/ohq8rDt4WbLOPkPctJOYQz+V17m1qaDgceDdsVbUlVVSUdBmH3Auq
nhcQMGRh1XJZ3jR4XY6JDwNLF8ZgGpdR7KeUSMjcdm3/5K8MA1pzBM0k0StlkhvE/CQ863PtQV7E
21QB5Nyh/FOGjz3O6ISoqWmCkEEHim3Z2naKfShXhbetD+huWuIUD8orbzDJAOlE7vJYPXCCLZkO
Cf6w55pFppT/RpL+xYoBFNU+0CLy3X9Jde0nvebkWaZAnx9k98phk23ugo7PtvO5uGXHGIlWo8C0
t6mpWIfg8Y6nIo7DwWD/24qtudfkowZLR9s9BWFqHJq3W0Es3scSQ3oD6dyezgmttouiG7B2Je8L
yqPaJhqX/dI3EeUpdenVmfyUmqZOCGaGiOPcQ4zxtlUhjXknx3kqKGrsCvOL+jRVDaTG44nlEox7
bNoQ4ffY7yrrMlU8wbPn19otc2kq2Vj3aMc4QHRZa/dq6/saGnBRvgCb5FVgS7qSX5VprooWjBHt
rJtnrelhJiqBla17tA2tvx4UJPhYJpcGR5DV8nqYVXQRYugRpLJJaeIP/1FhbZdWJ/vf9mnX/jUe
VMBI6BnETQZ2WoNWfW5Y4X67j94wTWClSCeKQ0XsescaI4GoqN1MVByqe+/Sq1bNG7z+Eqa5XnMJ
zapjijp40OOkqtU44bohxTKcd5BqON/kXgMAKdxIlpuZ9UQRlBL3qIA13k7ALbQNkgZu9JlHeWT1
sEz5ShzOrlioUijx+RwCMkRJ8cs1Xfqhdx5Y96RqgnQm0EUR1XjVFhakdHQOJ+CGqgmdHIFofxUo
TnWIgXz1CRzkx3Hn6CWsZ82Z54SdHwoXGQ19gVpq+6e9C/F4KtEH8U2jlDTyqgoYE5kYuNCcBqpq
cjMaMfUEvPUpKxx+2A2Pxajx2HSd49NfnDOVv8xwUPW8JGveNU8Hbp6QrUgXqHlVN3m5O4FRz2Ea
lzORn/AxcuXcEs3Yva2UpeVwqGYUeXMjH7i00FadXVEkQoqVRfD//en0XnfvvdvEkhaaawvfGGwn
90VJX8LkT0r+K/ch6cj7Xyd8tzslwMx+U639SOhD5ASsGnIOGGlHxWBIYc+lmo3Nb60EN2Rudioi
mylXRBZuMm8Xmz9B2X/B3JrXwSSabPJ4SVb6xHRdBX93NZ3XBW/4B6RGMWbokI83nObSY5iBFJnb
ty8SHN6VDp+7ixKOC95jExYbDgeMJ4Tp8MCVYKAE0zR2tkB0hdL++QNwqNz1xjEPuw8j0PK/4RkE
uYq4hoPQd7CGfEkGjAHAq7l5q2YH6L42FU341DxCM2yWxHb2FoA+obgGXjvEQIgTTnIJBvNQTxSs
6yXsqCF+x3+E6h2gVQuKWJDbcdKId7GRbxTUdSp2xDK3XjJFpFLad1OczUKzYIPtJdUv8Lw1e7rq
OEn4ouibE6uexF5Xv45j6b+2iMqfs4cmrsC/tijuX9rXSrRxjBrDRPsrzQhP6yY0kAm7baJKeGB6
5PqtjHknw26x7OSHVSE5OofTVZV1oWUTn8fdQ2CVgsbnabbKtY+/GknWLzVvPzbI0EjfUC/MG7v/
eJiPB9aJATjAPwaUMyFIRlJUJOCEp9Pbfj+sYMSdn+gV3PC8su2vOEbe8OrISVq5I90N0R1hrZ4w
eOr8EHCF91NWBIHJ9dmSJ/L7WgAkHj5nG1RRvHtOM1zlDaOcnj9JRmoyQNkGMAt0zxnKVTTxAmbh
5J3QcCXvjwLDrk0JTKQutg5Ft5KiF66NOowhPZAhhABtV+TCPAJabPLcOyUvVt6lutgAxcn1K6l/
NvTs5c94MDhp2UdK/CHDg1PwVdfAGDPnWnjlnboJ/IrNOU4cO+7XKKvGKTkA0g/6N8RyvBPZ0TdC
Gow8KiXa4izQs7yTr2dEUlONG5h5yILx+mDc+zHZXceTjSH2FhxABhAOItrXI2a6PLE96LqELa/T
WVivn8x7lfYE5TzJfgzgkHzrwf0L0FW6XGmbRUcEQsnjrluMv9LiyRfZC79yYPe3uNkqtRM4qWgz
S5X0+C+TbOWiTnDr/zkXwyl9g4VqVjokvxs2iSqEMEzFIltGclb5Pql0+QAMRPuQ15WtJnkV+MEI
Pf+6O4vNT1pqU/aJREy2Cr293A4qXo29iNGpydJQYg40btljzqH40cu6qxShgjlIk8IJkOCwnTIt
odz1RZulT4W/YTamn9vhsbhBmGj7rVcCyzmqGpQJv3YJfozsewAegbImBa7aNK286c3Il6x4hIS1
NR/HCgKHmTBUJwanaxi9GGjGV5Ynt4H98xmmzVaKCavhkNqLlzpxW8c7eiWPHm8M6/UYtFM1zJpz
lvuAS6IdOdRu2BIZyvFGBYl+wFVe1QT6eQD5zX794PR+b97xeAE+eBkafmWCNN1POVXjusIcMabu
ZRvGaXFLHU9rMxErsT2M77EjmfOwkDKl7Zrz/CR5dWdQneLUyrIqI7JsBlOqiKderA+xumFVwJu8
MxHmJ/0lVWnd8nX4xh8Hcl5+rhqrT5GuwzG6sKkRPwQtsqI+d2pKgGigFyXuY8onAaYw1YpCljFd
hfaVjHn8Oo1vYgH/V5Xc3j9Z0Rjx2Yzg0CirW60oi2PQ8jdaKG5LFJPMY8Ne6TC3VGC5SIvk3iSJ
ztSgHg6cyKAeAwQGxXCTImp4JpsnlF0zJmF6qv5YME6fKfgboWmtm7uIgXLEtFBRJrAgBWwV2uLf
ajlaR7wZ8CoQCMwPFBT6YSNfl3thSfre2MBONY95tASJPMDpwKFfV+Hl4opZos6REt90Ss58rcp0
4nfTcuUkFkoprUPw/hmM1eFQK/+9Q1Lnd9z3VJ+AMuloFEpgpS9O6yGUOjSc3vjwVFtIadgfloEz
wfSwfK2sagFCnsbpRRL53gkD4UdGxuqe+CRaLy/Cmap7FWdHm0UydIeoUds9hyD2Ma+gPi7zJcq4
oBmImUNJoDDd+dGBmUxFlkJzvIKalHhfdj0NLVVx487dYckdtprNjSALqGt4wTKej1bb2RniKJys
GdDrWxJ23Ow/kGmebJ9uEob41qUsUjoBPHfzOUY7eXOQPSe0xcFXqC9T0/qAvE11rzWywXVXnAwf
6jTEADvpcngWcstrZ3JmRDMSfWaFEaG2W1cUkLucfZmeOpwTO4ILVReFDaVwLZALnWPQyySJycTa
AGtm0JaKAcXOhIWgqt4iiZ5yzOiVqISrxrklIw5AJwKL7gk8Itfplpylp3nhIejrw3I9D2+Qs7bT
ib+iArNcfEnTA1bWbZ5tjIAWU1AtP+xTucoftc92fCTIfsywE7/BEl3BE1NbHQnE/r6JsSKoBYXk
4QNjq144QY2HS+p+asvF/1a78xAEKJUbg19Sifoxe5783LXWRI+7f0Ndo968i3JdoOv11nkrF6Wt
ODQqpW8MUZep/wYA90aENz29pEzdzcf8QvCFEWdwPv/dARtzEkTvrAALR89UXcPtEm9R4J70nZeW
fxVud8ujFHqNnPu8EanELNGUWGxOUfkI6vpwuawYS/e/Aq7apkFX423zxHNbe3oE3q7d2o8AazNt
2CxBxGA5r3c06LkxaN5GpoXeNkw0P+2Zy9pMGG5S0G5fcb0ukOSSfnWeLdOnZPHvnSMhnEJDOsi6
UNdtMLoKtudgrHMQlzmrlpR4zerFSf5nxgRsKHJzk1D5V3KTIbTuXu2wHTv9DdxBK5nrWLiBG40E
hMN4u+3/9kmOryG/EWOdcZdDeqVV+lrAE1sF+gIv9lbUoMyQCgH8atCMozwTMjvLWbpy0CwYcvKf
cyi1+iHAozJsUMHnNHFTxfWg3uOTyUXFkG8wArcnpUbEGHC2Jp32sESyMBIbEcvpGAwzVsi6JyRK
N61KUtLTYooyzBUdYdRq62YdIj2OmyTUqtVpZei5YE4utVi4Na+40ixZdVqHX+zeMBdeYTwjMOhw
sZ8YfEOS6D29ruAWYmUIMBMswAnfAGLr+FRcUo7o96k8f7Gq1WZJuFA3dzT+o0jE+mIRXbbLVLHg
pQfCkFmCUz4iXlnLwtjFyIUm6qwEUh2bxNw49zQmZnpnCG492CbLwtnEzz9rVEDH6zXBJaK7UfWf
XON7f2/ZUqnz0godQ2adAkKK8mDCpDUmxnpw/bOwzUopZFKy03GVML2W63UnL4iLj0r5xwznhJcu
C3OMqpKQL9ONZ29eibLJtnaC5YB1aP+gxDnrIXU2hVa3W5ToXvtOSFw6jB5FQrjux+iCRL6hZkA/
BimAIA2eqQljIggujDu5Tkr2844hao3/xJqi2N5EvhK/+kdAHiSM62XEniA4mrywvMcSOxDaALMR
KtSkjE9iB2ziYu8pCbDWudTmWxsGHODVVHLLKNLIgmGfJbnkeV1UEYoI2vrlztKX8c576Fbw0cFt
KaN2ZbE8+YnZZoLnLGjyOXf+U6A1TVS4hJmjIc8R8BFs+x0GjqkDf4NnvSCLIwopaCOJhkZ15cZD
FaHbr2y8jmreVr7ERi6W2gew/4HvP7oyNSk2kFHmQSAZm8dCWDWdmm/yhyMlT03dU64l5x5sCqRu
2gO+v0k7j2ILfir3r3Wf4uUs4HcwrIxUwOU5xhtr4AdSTak1WHoRrDQ7CTjQ8bmawspHVRqUTePH
jfQQX3qz870++vJMg7MEyOT0Tk6SNTHny4+JAJAqEruTGoEpyODXGfV6fwVeplNSTNgmkGwMeZEG
NfV9qOrFettM7c5cS75i9SIbKWjCZscBvdni7CxXXGn3W+6o5tFODgu0JhkFGQ0Qbj2cvwQVRSuP
ypGDNFlhexmMbhokNI5Gbvb5FlvUak2hfqZq1y6BRUN9HQT2K2nyIvSAcfR9hlrQLwvjfkxhd5YD
/Xlx/Vfs5+o18HjY/IYu7MXCdFhwAvv3qvN7xMdcR24Fjb2dPpErDfJQfY0FUlaJxgSOA5EsQsdE
+VajO49A0BjgthfD5oOh9yfECg/3+nsDmVlRCeNdvomtUbjDO13MP8YsQ0cyyDrPzd2ioxHoZXov
E+jfLExlIdSq+1BMgzCeM/EZ27x6UabYn/htgRkKvQ3L5iitW/LOYU3o7hVLnG6Pq5/8Q5zYGeur
UsJVZcUCchgqpVHDCFarozWKyQAlhLcF5ZCtOD+Q9aVNtZ100hqah4RBJYSPoASO+ft7yHblg2Ok
6V2r1PClQI7MiYWmbqO0pNrezTV9lX24OhLYtfOjk6y9SHYbNrxserkAPLXrTDd6ERAn4fJOB+gM
KfBL/+qstbfb4BCLTAAesgoAgUtQfNms5A+v57dG8QAe+sT7Wg8G+8KGzspbXdmiJ+zthMu3o/Pt
qJQn2QLq01E62pFN5eXJEXaE6ssIu8piy8MCrlUC0X+8/EVU5AWmmN2JzWkJSCy2Ml4fg7Wgp14g
MpjpNK4he0WwGHkoB28MSoNA5TUREdZI3tzvb3potq+CunL5SAoSZ1RPw00G/DK3lRmrB78/yEAd
0uvI2HkmS/V3Ce9YB1fqqiy9zF+qNQ18oiiHn6/xR3yRvr3faV4a2bBErF4Gt7x1QlMkR1Bw79kX
yTTM2jRq0dI3Wq0TxmkkKkpkFtoCU7GuN+N0wDCCHzBa36IEQWPzJypZINlucFb9cB+4Odl2Ff8c
527blzzMC39D6vY9UYcjJb2R70gcghh0z+vd1Nhc0NLZ7vYxB6ESerfei19Pt7kIEy+H35BYMhQP
NxPFZVMxmq3ypSW2PFka5bbHtiFQtlF+QortQpkvNxNimPnYTlQjgiIumaXGYoBFXbw9eUcU7dC+
C6MjZESQoZtypHs465bwKobQAKFMoeCHyC4Vcn7lsCDGW528tV2Q/yffioZO8HbY6X/FzoeA8UOX
5lUTAeqBO44lSyXz5k8dJ7GxdAeJBOxYyqxNI49z94KNmWw/3j8E79JfldcvwRJSExleyYhIGn3H
KIQMtO0xkxHBDSkgYeqsLHM+QSSGvNlJ4MZ5acXo9wSYixe72x1Omc66Hmx4N/MTGiWPYx/f3vWN
cuZlDPzGz5YYR1bfz6gnI6SrtxI39DVKdnsA6LLNsVsAElOb4XKIkFYXfugMEE3rhckkVEFpVk67
bgqAHTQlC0clx43LmYkOTGD/N20+dzqCohfmWNtY0pWmq0N3l/9wHnn9QxdCScgSWEL3gSVo+ohG
zmCi2sIF4gdUCWQ4sczs3M9qeThMmDdbHCfb+XhN3rhWXEzfPrMz5/cJHuPOjOxnFjD0scHLXAXS
Bi+M9iwFEkcKtdBTdXgpWhP++zCXSjY1y8OCArhpVUegKBvQnzb3RbvuzXomdZOrtWEA6vAMJAtk
u9A8ktmRs4RYkdnZ6yOwEMsJVpqp1M8YnZ9+S7ynoMIn3IqhedHfwDtjh11+bTVy7gskzglgovT9
EXEw0eabIAaTu7wTc+5htYwF7MvnYnEdmu4oJfAW9xD++snteVCipKj8MRgjTSvr11m20vInM5yl
Yp9U+IhDvLSZNMMCc0iMvviaJZLZGpG5Ea7OIs4c62sMqOeZib61NbUsmK43Cb5Rma0ySjHEZXtK
35p9C7WIjiVPS/NvckGhUzJZbAtduusHshav8YEYHOe+YlGYRkXcgO0YDlfZlVq7cV8IhHv/TM9O
D3kgKiefXUVVvA4k55+tyQ34U+zS2lQU1SbAytBpiZDCnvTnMj930PxtRY3R+I8KvCSrsR22kJ9a
SzMYFvyH/bk4dwv+TbILLKYeLhE3rquEKx7aE3475ZM1ry37SF7BLNgzxB1924ijlntdn+4UV9jr
O2XrIK9EJiGcwuxzBnVwMtw/XAnumw+ROnN/+14iSsqVvBUgqKBgsuvXYMVzpLd2m/uYQD3gcTPk
IUsfww36E2DdVprWqIxmzqpHD3RVqQDmPFZ6vDlk9e3aPQy0agCdQFf0zr+w+aotwpfVNp5oqZky
6fRNs+ngv4qB6txwcfDDkWutZLMiTJ048wT/MU4lz3jwkxOfob3rc7/12QRfSx94c+eQnM3LBVz8
8QRKaTL6kLBM+i9a1u4rt7Ed0nqSiLuQ2d9IH9JsAbM/shshCCFelo8hX6MFRpuSF7Yp1jjDFFRN
PODYcv8OWnZ5591RH1dIgJ5ko2XiY5atrYk9jX4Gm3rUBP42bNi1uPQx2yMWbLJnnFMTwhv0IcaS
4K9I+dutGLST6hoBYQKfr41GXwSxgJtlv+SKkkvG58Q9kO4GT6GkMoIfiM/MOQCfWieXF4Vk5Hg7
j7R4dPyr83ee/H0Hb+cSgJV1OOKHgFVwyD4E850FfyeFEV2+wkh0UEV4U8rg9BudsEkO7Z8/5EFF
GcL7KnYFWLbf6ILXZ4LFluSz8BSU6CQHcxjqWTE+flPx4vzZtO+OysFRJZX/A1h6ntK17pr38Yjc
/gDRvXXXmh1SqGngwbINtAqKtzBkaBdtNrRu8Ft3pmlKZc4bOpCXwALIYGMpdtbQTh3DAgaxOYb8
S+KaV6ehg3yIDbLTr35n974OHcp/Z/9Ma6NIZyuIXdF7N6OBvldAIwV4cMRGcG8Gg+MaThi/weGF
YKi5oPZnZn5gjJegpdAu1lBAGLSM42yIoIvFXF7+DpFmKsaCeEVM8c6aEHmxq6GJrfF9jGyfN50N
fOP8a5zcJW4xDTMzILPjL+WlfqkWtcLiBBc5tv5C2lkcID7xq7TNh8Xcps8I6LYiDqvdPu7rj2z5
lj0YTqvl5oUgsaapISCRJueFnU5hMTIrdhtak4UIezFwsocgejUwb6NZQG+r3Ylg0qx1P9qm+HaX
zaMRIm5t/+kckxpMY7RBFigRim7XTCblcaXvYv4t7b3vjLoG7yYCxCtsjPJv9ObcR4QIxt/O/S8F
MMNxhTFoX7t0I4kdhY2Oc16IGiVndTi2GF6l2uQ3weTVcBvrBStjaVLzfm4d4SjRKYfozynXWG+T
sEOzvZNF2invJJtjnWN/k5P6Wt+Jl0AGMQsr7+Os+EpRs8UfD51XcbJwqeW+VwsKdaGcxyLKirHh
aT3WcVFVtBnmALDPbFXhNMRzNrioZsAS2glWpyk6kscbDwnNahhh46WI+szuIvcUVQRQYEnoIgMG
Pech2XK1wvuuD9us7briNNujD7bxvsFqVzrYV9Ks1tbxqreS7KJYhcFucC3L6kLl+fhkXxQaDhYw
CahEbNeMtEGwgVUS9DTNDaLKgoskeq59qxHsoqOoEJaxoVBgw1edwV/JAHWtpK1apOygcUWlBHio
Twq6yfOaix4DdGENgml0tfD2rAXViWwEmJz9c8zm1g/++CEzGAHeYrP8UF+p9/WQ7+sE6vZytvTD
ahVFcwCdKI4wlUaw5tr5t3TWZNciqi2BBwynCsA4Od5pL+2YY2UMF4p2QG+JEv5SFfSZu/NZ/M/Y
Jz2L2/NdwZobcKjpEt3vpcPmNjMc0uaC8scomQBzxXL4ocHXav19xuFc4gUAtjAEXyPfowccRQdN
BLgPQOh7F2iMHzGf2mWQrzfipvKzMrqWOASscYiZeMBNI7odJjHf9kYhTAAvA67d+KwxeLOuurCB
6h20AxXkPq3xnzHLoj6fmQY4lqLxOvatbPZYiQxq8sl/TlRGqZzlPEvjPuRfTUHboq0m3OtwydDJ
yI06ol1BLeDUmaetzpzQlXUmDil2TwS0zrs/CvkOFzuKgawpjLRYgvUrGMW3zJd8w2kbuS5fvzIC
jm4rGs+MOw4qWXj/6nc5D/Q9qyXAyNlTG7w8OJfuFkzHDhm5vF7UtR/2SSWLKN2nActALoZawYj+
1LD+iBUVzF14z0DRk0hIltSE+UxBT//mCzBLlg0lJ3/u2lsi1pbv/mbfwqUCbd98Hu7rmerGGnEQ
uHqkENM8jvAAGq+nxuye9QcYq985w1pwneT7y0ehFm1FWX4wex2rQK4L+Z+P+SzIxHHOdlf6oLug
rdkBCogKzdhVaV1FoIIRJrKPogoyiE9EiKot0n26hgs2vlU+zfddtdYa/bmDnhwHCahfR/7JlQmK
y0mxW6a+92sKRR/zvyipY/05wSWwM2bPfLPjw9DfQ9ouGrqJLUTSYmz+irhfg0kjGY9NDNfTzqnM
ez/ks/YxETXd0rHxr4XpC/tV/mWycDJIplra/oYS7eV3S4htJpr+K46kmdttBsms3cQLgLEqj3Yk
bjEI/0FnngrRTSke73RIP5S6BJK/aWl3qpCRQGNnAldrFg3U41q67GVsZ6N1GaTLeFFPLGJ10YUG
S5/HS6/KlLYYGbqgT/pHaNy0pR9BY2o0Pa2Oz61ct+V15SDH6tOOzkJFZj0wIvedML2Y7TcArLkh
W59Ayub6tgmJd9HlkKbu4dYpxf6D4g2vDbLHxdMpYcNQuQO2mfILmffZXHw3k0jIj4vViKf+O+kq
H26hqiNssLrVXri+9okJPXKp0P/PIjJULFafnirdwKMGcTkmD/NOPYec4KU97+XDAKWtE9vlzTpR
5ruLSAR6HBD1CQqQYlEG+rThJf3OLPJp+tvw3KA/g0YCA8+AiESGb2VCxSuQ+Bog5L/xrig1ntwb
ZJ1QlPdCDB8rnCDnDrrR07qeJrHrF7D2rnJ3Qw4+bvDFaM+rBVWJe33vNMDms5pDB5IWSzIp+E6O
64QrmJE2Fd7XmIDbVnFIjIrITc63M0PUqCGnkFrvAfTGKnGO5ofoVQe9+qUYJ1PJK/6+S/tatDXP
iRIL3BY9/7DrtFeST+JWU9Wjd8tgnK3UIqdGIEiKj2UlZLseIAjZufn+GMb0Ochjuxlte8AtkUjk
S/SeOn9tWfwDt2T7DDK5MjnoPhfXaN8AyqjDHDOR7lK2L0WI3KDRQJBrRxHjrJITvZLEDfBUnnnj
Trd/U1L2WXhrG06AJro0xVfW9goO+N9CtVIul3F9vFG3GQmTgg1siF8+YCVju+gRrPIc43K1UbkH
iMFZwlg+ocLxMl3CzFonEqpbfCQL0Tbpfz865sSR662OSb6NDkjiErhnws7dIm4BIS7mLTdXm06V
aZjqRhT9Lvc1aEKYBGxlnza8AbHtOWjXFnX4aIN7y/DTC8UYOFc5CTRKOCb62/spRLl3LR3JLl2X
FeC9KV37K5RXrUtcQw2NQPYyc1AUGwbp2p/su5SP/XDlN3II+cjKed3hBtn4QkRD9xLkEKJuRfQb
IxUMm91bIxeGQ7X/Y6kFB+JQ7EbRaFZiqFIfkc1CZTXHmQieWGIOxaap91lKugvjrdTOU2LvsCAT
RCaVUpEjDqnpP2SbNZQANQcBypoDqfN3woUZnvafoj8aqI4WoBL0OwCfCXkCjPc+SQN4cxD3acA+
xnaDffsAygz2ivKYGn224TX5C2CRRo1/lrfqz82xpHRMtg8yNry3zI3RRl4YWOUo5JnzWdLT6EHn
jVRDEY/7Ifi5iCvrn2dQrNfXHGYUMuYfuvqEbjjUnbpuv0LnijAbjg5Iyvn1Hm1N9BiP5pzs8o4Y
CyNlslTeopyn7yN31CzoqA5O13zqQCOmRoxlPZJzcvdk+YaMZ2iCn0AVciEMuBgI8Zxi24nVBCwL
uLY0STwi4jViN5unmvLG+T20kF/0AWevpcRVSU6ztCNZGrNl8N3TTPy4HcvkafrUE8XggEHrJh8W
e4E01FJyzWAkjxrEblZd0i3as1Xy1cr47bfiIf0ZLPtFoe9UM2mDVFvtPgGpufO8J0DVGsdPJzjt
t3MhIrb+KIkDmMAeZGXlqDc/1+5YVSv1Sq+r4w/1j+Az2GxXAx/NvILSo8iV2qIyhC5eT/gkS388
iXWJk60h8B4lNcjC7Ax7WlJMcmYauegAZkea1Mi3EJQmOxU4AqHUtpi0SBIHNqmffr/L+Qd5ISg+
OFJ1bscnficbk0uwZuxDTtAaWP+FJ2IOmUjVb2dHNXUlsw5ABFf1YLxCl2DlLA2X1HNw7OKQbTQI
LD1a2wVLe9rTPFMkinYFdmMbKhygqcJnJKrqTows29NIxZq2WOhlMWfowcGdQnZS7PzGgkISiUUK
xONtbcMCKCiI801u9h5pESCa13HRlIv7JBTUmyVgXJsGwZHWLqR7zfyyEZ9xaq6fdJOiJZOaCToc
PW/yjGM6pFYXn1vbcWWC15JxxisWum6+t/8O7MkuysELs3OMp4ZVacGaPhkIkqvLqv25j5ax0BY6
9c3CR3fyzDxabG7FzZCKokqP51uGFqffDVmLlGDyJ7Saj5iup4CcQ8on6gqV+sPeCyx3WDCQ+bIr
K5VSfSRo7Shxv7/k/pkgFfJiXyvNJHBzaYvT1LKZ1/IDB0UcGNOrcEKvTE/fcb8kqg6bNhj8aq7s
4yYVmklK2ze4Hl7gKAzU81WoW+o63vQ65Uob8UD/MERwF9DT+n3hpT0qRciHDj+UBtVWxBjpVI/r
1n8tBRVzz7qhQByZBzFjXkKzOXIVEorLzycgLI90G+CgbkabYBlGSBe8zkO7Hm37aQPr0VoNX8Jb
7rP/Uh+MsSdJN/Dxyvf+0kR1iXjpvM/it2Gbr7ruHGX/dZuj+JdQ2IRk18lLVzd9s/89YHoFSL4R
Jko8gTpjMDHDt6ouNF7e/jpY6BXq4FzgME5cjMfzRJ0xmaBIPC1gZvqvVvc3t9MdxAkR02B2D2/i
seK92CcDpqlQxTANMXwO3ZduDT4T78EdCLoak9wgEgxrRrvxmZAtjzvpRRNoIoDSc5Lr7Uzm4Foo
y7qRiXTy4wke5vBSCZKKKzzSORxtY2sJx5aAKvARuRsw6pzfQDzPwZuiiTJh1zvLXs0fcGua4PFM
rX6SdR0Pf87DY4LgO8uEF4emvf9taqntfUal+4622YDODG75kuzDOkrziKu9lnAeP5UpwI21z2Kf
2n5QlTvIpAKa5CHS2hL4CLnOO36x0nSak+F0cXWQgzoDUJDzv4HErhN9eVU/jakco0HYYWKEkZCD
sIEcPi095G++W61pH4XA6yI22WbGUlN3NcMw0ceB+cxITYmuU/jRWltTBDbSVwkmfu7q8OybwyX1
h1R5k9FjZrR+p/5s508G+LpBJIKJk1IrbU0uSZwigNDP22KJ09t1hkkpNb7LWoCtpLXisP/7RpBU
5qFwE+elhvK32u+DGf1nMVE2xtWP68ehOBNdnjnnUeCEq4VUZKMvVZWII9koKAc6lQ86TNj00gIe
cvEv7uPe8FxEsthoXA/qiAA6jgvKt3iZ8lVk1YfqVHuqCXbkzxJkTzfjGnF28YFXNEFOB+Zc1Tg1
VoYYu/s/siMLlM4hp2/zAbqx1V++ay+mo+li9CKGPnZyTtmjoPtbGqElFaXmkzAzoQ0SoMhpQJsH
nQl1W7x9hMOgVX0imvcx+KFucaaXScs/n2bRVb+Ocz3WjOxJJW1zvUjl0Ti1kPGQqxgvC2z1P4kx
yyQHfW+bBAE8hKT5yIIhV5O/Y8LCYwLt7evUs3jRMdVbUO8xSjP6tX3L441ajlv8wWx0XHt/EH/N
oPc9FqGisR6iWC4z/lgIzHqh0bEiXZr2wQtNBQ9gnRQssD6mR70KnxpY0YGdR7cKIBjt9OkK/lyT
6sUy/VBl8dYI4tw1XG00jhfFXiUP7slAFIS1w/oKeYLX8g8nw7HI7xVauXV+VoofEkhuI6bn9G7O
KlEn3vvgO+QB7Cyufi6dM7gdohUDTMjdnrbbHPLt5a/smsQ/X43J8WeWAuRFy9jGLKjZHHmLMaqb
nQq2mfRs1xCCehihKdnA2v2Nbszyh+yIR5c6WpvO6z+ublQnb8wEiXZ47L/8matVQ7YlRlWGpFbs
LRdLd0i8tT9UpQwj+jEfU270Ciz5hWUZ0QbLz2UedXrAb3V9OkFkonOJHQUFuFsWlRHT/VMiKm6l
UvYilFTDrUw//eie+S4PjFwuAb1WCXOMwu8jU21UHkJO79DCBY9NLzjzq/UGk8y9v1hm3rDs1dwR
tq9NqTNgUcPExcn+8ENIMiQLzNapy9MEs6cRv6suS7dtUs8m1TaT7Xc7sV2C9HwuOS1dggIbIGrp
2Pqw+QJOjTOVYVw625l0rfrOksIgCZQGP0pXJrc+IhWlkorrll0i+4D50wiW59MCM0uXH3eQ/EqT
6BMzqKJAY01duvi2Ig63N9/BK9A21ODlnxgKrnd8GVMSUVe0KhjFLcvd88N36Yc0okSbqMLLt5pB
x8sev9+0/Zs6L/Z7auLMA7Y4aFElOoKH7QeD+jaXCuD3wpK0PxlLqYbkVZRS0q7BcDn3sqZyXLeN
ivuBieCHtGr3nBd6l19Feo0fcpTolciunU0ZGhy79Z7yIK9YD3eL9ILPNuvP8LsnX1vW1a9NUcl2
3pRe3zUiKqofu5vsxdSxQOmegHNSpAe3X9HHN72f9sESNR34n9DFXZpqL6N2eud7j9iE95gTdHh1
dkAz7smWosbKCnC9xGeDUh3dC+QHRJ/nv7FI1uCe6WCaCWXvobyEnKafPDRqbXKxMF3BFYJ+dLdx
RmKX5PZq7lzvdkXIj7t3DFJJM0AtEYqPuo8xd53V9V1XX/DcImhfdu23z9AzvwXoermA3b82BWTd
9RWKG9JripOcBJGST8kdr7eBTWNX/RS3y0VZJOInPuHwvY3TfKwkvB2pRqxc5484gubEHeo6uvqZ
BTRS1ivVMR90sZDUJmWi4Xih5LDnsWcsiY946zmGdes2owJgVLxl1eGJg8xLeIfZMNJnlwW+y1MR
oKnMWq50b09GjhbD86d+I91BxzIbL/VPe/Pg++kEtEHEkG6IW66F+W/AvPsv00fva28U/T5NQNjS
cvLErjJl4e+Nfm7qOasWv5fK1cv6nPtO4jTv4cBhfz5wYWSc8Z1oLKDqO+OGPvzlm2TB/g5Bin82
71RSbzI0dkAyW9uChQFbEWjMcmuGvLwRbFauCzTBNEmQ/v++rlY1SFCYAiY39gF0Nn0ZZZPxrd72
lyM2eNnvLEEDsV5TMvWjL0oid1SS73Wynl9R4YDiOfgLpooNMlgvPJKKoswOxJtoHzzNnRp3siy4
L2+6yjV6NFjlMKPgGitRflgpsjSD92tHqPLG9MkCsqPORnmp1FRcZL09KTDbvBPLy+IDbosnYTdc
B97Fbxtds0FBPcmv9lz3oa28k5y66x3rectDhfvYS4glxGAdhAaErYHrnIfax3KdIEK6JIkh9O8o
hEcB8wA5gkWkNkcda0DWH+5FCmWJrLPMRDUc0iXdDJ6IPkafuHCNZFrdi2CrJSjH5oDlTauPi9Xr
mec/+v+dPw8TZ+IynK7yXaEU0Ljj71vB662UzB43KUdjI3qAlZ/IUbrwnFZxOVPie0D4IT9ELUYk
wiC9u6bybmCILB5Cf56RY2f1xNzWUNThe9z0cALR6hce6NAQ9uo0EobTiCQK2iUKUhQxKRAqLWeX
82qulZDrVjiJT12ASl+I6ojbp+/SqON7WlSXfmdDUm79Ee6NUyy/HCMAcvJ4avwuPkjsx0SZXTE6
atF9Ab4T+BOsPfFNfst8kaY0sSA8iHaltT53jFJNMWWRtCyK7bRq1uwEE6EI/YYERyX03At+SjP5
lKmfvMqK93sXGRY3/hGhmeC761u1fXE1x3l9xMnCxaUVrjetIOnQruFP3XcTobh7pXKHHjczGHcu
Yx5bXjHkAnr5k/gTfEwqnDw66nI5uP10WRvWuKbcb5ZR169cTUw+JkoP7CDrGOj0blQ+87LBen8M
tyFsjvklIjL2bccO5Rx6sW/Ulc/qDzhs+kzKGpkCyIbvhIJ/6N9E22A4SdxmDPymhKBJefFfEgmh
vfeX6szkFzjU5ydNY/7JobtkIW511RQ3tvTdXj61ea7ByxVKndDSkdFBHimct5SDiWMA493fgIP3
aRxbn5JwCt5N0VD2vXQmWXDzIz1eLd6hQZXSh/qS66s3/6QNSfW9U12seUra+LsmTGNpNJFdYyE6
IoRFkIEvV9Tu99nQFcoqLQzL35oYX0ihJam1X1W77uvqhd1q5B7c+f6/ZLqBa2cChWTAnNuWFqSc
FazSQtKdpLNYJmPwCGA8tc0sVWz4WyfxcqyJSBmzCb3DbvJ8XIbsq8QOMz3V+ndUAHeg3VK+/HS7
NyrsjI8J8kYchIEqi9c4gZcjbqSeOGlpqBefqnH7oVNdVTeFkuqloOQX7UxSDp8gBw7qm5+aMbX9
UtN6G8hSFSwDneCc6IHZw2WzNIqq9LuqD+g/0v6AoNRrz6CbBAYSpA8KCSfOFaeBZL0seKK2SwTx
LV8l7ukIub5TqKHJCmNWRNzFtw1A0xkQbojjY1hRHw9/fQumwRETXYki6iXepHtqK5xMBGgvBJ+p
rmn4fsNH0hLlo+G7B9KkgJK40UGvv8M6XUC8LTkY0Y/zQJwZXFCL+6MT9VIjDyJ0/Rm2qSEluJDv
CjPPgMM2AdZeNRvTeGx8Nt2aN0MNLDInkinOJWLb77FHUtlX84pUlDtQcpooTH/YIxeiX4PG2VML
69Scl8lKqW/0yjH8yj9uKwru8X+E1nvsyiYibOyN9VDwLVeE9ctA2pVXLahSn2D6dfQeeMjkViBh
o1b7pPtgvnXcvsdBGAmfMrZZI1wt/PcarpANbWbPkU1OX6wwOSyWKxUm/gC7MbwTC4soy7pj5f6C
hlXlL+HQDK0x9dToHX7x62vxKVcIBLqeEXKj7epT/hPE/fhOvS2QKLNgGHaGXeQGDWjAzgv6CxmH
UM4Uw2qDq6laHjDS7ODAEwlpCoKKVPdGZ/epdnjgwd3CmVf3By1/XItWAeFyB0cSOp9fOzOiyfta
UNEjqnHDyojv6B7l5PFOgk4c6V/pIxNktv+9WaQ8HLO3B03Se6aOjbDsJoy2T03FFH4lPS0s8mHe
e18wowI+UlL8uqbQ3+ArsGvIvmfIiW7xBJW69P4hG3xsWNevH9p+9lswq2c/ioOG+uxIQNeT9Va/
Ki9oCTEk0ZcK526xoJUilteL8oKWFQvoqzjRzIMJwVd6ZLbD4RfHgaxu7p0cPHDYV75SNlTlR28n
eNvUnQlZUXU7vULV9pzkB0MAcIfIF0/MuAE3UKry/0zasqmCWt6zumNFlPBT724o4Fitkvr/N/9g
tKCerQwSRpO0hzZJliJQShUCVQtdTZcTY2nOHBJ4Px1YbeI9Bqw3qLGajLbCQZ3Ten1F6UyQOz2s
Hshf0KwVCw7aoRlXHPTLPOs2e+8ZKG1bvWmRHmQ4FjqPCphCY8XM/GYBhnyo207ciT3uBONGWFOe
e2hZwpJfmUxSznnL/sRCANRMy78yuEffPm351KwbMYqphe536RgLg4gXd+QGYjVB/YX6TXpb6Jfp
kp085Fe7SrqKlAtgOAFyNAI46M+tsk870J15wdgd7oyF0RHt/ENx8KRpIkpEEhEDUnpk3CjazAJd
9ffXCu5w/RDGypZ4EjjY7K0Ao3ZUkf8UQKVuAPnA0mEvUKFANk1cuYDKizwEUce8Nzy+bK6nYjG3
aM62bqVPdA/FQq4gCEvrfa5eQn6Og7GrED1HPXZsLmG/Ah9IRk0DRJ84/lHe1kgrsN2hICE7dfve
PtRCOlXaz5iCFLkYQa96gmGd3g+GamcJ/FChz+5+fyn+JPfsWtvyO9CjUsk++ucEkDcTO0OZCXjo
APYpSlfrzKsesJWknLKvGo3vESBQXHoDKd1rSyIHsu6oz+xgqJwy7Bg0Vbf+RxvNUFMHAJiUtP0q
qjJ9C5m1PuktD+bWtASd86EN4tPEetK5G9DGJ3uilHQZPoeaetQnYu+Oxrd2LnFML+/qRmVYbrBS
y0kDilkKTCaDSzbTmxt0VIydyYlVBeH+Hho/VQe51LwEa/4jaxtvhwQFjrFpLDpPxfyyV3zj433p
eQRGq6vVEu8SXQV1LxcsxJu1p0QR70f/+Di2eANuzqlj7Rw4aay0poQvawMi55MozhH4o8HB3u6n
oudHbAYVnVEoQQzf6XLCbPkKo9IKyzq3diO0jTYzkA/jnC//HvFAWkF03u3xJDDcjTUeIebLvcod
YltPnOzXVnOOZaNjvxjL0K2py+HA4LgMRnnefRG2Zp9ERDOryMgO/Tcc827GfioIt1q22cjOuisi
LgRrJcuUDRqR2CwUr0oXow/AcVL0Mu3KG+aMBEfgMFk0dHiMGtuHGNn6zboXF/TRbJfkVDIV0nyB
5bOPwVd1SQdXxizQZLghBJCn0eMf7EnvormuXBgEWN5rRnfFOKqLsAdlnt28asGuO2PCiUfAbn2E
I8JddSR3ThBeznYI/cnUtwlD5yyW2LF7kW1qb2Lu6vCqf1LpozK13QAYboaJShxY25Hht+hzcsFP
oTDaK2aU12/8PX4dZwahPtKbnPOp1UJnV7VFokywF8eTsvogMDUXJZHL77xChK3f+3mCgvNpRIlJ
qsSUkCTOKnmG7+0RSr2h33J+lZem022hS7LLl9bUDVVLiHNJyy2dbPXdYJvk3vwU9D4mXlkbnfLk
oF6v/5LWZsw//FFkoIiKSrHcBVfcJwLKNcB3mysK3vtMDD5DcJplzyR4IU66a5lSSgTbHzUJquaE
6vKUYQvv8OyMwWpiATnmQVuTN7osQ4dV7Jupm3Gt2fdl+c/CRY/kNlXCP49kKb3zuZ4HZUCWU7vn
N0WB+fz+hPprcjEiRPeuytXwI5sVRjhzLwOYCYmmDKP5w/2+y3Vebq2eUsFvSIJlhkYgcN0wl+Tv
ecl07D4jTQato9lu5h6xJFSjoytXp5n1uV8C3B4gBKptfg17nwL8TO+F8XEUkaxuZXhfRe52OkAL
hY4ihgZYJS+AQ+DLmEp3hZKeLT4AAOnJEomtRT3zAKVtuiXe4/mCoirVsAhrFqchIuJARGRpobfD
L1vO/cNr4D+/T3WZaWUXpKikWu+N6rXeZot4jwrf6V8BcQa2LeVtNHXKGwqGHfbV0cdhFBROFq+B
kmD1FqFwoEAXs7r9sIkirCZ0okwffr+kqG96ZDyJYL7o+kaHuUTuvF+jdw2jmvhvPo+q1NOvv2+z
LIdyNPWyxa4BtihG61chm/5sv0IaFx87r6Dml0IUxpxS/t1p66h4ZUlcCIzJxZPB1eN026DZAvJV
6vQDjJd+qFO/4JL7hbbfI46p3n5q90PkPY7Bn0L/azckQyGej3axDCQzQzy7bXO0xzMxLdKmWYIt
0CMfaUYX84w3Ex4G/9ULv5yc6FE97YkYbMmBZVBj17vdIyNaVtTadbw/0EF2hkY02ddQtCGVwxIl
CJIsDbqOk0JGBjcUdRPvBhjyBDZ58zKBk/J7W1hyqzPye95/7N0Casbo5yYzlKeJDbuiWBU321FM
1l8mc5dI3xLX/S4RIjNnAw8nZo+HEvqEXwn2OpqadxkhQ5jw2vZjHAvcqrE+LEyaj0Lth5S5u5bK
wWrYl7knLgDKppRstS+bmj9kz8fcLP5CC8weAeo2TRSHAaCE9aOuSeYFEYU+tQzTI9S5a5RqY68C
V7VX9XbYxbLw9k5MOoAkVH+kzsxTOvRebqo0d9xE3wv4zrDM5U9c3EmV+z9Nik9gSUwUbwkOIYZX
Wss3Njp2LFsHRAHpVyek28Z6e67ieOtV5q7KUT1+eAXMevEm0dWmra/LfugmsjIs7tCJXBXZ+rBd
lJLiK//j2Za3UKhrh8yCnP6Bji/XQhAIwRd7GCYyuNb+NmOQWd9ABq3CnbAJwBhXjet14/yJrEZh
HlPw8xSlmtvd58R0E8Iy4RHIBWAz86XKARCmJesuF7bUyXmAohyIIIh7cgfjfbyPrxZuEhMdXRJj
a6EcDTXFLxBc4BtpsUTbviJ7feuAhdaS+pHzuEJlFVKvSbPsW07zwVM2XRMf3taprPnTASR88we7
Mhlw9kRjliZJIpgSY5GfG5V7yAbynhsSCcMWaVXKwHqANPKc3TeEvImxqdV3fu6jwb6XWhetmbmf
fadDlGGpmJBFj7u4wbm0O58sEi43irmAtHGG/n/ZctcbKSxlODYNbfzmSjftOM1OEyNTxvrcpQ/7
huKVWHfF5u2WbhsWpMuOCPr677QYyfDoRWpKiH/0B4ZssqGNw9dZQocq9XAUV+N9QboCsiTrO803
alzOyhjfDST5LXCaAMf6iMOF5qGYHNWhyUZIBw0N/aXES2QpxMtZ5rxjB8yqZgwn8FPVMbpdX6J9
VLS2bm4ZPymRLB6Nr10V4J+wuAkggEOOS54aeYUqPhSisO+WmrJBoYGPbr3tuv9MWyorH3+qBxX0
JhV2atGSO5HkHtpaQ7mQGRLoWwh6xqhlnGAv0lqyGQIHPNWUddqS3Csho+6u6CcLwc1sTT1jTQk1
UTUZYU1Ruwb04B7/BX6BQPr6MBju4TfXONUrkNtOEmnk6I40+PRz5iAPErhvhZlwM0cYH0fYpJJ7
4HtfFETligDVmSMGsbcDLSgtxP+gqxMFyd7WFXbcGzuQ6nh3VIRm+xa2c1UpxdwrB9s4v9rztKbl
Z5xuNdVnxgx+w2govUyyvdzQq2b4X4GKTcohj4wZKL7+uJz2VCCVUqJV4kSDf/LM/Rmvkthy5/Gi
T2EVF1zPugU8T1/esuNpVRPHj5oyYpPk6Jo+l9NlbhDXTFfSypYpiSuYCGCbIlYWD07N8qr84lwt
SWQqt2IPx/t6OjUGDWirRSDtDEuYe58Pjl07cpW00Co2aVe3aJaFEFGBZZuZ7cvAws3lMQoqINLv
je2j9EZYl9xSHnVuABZ/fx6N7htbg1rKFNdripcBVvCQCiLR8KruLiCVhDz3FzlrLbRXPmJI7BIJ
TIKnaIZxD5ULyX/51YX7yFTGwmYhUkxQ4Tc7Zw09zdZdXV0evM4J7IfPzPGFCKriRGeI7o9p1xZ5
dZpTdQHlj7Nu8lHi1FMqEJEMHx7mBY0Vzy1ACjr/+eMb3/0e7nmvycZxNkC/oU9uFIboC23LLVdS
aGvQb7luhwZjBXgHghs80w8rti5gSomr633Q/AN/tWvRx1flmYq0rp8mmQFJjfxwnrt7SaFLzhSc
SMTyJC25qkzhta0IdI+6SHwX0OIweEIK/qDMakZf+k8jGUcKzR++676YTIiLftsZA/KHnGB9a+jB
bu/sXo1/B0B8f2hj45ME/5luHVVrhaXvExMtNeIQ7gEzwcHhBFdEd8OGty/XmU5FmJYKvWPgHhxR
x0kkYliFVG490LwmjjXYRU9puvBDuu7I7y+ifktPf1/V/MB7uJAJ9FqroNR2yxHHKZ2DIC8DoAMl
eVXHbuynje1BV4B5zv7jUmkGxnpEVF5mKQimBOQBUhqZtkDpjlGa81kNOmzspzC7ue+m6P48BEfP
GyoUXoNU89eItqbgSdq5r1KWcNVk/TxfsHNgDFPn4kJrS/b4eKev/UwytdQXBeCrreO75vr7MnKP
x9epCmhDnqcbvltk8U2aq99UIFaQbfNueymx0YckZiwuE6oxuqM8SWChVsUJzPX/xjFqTDN7vmrc
lVAy+kO9FmBtNdWHbp+oU9roO+WmaTSEgJvL4/ZLKhwTNJRvIuoP23ys2oCOaP0lWJyPN47XnOBO
T8thf/Pq+iXOw4/A+eXZOpgUcBNSwhPZttRZSeQrpGVmX5nHebE4Gtsm/otw+liGVQNHGDbn6k0T
D5rZzcOt+yG04NTYiUfhuNzFC3td/4FQHLOaJr9DJ6Gp+0lL8vSQAlV1gtTfyzhd6yTpYAItheL4
8EGQBLXN0owW1Od6hHHOTlKsu0mk07Z2WwA4HCWe1S5Fqi1ZmMuJo6YHSAmWEDAsfwTjmBxZtCHY
tSGjaiZakzejIe4+sihhllj9AVdqmgUr/BFiWSRDRqOkl4507c01x5RUvQYYDLTvaVkOykZ5a0Hi
907CRjZUYSBdI3Gm3hhVOy3/09bjcCjKspIDPaJ3DpuGrxul6YdQeMuN6gvmPc8IPxgyeF90ZQio
xtW+nQKIog+PmUAY+mAEd91P3BQHMvsyI54vlrP1DIZecrSBnn9YiW1DEs38euwdty1Y90xadRb1
+DCvZiJbHY1Rt53T2ad8re/J8xBbXByOwzC4mMwwYlmIdH2QzWkOPZN7ydVPELAY+vt7iuDWt4JW
6M/7qBZWz0yz8J2H1iWP+deoA4dA8m3VWfpaGg2bvsluT13mpeYLp5ZGFmY7vdIcPMv8ZvImC6D4
9R+5LJDlNgXALP1WYZ0XX2itpwoQkLZWB9OlnGAfONrJ9AGt6zRbaSo5mCE+SjgMYc5BhVltjBfH
2Iaik2QqPnAGbKGrVb9eI38EnNLaK8zQ9pjSNqCqhKNp3BFoPbeoF4DNXjy64jukK2+uqwLxaxpP
RBnqxHwQKuK1Zl1AABxRIWtldhNPuKTjLrjtH0gcS/jD1xQb9FJobir274wKsOEv5O10h0vlKP7M
QC4a/VUlbSnhulv+D28/kecXrEx50qCvAW1nTmEY96sV6jEBT/zx13T/D9r+20YPWHtbQ33btGqR
egJAgWO6te7tY7XFLF60SdInM7K1G65r+47kK3r2G+lDDiLi3a+/H5dk0a3mKe69/Tet+YTf3L0u
o0K2tbtBBrhEPk+YZuJxMi3Oq/4iHURZTcZm4fQXkqHEDRCO/71q3o/LO5ZpVll6SHEj0CNB3IZ6
LRE0B6q6/VmwfF9qBVt1H6spc2MHAo/pcmemcPa8rGGCStOz24lle8ZV32ye0qB+85zBGVKpnx+m
sU8SBn3G6kkWI3g6AOXvQ3/4Wu3nN5aAtEf6ig/dAozLa33o+7qnghlT3+L3ps8s15tvaGUsOx+x
gIiaPgFUblwxNYCAWnZkq8y1WtPIduWucaxmkhboyFUe7+1asoANPt76Ylo2aWAswuI7QZelfLD2
7HvZ0yCPVUptT7W1inCSBFs9Du2g+BgNQJxpZiCRBOPBzoWlqJw1c7mguR+K7+bAHYvWYFnHP+HJ
CcZ/8xh6QOpsfDXP7sTzp4gTr1i5lT1+wyB1UnANc6g63dhCNudhi4arwKxXM+fB/IhdxHfcKe2w
cQ8a0qI1PPglficNo/KbQHZ/oJjbHXyUdnlvUd6VCXeaJWlwey+L+PIdBG2zcZZwcgCtVb4yU7GG
CXkNlIlBe4fe+qcxjSvgg54f+HhoEwPRGvhLC8PoKoUvQIq0/OAOR++F+hKdTczyKBdE9W8/PUZe
TrchtjMGtZk9DRwbGTEykYsJOdSXGXNpIetdOdsjzPRCkw9jeduT3bCvFJ4NUECU4qSU1evIltGy
ErvqUIN0rLsBfaGZa2DuvzuHqzulOCIKCI0DXu76ytOZPMI8u0uRr2zlLa1G3ork+3i6eq6Bfpmq
GAflNepDse065EzP7hZhMQP24koDnO+e9g8gpBXzTmMUsKLZky9fh6d38zJLU66a5l6F59wMOaEk
D6krn+JtByMqXRmv/RAd8nj4zfMfkPWpShTNOK72Nkwni2ZRcD6OKVNRvSnRys1S/VJ/AnB9Ux1C
rec1IdF9rLj4vYSxc1gtfNQhxQiivuCurAWrFWmr6yPxh+j93ILU2RohdJS8UepaYtM7aouysWS/
8fEGjzsLfgvUeUuNNwzpe94vdDi90ftOs6u3xAWswHJsq3QGw6o8rhMbEvbufRn6UnoqL8CZIhyy
qworERB75xlDIVqRPo8kbe+8sJEz4riulNzOUwe+oONpIr6tdRf2z8NNDjkknH/5EVcNSqyjd9Hs
kxk+RVayiw8RdARGmZ6qp/Dw6iVnTWVRevu26h/EImtyKbswXOAUy/VsngUtxY6doLuOLh/yX1mZ
iehLBD85KftFwBKsWHT/KMrQslhT+UGQwZadfR9Cb0tA956ZHn1ta3Aza8rwB6pmM1pywNp/6BRq
EvedFcJGd8T9kdZNxiWFtUViMOApYAsmy2aT1aXbVUlyLVYRnHKq3j+lDpt2FgvvxeMCO6QF666K
kOSPrpL2N4tb5h2WwciZbJy/lJt90in89wvcWX9367Yjx9pRaKg9cfYW+E/vgA+sGqu7IHMSyM26
jJ6E7oSAEYRqQD/kn9unU3CvwAHt37EL/G8mPeFX84tQM+Q49VQHTrqIQqGwrrgQjgLFu6QT5duP
5GuRtmFIyxxUryueGO44iPJvro1BB49nhV9pL/PpmQPuzS5lHbHJRcjSCp+uZgwRqbMLWesLgtvf
YokAvpB+FPeyL6TiePMekZuOKraXDnLh+C36t3eaIlojdsP/hogkZjZvRQnjdZAiM6H/A+EvDGeZ
DMul3kFgw+uHzL3l27UoqBCh9uuHjDeHJqt/Ag6smOKdeCn9swijZex5z8r25etNIUJHax4nrDCK
EmPftXO3TBeo1scnuS++RnE7l2TpZtkvBad89pHb5O/3pWiX7YdSCsdN/3tiW53PdwPxJsyd+4E7
zpZtLu04DFL0ODlkqW2EfOhrXKlMzcQ3WnnDFBDPzCH4QQwGFv8pBIT9BRCkO95QJWTs1jGweqyz
D6QQ+rRwXHCe7XHNb4zADHGjS7E5dJEzsqNUaCVBzWGn4tibPCUpP6QvSQhsQIlgxqx2CgqU/bEs
fLVmNnWs/z4UKGPu32VoKAKcrmGLRCKX3tlSyzmB9xiMAL+0ACD9wtATniYq+7QNKYKGYMJ2Yhcq
8vPFV/8IVmpwFJx6/9xndFk1aAy6+vhnlkbkxhnO29CZzEau5RrvSKNSGWDENEYMjJywMypPic76
dIJslN0yYuRK1fHL9HxsF5Df7zMquXkcvKMbIy8WbYXUni5kbD9kUb96CyY6/q1eKd6Uv9qAAY2l
P8gRG7oDEstPkMlCxTTnmilUC8Hl7FFD52rzHLTrMn362Xq5GZ5IXUqOecsUSWUtGiAcEvx+Ht5d
R7pWCFzskIm4nUkc+czZJGYaktdX7Opivy6H289YJ85WnaErf3AWSJjUnIAMAwC0QNl7/6hOtDL6
vUBPkn4j5BlRnZXkHpcZv0lmP5WugKJ6Ifan1JJcBAPrFwQMimB0Yu5RujWP6xqfWsYUY/UmKJ23
GkcQeFk5/ItpipZKaHCRRvXtDzoQuaUKLEgq9jqfTzSxlCtgwxevK2Sf76Yqls7VZCuEiiXd1ovP
K7w3P0Jhl7B+Ul0c2gdO2828gujORosggrn1oIgb391eNvwwljXtJEn0eu4A5ZCPIceB+i1+c1di
DTb3uVnfu5rzr9KkSDrpmUBLVjc5h8mCRKF4Z3AYsWgCmn40yDYAG3Wxxi+erK0e8d5YjwoXxxAm
ECxDI7iWok/u6GRcUaft/JByqJHwsusllEP0qCpQGsv6FBOJMmMbRjO4kKNmcmU+sXXUHIgPepKz
xCuP3xakcbdqA4KrB17Ng8uhHl86oyomSn/e+u+Lxz/gSaZp/1amveekIbLCmwXubDNK3AU7hRFb
ndAKU3c+m1AcMJtko0O0PaPJOAY2TbZ3KZeRBbpt6pfHtFqEqKL1Ka/0/ruLZb72acQuoPoNKbWn
VEhyY/sZltpO0FNlj+TYVOfzadN9erjSGBoyzCZCQPo/SLjqPr/KTunLw0iaBale5TIHt+79KlSJ
5uUVNHPytA+pqY4XxfGUmP3giJPjjDKWMkGwGhPa2q0/DRwti4HCZXHjwueiGBCLdA3RFSnTdByn
ujKSEXFD8TB2dTdH0lJZGOZtRQWdBk/5LI44A+VX4oR5JO/ZifKkBcFWGbOrLQ6zzL8uUoizpGGU
1AEa362ioU6dLRPGBQsXbXw1ZeU3vMNouZ1p0mtAFrQ7SaaFW2IuXHDFHQMumx4V7URFURKGlmrQ
h+rTVsMG+MDEwhvI9rS7G5wD5BZfVARYhzPx5Jft7p30ezkiPdU+SwFDNsOPk9bpiXwd1uzlZAtP
UQ+q42f3dYlOCNGdx/3WkvlEnWj/GmtGqzoxlqL9F5n1uRNNUGqt78SOenrgYWsnNhH6LCNgZUb/
3SIJ5aMV4jAByREccCNvgyV4E/5wCeO1Qri7yKZGGljDd6b9AhYOUL/B1foI0cSpv6KnTWSQ6hHY
agVGAGi0sHnsjRGu3o8uD+rKNH0A1awR6Zq0TaV1e3eEFzHaezLOzwAX1DO4D1bXtUjsFP2FVDwc
1afRWRJbBy0SpEfLpUcen5G/OTZBo6dAE4ABf0WFV+m5R/FKGQNt8N3RPQw/4QJbrBoRJGM8ARdp
WibguwxAOYvDTbdcCjgRJN/T5yUBTM4ZT7KBjx912+gYtt3sTA9AKwlAtD2Il5h2o+JkbYv7z7uq
KhGTDYRngG6Rsms6NWJXCHiQOHFJgTp+0WCanx7ub/dJtRflsr+IOYS84lwKb940xvw4EV4KZuKh
oosKQv22L8MLLrK3dBJQ1hJUCNRr/t4v03AAPym5uy6GG6QqsdGnXL65OMmWR47TJMUz1jo/6iat
UUoTPcwL4fnKYassGZemuAf7PDbhjBa8fJxHN7E+J8MrM0uMN/K/mYwijqbp/BG/ZSj8ouMtUPi0
kYP9eperZ0/9C2ODmrugCr+K5Gvxbl6GsCAYpkpCHMOw8SbIGfGKBewI60ZeeY4KV+tiiv4S+YBJ
AmpN9yUN5Txn4HZVkRZa+/jNFRtTw25IdPI6yLvTOogXHU0zZOd57age16YHVnqJ1w/0SqP4YQfU
BxpZ8Xvrfa9X3KTYp1OJumZGoan8vdv2TuDM2rrdgxf2LCQvRQ+M4L3nBeVojaGB9ckqn179SnxP
t0fDFS6XeZmommLHujfOJUoxTQc1H1vt4BzMWekHgj97vmWzZPJ6YqKZIzpXSbF/ItxCYHXYDcfM
e3WbOhOmPBiQm3YXx9YEdKkyFEGm8fPpkjGP3NkNlU4t3ifkB6Y7WxpNwj14qwxna7CsGep4dWmD
Gb/XA93pMCW9esYC5XIVvMF6Td3ABLNypT64b7QYlJRUlQNdzeKOSaG4kfHtpoqqeWlETOAcxlGw
7sYEXfur1PXQt89314xk3gVQUlGkwITSfFu4q7QWykg1r9wB1qekbZZbf6j91BGAS9T+tABaD4bB
76Itn2yCFbx269bH0uzB3VbcHX5vOQzOakmnRnmE9GFm2vXr5KXoMuZrMl/nESbm5DBbWu8Fycp0
Avh9sk7wqdoAXGQOHdjR302EcaRV5bQ6h2SbtmK1uCtINoHfTREasecUtjiFbwhNEp7q4dyE2jU3
wQjWJz/+aVpATQ0BPr0SuZxOy9mpLX/0r9Go2JJMOpYRvHUlvIBAfPNHRqkvlxnFnrJgXdzJUYoB
009v8ivsgSQdTkvmI3S3KMxKbJJcAzkkUIyhdlUyckcXgA63muF/aA+jqBqTT+gNVqJpT+4iu2I7
FDZFhnxAlou+z6zfJZphAi6IsRoTkP8ds6BnA1LED6ndrwEEMdkezLn7I/wA1XgMPklG5ia6HdPK
2Op7xRXT094sLvVNlGNWFF7Pp2gg7oOM5xn+s5psn0thy42gnNuUjaDA8zglrUdlQx1QNC+iO9D9
y1orya2TU/Et0p4sbvdq6lCKs7XTuu6o5Lbh62H9+hhrasm2waxpfRgrQPq0ihoZb/ebfhQjgmez
ImPpab9k7FQC4NQ5rmOcXejPitBiGdsaTZcMTCi/mo8lvWBgmPdfPN6VI923LglfDuvtYfPq3l/0
kuTzVoz2JYvQ86dxbYsmS97vCs0etkhARABDZBhLO6I1mTqfunhMyzVHe+AfsvjObYUpde4mP/v/
xHMSDmCAPp8MBq/akpX8uPfkbLc/aKDmZkX3+JRFBn5ztczHn4O9oeY1DxXAecUjRWpVU0mMqkzM
2mCpQh8DufTWu8iWZs1sR18h8O+ChMmNmFGg75EwGcWe+bQ3XjwJZymcAl2vpfCi9tSgg1tTchbO
UERCa25KY988eaBsAIsJ4k0KMy+AFAnSf7TTCe0FQdLqfa0ZVDnZ+OSEp+/yHcCU2HyDmoMRcPkn
nhlwnxH9qKAjrfNEleS4B/uQAtwcoFdmKg1e2k4I64UA3eEsPbZOStiTiepfUTQpnAw2lJHPA1as
3tMywzgo/xlUppHXcyie6O4dRR36mpfVEWwr8vpTIVihro23MiiSoMdiIGnjrwou/lPYmO7Jzn+f
3jULAir6nzH7vulBCG8biRZv/GV2/EIDJA1wbF82DaHPIEkj/QBXhzLXVDVkc9Dspk/gek8zK85u
0ptQ8UgBAjmmlF6CfMKyyDYTfJvBEWjZ9KvM8S7CKio/m1l6KBvm74cxrLFTQyW7uQWoNeJjxwb4
iER2fpAezJDHSrA5dyAePpOnQklKrsc5N8ofIU52sS3+1enZpwpQzVTiUVQ/shWeY0C0dIWNN/Zf
BXBZD2buz6No8KN1cZRprmsGSHvrILvtjFyYXmO5bR5BJMZcBNrvqainSEjm8xrVlil/OS1+WtjP
4tUr9csgEHNfg7UuWX76yYDlBCElPU5ZBRN665eLWCfvEHiZEDZ3m/qiLyOYoCY887SXT8PpLeyL
vbqMi7GZd16NXk7qi2oJMgMGD/KdMpuc+McFIIEapVUfsBvGEWbfb07DZAAk0+1/s7mu7dP0fU8o
chV2SQUQAb/aXrWE1xOcS5JigUmlXa/3nA2y+RJcnxWy8qCsUtjKHWW8LEzACFL30u7PPVJ/H7qR
/Kyy7uG3ecO2+nrZeHuRscGGLjho4INUNA0UUmgO07VrGczZM0ml2zgaODRmDcP4bmDUNkBrElyy
qBROxdOiOgvnHXBeP1BTOuTFUxgxceYRkoSqkOxkMrGOGqybpEoBOqN8UjCE2L1EV6Xb9hB/J7yC
5DnXKux9y21BhPCA2WTZA3DvjV918lxukbMMg5fLO+3mZjx/4vdYbRMsvRARYKo23CqMxpFFXE2a
1kFwgvz8u8tjdg+05R17rQiYsfmTjRDi4Tw/Vu9CCVIwq8YJS6AJypVqky27vATiBhyiZVff6E4f
IyBcJMQ8EiTHwqaBTTzr+yrwcNVMaJ96opU1gje11hrV6DegXTedcPvEhdd5BJrM8rN2yH52sBPY
Ip/1vpss1oNqyuz6zDMhMWymE7/zlsJifXrMho0gNpZNgsPT76ZJzPBANRQ9HRUfDM92xfZj4cvz
GbQomJvEdC+MlvzCo10MsmCaqz47PhPZlVRC0JJeKd6iRarVhrHnU7gkB8v0rh29n/bhtpU5wqAf
dNJPEjfwGOMgzmlY0y5HgVxRxZ/ualNMMpIAFPXxqNcVM7i3lAqdQ6fik8h1URD1LSPcUk6h6+jU
j/rcRwwkGHC8fOtQHiwDbpUigeojWqPJj2MijV9TTlw8G+5ejjpEYo1X1eIRv/rxZRzoClpq9nEk
gd4FCCaKprEnpOJcVRYhdqyq/f5W3Jo0LGm6HtuX9IeEHCca5t//8/HPYFXaEKOtT+laBeFsSjSR
rb0ht2QuhggW80itUR0iwfer+h1CCI2kFBVJfG9ihEnjgsv3rnnp2TBTneWr/WC8Np7WN2rW5+MX
YrK/BUD/wW1Qomzv2NEnLeGDL9YtkudZfxwdHnnOk1AR0f0ij1LARa68ggMsc33A/pseug+v/VoI
hk/rFNfQ4Qw9XVfv/D3HsAkgQWSxrTlEL+RE8AWQFuZVMP1Gw6lADmp5kmlJWf86PmxsrIdN6c17
Zq2LrpF6H5qv0ZSL0QMwT5y47zzFtPf2LvvEdUZ45e019s8LrPCPeXs64q+84Dpj3Pw9/Hcp3XWQ
2O9dz4lRu9xxD16kVPITJpLA9gBcxWYuzYJYLi8P+2pWYO3XbNtpvkthsTxMi6/6ahRySrVkOxnE
c/lxEoV4CZMG+Vj8WPYZ45fy2ALRrNbBzKhuy5vuemqKAIHJXctZtd1GxrM9RQ9bEieyKeN5YKkt
5Uz/Gg0naVH1He8xF+/PyIiVVrenJ16nVj3j3tCFi3P/h/HLMr7Z+FVfC8pqbSvT7vSXaPWzJ61X
d5eA7hVHE1D3gSaw2vQnaHMwqTuEx5i/jZbonbCJYlnWPbdqo77UuFy6B07v62Zf26ya9DyYZ+Ui
3hhtkcdAR1XLOCGxDlh6RGh6AoZ+nFwE1GjLbdBVRPK6fGzAmsClDuSGBg0Sj8QCkGW03l0f+6T9
589ap6bzpxF68wwG11K3uGDKfPnSgZNCpAqytmH0+RNgcvrg3FKgWHf4t+9xMgqrwRX/4lmkn40W
Du5geH6Vs4rRGie/ZQpSvn6wSqfAODqme+3Vy5iy9K0BwTPmMA3CIJKL86TL7Aom/zvzCxgNXdtK
cu9mYcW4KnWfzgTbB5bgglwNlD1UX4A8PrzG8AjrSRl6SxHQRBwKlZtoCt3VH4/dB0sWGGo1WNna
/nc7uq83fsiA9hhcH74JzKEh2AW9CiCH9hJEtzOq/gbw0pO3tyoMPSAfjjdZTGC5QDUiPFFZux/P
K9WdPpITdr8c5XbdappHTGGiAeWWb+kK42TtoWi4fwNWCWJnLfyZou/MZF6OSdHwrnvDK6U4AUky
XmNeISayIoJil9OdC3ihAAprsTjlQeqUZ/p1b/i/GrsiFjUa0RdyulgLn8P7z1sYGELzeadjkqIe
yPkdR4084ew9OFA5GC6dQx+C8rDij9PdYGOkSHw1yeSXkVjyy9dSnbTyVbj+n/B8cMaUPGWkGzqy
MgXX9D+kxo8nAw1EDGbaatyrXlKVDeaqFEhKeCAm/xbSOrB4myKk1E5rMiTDnfLY9Ff7UH8NN98P
VwClKKZ/opsbpfiLvz8p71pXaaDVpzLD2e/VoIN7pUc/IXHTJUtsq16v8qOuuouYxKSuI6T602E6
0Kh8MXqWqjLYYkrWr4AHih2U/Kd2WrkVZdf0Unem3o7MbEZqwoqqAUAlq+V40POCgJ7DF/Ee8/2K
SOnCbAKx4HoWC3putFpLRf/EEww/190+Lr8603i1lFEJihDuCB6xEP/I13bplhbwbXNdCe0QdBVN
wQ5yEoBN/5bgGCfD6oPfwQ+uikfKEHh9OLE5wIjDEJ7ePk4NSwF/UZg/t8a5FprChg/N46BsKAOQ
uT0lB+tBC9EXnfBK0fe78MkcOysqP9+R5Hb6eEe+gTdgIJFJZmga5cKlaktKjeu09GQzbpw5awLu
39Lotq/XBJqQ7sK/2G2G/z4l5xGUB+m6CFKdPI9AeNEiQ40HVbxqU9EZrfZOXTASDwUltxnzYnCQ
lSgVPk/eVE1u0vuMFZ7vG/rCD2fVqtZzO2+PesqbwNda0KA93ii8rY09jyABI+h4wiPlpS+1bNCc
n0MgEiwXu/fl6XWHjZSjc535clcnJXjzozx2pGaPMTeyEeLqZ5c/or2YMOgdcITWQb2WdlMODC30
uHPeYiCqH93bpJB8ARLhEfM5+Z66eqbbXo/XCLn+6ZW+ErhB6tPVJyux9HCtM7Vb5TGiplle35PD
Pk9l8neoes3OjL5UAGmfq3noIiwcbdan9MOkfGWQ7x9vnvriFb77Upy6igrAuXSzV1rzjkvvulP1
B65SKDQM/LhEsVQWwfl/ywm4ZawPYVo5o8nP+RAqThphNih2E5txBm+dN5bPtR4oqEyk6SWNgeRa
mIwa8yJKzWl4woans02y49ckqShmStPoYJo93UuXZWy2KlRjffbgVqN4/+RXEJLiryJzbaUL79w/
GJGYTqT++Jf4yp/0KRn5V1pyB6B6gjaw93dig1jBkzOSj/P5LqEuOlcAAQ3z3h+Xg3R6ks9EMWkC
z7ZvZxODKNmIZVgAouB89/x60Tx8bv4/yJeYqd5GO+yRq+912/HoU1836y0vZHpWm5/h8I99Taxn
LuHDxw2u34LlRwq5agIJrwLhUG1OMLEjZspguHo5ALcyfhmvVuivV0B0A2HDjg8KBMPzabcJU8kt
L8iWYpFTtZsvBShv4eUhwO/8ydS5IzUYp0kAUhVjErbZZOrcBaKqZyVlg6UYhVA+nk+fFsot7nYd
BYBjDJJqMHln+UZ6TdN4UdaqIV7ULReGB+7nO3K8CNpjg9IbNGLwxzc6SbLeLEZoo2yOJ4rrfQyn
+18qR/5FrXqWamxEICq1XhXgOkjLRERa4yV4VCIQ09wac2Pwf8h1HNxMrLOrtM+MTt0M0G+Szaft
vx/rBMWIC90/pqDYrlWl5RsRXN2JNNfW6Bssz9tcyd76nUf7Q5O6alkjuhyPHb8TEJkr5HRMwaNV
SRXkQLv6TRkpeTJFp8CrQiM72g7uxXCDg24H1tWY97GabzK9s5NV7/dJqihD1knCMJ2jDTynrs2n
6le7uFaw2MEIIgrgirtKSWeM1CQw5lnqLmAjRKLXvVWH9cQHPZuQz1Gvfz818/uwSFUYjS6g8j/q
0Yz2I4LwQ7QLozPk32g2xPJOk9nMKYnX/tlw/bt1OFMfGwDokj9J3hW+xKKyg0DODELdkNrhaOkh
6xgYbZwQej+BsVlQXalmb8RLcxcxWoGDwvKjTeLT4im41p/fWflo9YVxImMreRBb6k1rBJga2ya9
rAZA4oZD+gkLgtdpaeF6YHW2LZFL1w3C20nTqvJfNXzXxJ56yb+cLRXZ7EvI2DVuQ19+S4xUtRbt
CXoB3qsxjLy90aRKzTtfgwYC1qFx08Qv9PyyG8XxWh7z9RPOfXhO/ShnCjL8NjT+6QAfrOy7VMU8
pVItI7VvuT55FjOU7qYqI/Zwf2A6Ho4gt109AJdncvQn028ZenNl2dgxbDX62zzy8PSo/mPcgj7+
MsLm2SA844arycoa/XPvvACvs7CcUzsoAQuMlzf1PPY8qHRx2u3dLUFiXYzZyW+T+L1Gkc9nMjg7
AYS/FJU+/g1jCaDVricsvx6wZb1emv/0x7Xtx7HFZmitzYBahvdBIy9O5K8K6s6kppsiuEAS+gOT
OtDAGdy/qW1MtasUXPJ08GvAM0iF75l+CxJevtTzd8ds+8TjgL8LdIhJRU9Nr3/74dp2D7wV2NTp
h6ARicN6TG+sWLtOxCklhfMOZOa63/VaeWRYNpmgivkb/AhXY1fGeB4oBWyVPfHpjiUprqkD6PpY
6pEetE9NBFo3VOew7VPld4waKNthzg+ncjvReggAgEoWh0hFoZZiCE1PmJiOauxdiiqdh2fBxQp3
vrdcOu+uHxZsRUQ5vtdleS6e2LBnyuCEXQA5us01Crnzx4cVAvYOIXYn1r88o6Lg3Z7AsZL+UVPD
icWRHptZQdFdSetoyBgNCUNxbnbRfxqNyvgF1rtx9okNQSTbbL6A+h3jxBjUflt2ARTdeCJN1OSp
Ncj1Il8mvlV3wK7N7nwxG8kHyDGpn1nYL6Co9PQm309CaKY6gpTRdXZqTy5Ynm/q34LDaZ1easSh
fWSV87OMNM3k7ExFWVbmRym8e+UA/wU9CA57Wp9rdFZQmqzxZe+iFBxDsZPnL8KZSXRwcg7M8/UN
4wT7WNiTogPpj/Epjis24rqg/ot/wEzwKqa1CUtybdVdSvsI5aHs0DvztdK0/nuUBHCaBNi/oRpF
uTnGk3vi8sEgoDac/BS0l3Lv4UNbq7k7V9cFGwzZUSV4CT8OXPN+npcACqmXOd2F9lLgT+wnhl4y
LJFG490eFNZnakEGW8AEKunMEhmvjQNPyBY6QkArgTZGVAVeP/Ma9uU7eBKkT+zpwQYq4oYjx9h6
IkzLYYZQTZmTtcLJlZY7cVAR2XjFvIVI5jiZBzt/Hvd0FuYpVOuZ29kgnO3Lq6e2qbYIH1576IZp
YqPnm/EfInsbnR9AGbCLjx0pAPxB1/eYwh1HvuTMojTgQBYJtw/OjjnKWjSYgY/ntEAyzpdTAmVp
UUhVVDStsuRGBUExYhfokgKdQdYgrJn66CC84wwwAgs2kDaauW5iAQZ/51d357iSNHusCUANvK1H
Gv6BBdKFiTCqNxfW5a/iYfUdjp81eJDHtQS3OgAtWjek5t8vZYUjp9hRSkVdCsnwk+7KbMiUFmBq
/PI1Vc8vzjBXwkEDYA/b9XqymdP8kKbL4ONtS7wIsC7CzdkymKvrTfV5GvfLiUASKv5HWf0jwump
JyV0zT4uN4y0G27hoEu/iG4HbK+0pXdMXeMYwJ8q6LBL0D0H9swytDyuUv5jUQ51k86khPL69QrB
C5Arfon9ykSUeHyOzMMAQ6qyQbo2h86Jjh/BDjVuGlN+tHbi4a2Au5/y8dW4rNESrpjnesaRTiwB
QliLYMyLB/WjSfEusa3QzL/BiIYCsIEDJC0KGLO7dm4xAet2W2MJVzbPNqWQjRc50o6t2HljJ8pu
rkEFV5ul/YvQcoJy/yjUQjQ0ydJi3L4Y2UCCmOd+JXTOTpFtScbR5FGISVEKf3q9OerfsuUQyk9L
qNzabGqg/OpeVket+Ii1pScF0hMWQiMrgj9x/SCa1q0YrEHSpYkz1iyWxFraL+r8aIO8nbXPOYef
4kfVM006+FhIGbyPlTP8XN9t+mgJedz0ZC/FDL1vxtj8qtZhD1L3ASyyfxXb53HWqXNGz2Q2HYRT
yiWx5/oRuXx04FDXNUlotRZpWBCaTP+QXDeGeBXhXGT1mfmx2gKYHebSR2FjNVjM6oqYQT5x1AKc
xjWwEiKRdUqUFYQSCKSeX7f8VnKwgnMHVOtXMgdmnL84FQdQyrsck/8aXL7Y8PP4gwM9+Et40O85
IY7hr98P03Ee5erJpboirRqjON3T4OOJE9N1VqxQBTasi5r+SSDcem2rgpRKLEPXC351tBnskSOF
BTUG4Uk7dRwdONKafDzRrGOYV/atappE0WxXhfDYQoqENFCqLLOLa3esNQsQETLGb+iC0MW8Ra+t
lGeiJ+EFbHJpgn8D7wsNo2WWSBkvyQyE+91Sbq78bpRMwDENTC7nvUG2brUxanEUS8iiVMz+KcA7
USAIieNLyaGPB/5GgrHZ7Xc3PIItm52rRgcdCAQkL3lAHLb7OMFrXHII00wRswfRvu3M5YN578Ch
2T0CQYrz3UGQyn6o/LyJxhhwVFw/8idSHYKi+pWB92ryKkTIv5W902/hReq1i4T0wOsk9voc6U/M
8dHatAMDcvskwr06eWbXmBjc/8703PLxK15JGqbhNxW66ws97m3X/yXFtRVnWGKQ0OxiBXRkFGap
Xoe2ffaI5tQPXS4l77gjl6oUzb9Ichjvg05+EMirHpE4ZcXxR4DmIcJ/HZXiyI+h8/xajkNVRDNx
Bus59QKXOHJjfhK2XIqUAqJATPFgG0YyS9j6dPXxyA7iqFirkRjmGQpS5KHnZRRhAHt9fI4yO1Dd
LYlUUT/TWeorTfcSzjX4GUxujcpuvVpSCkXhmbQwbCW73jrfrHfUEbQrYRr6YzqIinvjLAXf9Nm3
529lKwUv6Z8wwMaL5uWN4++66BBJE13ICtuCGnqKS0s/mLz70HNj1oMPseZgneHLpQnWX7fTGMTn
d0Epyq0dy6rbk/4q1O6Z+H2DpeGuejeKSzXioIKzYzLvXx9tE+dsB4Ee38Yfna1vnmDOvhxXq/LV
1FC0rUby6B84GqcQiTt3pluIx1IVZl0hldQD0d7jrmqGkkJ9PWj3oVt4xYD8i0rRowIGqigFgIv7
3pRkmY8ymAYOHfbT1k0hq4ilsIyJZdL7LkTrStKjjpHMV83wW61qnZ20lQhNBtYE/93e2tkblIx3
7JYpKFrgA6zPKA+E8tSpey4JyRKmWTzSFOLtJt7VDdIh+dsj5Zy0QaK20vtyBu6YjRWbcRncSQlA
7QGYIU14akk+JHtZoaAMNFNEQ6+FcK1YAzcL0GNwbao1kTfknlkvbgyxm95f3MdDr1BpgyVnxR6s
4f6gkrdEV8ak+KXPB6l97vSQipimVZRcgISQMH7BgIqmcnArNtfgvYFnDI8ohQS7bXN7c0bHoHpE
g6F69MU0uPkoh7Nof1ghtwNcbfaN4sQmoOav6q3db5Z/YL9rjN3djl4VH2j3kk5R3laTfM6vt/d3
3RgIQr/ZdTouU47c7eZu6QkZ3eLGjJiex2LdwE0Fi7uTxlfo440g+HWgPj0wwz2L+D9x87aCGv78
Z3Qu/ZWnGnuVMG+wkX3kA7Ul3t1RQueFmsbkfG1el12Mz1UcSfljp56hISfoQWiNimBDS/2+2XZ7
ajctyw9b0cvJYgUdJz6ldqpW1t+yBz5PWOGL8uZtNEeud3AIPAy1wyE/C8Az6XziQCdqUS1G6HiN
DvD9/lv/N946aIj/7fCNI03xr5vaUaZHREzGp92F06unJXJ/SeRH+ZB+49OEnOI6vecRmlwu6eoi
neCByHfmePSQRqIWiA1xcJhMhaJS6/wYh8G2VosFI+PArDBDbq5Vt95qG2n50siRMEOkc82+jJeW
kOdqCXz1nwYliPjaZWikYYYUSX4KmhzE/diIskHDXYR4IdsCnnIGhgoP16K7c57siK5pw4+i1/Xb
CDJCYLJC+fVsWTBofdxYSm6SIQBi6KNr1fo//6vwf7dDhkGAmAJ1KATxWKTITMGMt2pxtKXpt5MF
xQu/YhJiUvuleoUyuOHOE88T9AtspSs1MSmD/DSoBROu7FChowYzR2PAh4cWBtvoqcRqjroNQRPj
BopFG0IrEjpwpRjeVyN/3fAxk7OvvmmAj7Gn5fJXlthsqqE1ULWQWc14XO60RlfUTW+OEsu2LVAX
QAXm78QWcygVkl7eYRzmOr2OxFucFNHL+BOyBhv02SGxwPZUBYhE3qJIlkfRaIaok2I3zTpXugnN
/WkJEvRhh6ZLss8hevm/aWvG3vMQLqtct5P20uvosoc+mcAiCWJMcE8tgD+AHODQTlfD95y48FI4
yv4oEvKqRpLNvZy6ATM9NMwoG5trj7CxGe7w2wKEy/p9XVkJfuCP+fDQmnPD6gU8BCHkegvjNiDz
u+g4T5uh9XzOOcP/nvlrmy7e5tUcLSUJfOEKeY6lYlWK86BNgnaovvH61mTN0yDqMM4y+O1HU4QP
/jXhyRehJ2MLRqV1Jow9K6tLgVepKhz6mjlZER7gs/Iv6BC5o55uoeahb89vEZaOHFvRQD6lHtTa
iE10heQsz2wmi4psfGVWOI3HZY9a9TJcvfFTHaBUhe3f2CXdhL9+nI6tG13lNppxJsC3xpqTtDuw
wrSlNZbi2lbGsWhO5eFZ6lATDUyU/a4cOzCNl01qvMx+Gq8LC7+Am/Hf2MqUcGOS1oYd15UN4Lze
XmlPEmsVaDrYLZLbS7rcaOruUXMjqqUgcXPg1QZjYldWTwAEDqxgPfHmeg24xxCZ2Zo2ETDKenM3
No9UtTFH2zaWmtBIewncI7YH/fJXAmN6xzFCv3KtVDmI5rG2SyhB1UKtxGpmrEMFIj3QXTRCI58E
5xKz/LmhIde5aMkz40aANDK+qkrO1VAL9lDzSprRP+ycoMqv8HSwTqjJ2be9WG2Iasc5PslQOQvG
EKDr0Eg0srL+slSrMOu51YK5zmgCiee3sd4nFsC7Nu+efFQaRNESzKu1/j2BzdYOuUwLLqXPdfn0
1CPk8U+DQV7Nqt4Mg/kqEj7Sfz96Kq2FtxIOrFWjj8aXx1hw02hfl0k9gL5VGHoAisxFaLd+jeRv
Xjj0VCvn48C9SfeVcSMKdDq4WmDuOZCnazsBHnhdevyiltNv7aFCeonk7bWtDXVUtx2i4m/yuArQ
11K+5ZKJrB2hPz4jNtIO2N1X2Yuu0USlVWLhHSxcAZa+4VMUydVYCn2NjoS+AJkoYTqgHcT7ODel
XyrpeCcuLai8E0MiNz5PGyjVallAcygSB1KRDNsfbzCdaRyMy1G/cO2/hg6deT9smc2/Cseu8pcS
MspKZhLkvYVHXk1X50qqov6bCrcSbwrwEIpkRh27RY6HDZ031NIjUySDVw1pRly6Xe2IZTmNvf3o
JwLPOTqFz4TUyLG/nnWgEPnaFNroZ3eW+NzmHr8yIE/58O5QCCk5uuJUhnhjNGz8ug/FqLQn9ViL
KtHw13j59YXD4BkbS8svd+VCTxr0Qe8qQCC3+eGrUv/WouTozFNAUd5215GA+YbYoDa6kMjUHPjD
+dotDIVJlc3O0MWAUHKI2oyFKHQp9ebaugOWLBZi4wSXGxbiN6Y/VwA0WO4CzmPUF7eE561pY/u4
mb1r262OP+4tEMpcpHDw2VgE3vRhwHGh8s1btyFi1f0qnA4o1LLEbCf5zwfjrC/7YdMPd+CIZNTV
5AOWNAI5kJzKGIopQEv0DLaN1nG4LUH3EyrdEfDigK04NGSxmCTRTDesXCwZ3UfCY+/X0i55kC+M
1zysVMpDOjl5v/qrdxYfcigRpbV9QS+dGnp574cSGWst6a2EL+WmRG8IDSv3hBWJBIT2ma/eA4vb
qYj6dxXu+02wCTmATP4DqYGy6KLRNxZ/BNbi6dESMDV+UYU8fm9laN94zSBUwqzld8xjD1nVR8Pe
hJbCwzLr+PR/rceIyR/0RO+J7ZN1QndrzEwqXpnofXVpqmCPcK4MAIgMdJxD1c26A8V2F9tnF8EB
AvPiZjlOT53u4WLUbNghHqHH4jT++Lqj6CsQRJL5EO/QZROxAXcnF2mDlP0Jnbbc/Gt2I3cOuRQL
mRVfP5WlZ90beRyi6OIOeEoZAUxTabP6wcB48+txvH1vcokFIpUN9cRn877qiMMfMxN1ydsvazMT
1ZRnLROeWX1MttbsSHFa+YjLE1pBq9DSL16WhGSo7aro2yj25HAVuD7nykZ2+Wji7ZR5EzBxbMfq
toz97JLkBfW/LMGf5yIpbeZL8OMILvYRFm7xpcfrFIS0IDbOmH3iKxf7/GcFKH8fAmo0uh0zDxfa
GCbJfwkWlFAAP85xCuQYi9IDODKjos1mSdfSvt7ShX95McJ3wyI7xN73vqi/qEMME/yApwv9CAT/
efdZAn0qeOLqb6B+swkDzRYarFjgDWy/0Au4SHAllRDdWbKL9SL58Jfeey4FsXdvmUb3IRCX/m6L
5Zx6k0RYghY9U1K/L9BvAoiDS+IO9YUI2zxojzqdmwD42NrmR1txpFdRNR86NZH05V2+zvTPlho0
/6AzCXDnr4MAB2Khtu/tpYEC/8eDvKbT4xByrOtOo85yN3pfyveNj5wHNgHABbyaQLP8YvlBZ72z
fuNDPgMbp/Ym7/ummILnbGmgVOVRQV1ijFyhHKct3NAHw0DL9deRTBSsEJWIHLzF8UpGg1Q3GEwA
4ScVELQCpTxuCkQHlcPnO8YKSw7M13QvvMleiH0d0LovLYs/Gnak8yX48rjjwVU60pK0a89XTAcC
WmShhjCbL8gUs3kBOaY3RyqnrcHUdtM5n0goo5LxcDeF+nls1jNfEuJXqRxgGrQJ2qzez5eE1hWu
4/K77OwJ1i6gSdGVDN15ur6rK+QLFL0lbs495szRIBeUratJ+oc8t+3KYenFtNWmP/PiG4oT+Mfz
dG0CKk8szgML8dCyts8Qtc89gg7kDV/RdhVhRPK/SOUewZR2LiEso0/mX6rrhis/Rx/G8IgDWRdf
i/pqEAd/6cOwfq1dv4VpJWCdrhdSChQYD+PM0mWCCFC0QlrDsOrMl0YU5QLW9k6ZuJwTr5ojT7Ss
WGCPidwfftYamHnccx9psigwTVyB8ExSNJor2UrDnqAs8cxlgXxjySxr9dmrx4Mb3ezrzVMMa4ZM
qRzqiKJ4hXpNXa4lkBnecmWrEWJzQWZLnXPiyh3BpTajMwSHVMw7dc+0v3nACqAXI/+nJM89e8N+
qf0JJsaw06MFFIxczE96dj/0l8vMJb2pZ2eH0nngGndZVtsH3TSjvVUtaifPIqGJzvPwGHWoss4y
HacNBr0B6B+kk3Br3uET7YWz5PdXDCy+Ro8Z/cXseo9RHkCezZqltRvkOkLLXSffoxgt/jw3GX9I
z49aIzeue+B66X9mI3LVYAAXEPginpNY/r1lPWCc++N8kVWgtcXoCtW2GzMD+tAAhO16Igqi+poa
XC669dwJgTxLt80UO4ja4M4PXhf38O3lzyxXS36PVvWV+9TgclilBuwSMjsKSjEr67u0sX/lD43Z
92im7QvNlGIaq0pg2wrC+VFt/fEq/x+MQi1PfhPYUFNra84dBjhzQgWDxsttDJ1JKUb0b++bhAOF
w17ZMTX0ITwXYFHDTUlH2vSShY9a5U/OaPZ0wDGQ4X97EkpVbtfZ6K1O2ZvkPunBLytjByxwCQpb
Y5YiW0B1xW3QkiX4mzbyolDCzDit6+S9X4KwBC37IQ+EQRaHvh/NglKlMUj+qpehX+9sKhoCYg9w
kjZxCQ04UYOd/0CI3ARk39E0L6J0TzsAQyondCbrAOIT3pbfWiKVrav0Yuj6QMd/khUI8+gYiGVk
BhAk1GibwMfUtcilyRmUlMjQ2uDlf0+QD5TWw1P7L3L5UE3XKyqF/Snor7wiFTj8ZGqfKyq64p/h
5VeaM2JTZ60BUyjAdjNQpoeVKcLz62bl07P06Z9Nd1FEnasq7eENwYQlBL2fg5tCawXzbhOaZKVY
8egK2NTWfs/GEV9/PLavCHZBWJ30VXVAD6uLvcq0adtBhBUqnA/FoEMKglKTG6K4LVcbnh2OgBGL
C6qBt0IIDtEQ3p6GPPQxZtlULDKhul2jHn7qCJ61LDKSdgzGUI8GB5/sWTQ2wSBmv1tvuR7WEt+V
/O8iylaZ77GSmWK/vaQdWkusU84THlOk2l6ptR7wtLhUjaMQ8N0LDomjtSpgWMU4N7izjQl+e/8x
GtdGtXltLMV0JpEQcK5KgiHPxiAbSv+cWzCGpZodQpXQSK3/jTTxm//qoNNrMWlwDwsgJ5eRMRSM
PPaAApEJT+IJqQoHUbl8EW42rRy7QdH0rbsbf2KUQuF8ArStTere6iFntAcoait8k7WLUi9RD8W4
tYo/7EXhwK4Qp4qKc188K2RH81iWWBRcCcU0UZQNub9E8TIOa2RzyVrr5ckgphT2kkUopOcowBtf
bIPceBkciyZtC0iyYso/2KK7gD2B2ZmmbEbMv2Q3s/RhacmcyILt1hOE0epBd/xq5fKbh6GKVo/T
i0ZcqlRxuAkwv3Q0/X6Pbicwom9uhUQakfByQS0bWT8+Z7taZ1QQzZq4NWxRxCJpBPIY7vvSYmqn
qY/6pWTjExG48OuUzBrY6GOP3EQ46w2p6u/yVWCwBBE72IoNFogqKYxzeUdvXA7ACAZYk5z6eWym
sClzCIHQPto/SVs+XZBBy8XmeXuFsV5ozJI/8YbJV9mOoddwR0meZgD4EefYPVCMvMr+i3+VMwdT
gZRieCtwOXmeWY1BOuPS3kEA7bshd1/5K2QPdwbUqI85EIzgYyKrqOjoDt9S0oVfTz3QRlrxrPvj
HSo2/7gU78OO5YW5KnIrb3jebdySuNvKozD26xc1FFEds5LHVJIg6jdBQeCY0EjoNGYnVeXPH/YB
oP9gkbhKpCUK679OfFFKF9/mmGh0Tr05GUq2zuL4NNcqEuQeNC4VZ685A6gb0HtuAvhsi6d6dXJW
lR/DZXVVLP3bMlyD7I36WeN+Qp5Oc+t+RKc6FF/naS46KBbHertX8qdkK7w+INJLJKIZZR1q1Vts
g5VtCnF/yt+kfqXDVZdxmy4QC5tLdQu+cOYzErNUdVJ+Ts+x0fG3jXNGr1BtXBp5d+DX0FUPpS55
qIqapReERhhAdHKkEkl3wzKdEQDPwGUWDUPOL7JFp/C799mADWaRnqoIC1mNAGez3BVhrMumFJqp
ILhgBKaKY04i1txKfXfrcEeNgbs/OMVTO3rzTpB4XPVC+J0FUkza5txtg0WMVNtpwj4+k/RKds8h
TDIQFjt6F0R3kiEao2FNMda+c7BxnFQKRwCEd8lQuDoyDyW1eWVVosYv/QmUZ4+w3YwfKnnzRBFX
vEyyliNm17HpJ3V3ZOdjcboCThyXOvQK8N+MTX7PTBsnnMhClX7bpnciEBVXK3yHMI7mL0Qaf9BY
1/6VulZ6BCzg5I0CslCmOhex4M2VVDw9ykNZldTalWnB1DM8EbB7fx/c6kgqKq+LDVcy6dqaR4F7
NYvWT2MYxhLZJgcPpbNZrZ1EiPul6/8qrSc9Cg6xCHokOFdoxHA1t1oKWe2JJMSyh5bp9Kxl5rPs
nljdaZyHFoFP5ZGwH/HFWeOxbiHT6g825+tC7Z2+Q3Xd+sVQ1IrORUacS0KNKMaNg8zoVKRvBbui
DiKkU3tvnbMRVSZiusQXaS0pHpIMZJm8VOk3gpqw/A3R2MaLHzatpLnj/WTZGTr8j5TLEh8CxbhS
eFVkcY00S2dXVIVklBj7jt4xcEvYZpr1uI/vMOvSYkwI26ZlkWpb9WRZNoMFIWmRKA2hCb8wytbS
NDjUy4yqpQdkGjz33RsNo5WxdgKxYE3kZ186SwtQnLguAmLzQLaTGQmVtwqKFyHuQs1CwVwEKqmj
Q8N9QnovFV+MPsdlO8sPowZGxsdynlzMPca1muD72FBhTmt8YCUMpSNjexMHhrjy36EKhwAJInyC
u9qrJrCo1JyNhOmzU2pI9Omt2D1VUm5q1X30Nxau214zBp21QLWTfT4L2kpF0eJ611f5JluHadwM
9tEs9POGtK3LiAwDHLiP5AF7dVrPDDf1XtvGZfLOltK6duKQOEJ3TAvYXS/73D4Sga/nX87XECuD
7f7qyfIuLqWUOIwMsyN8A7okJ4Cuw2Cps1WOXm3AoQncMqmVWRnzaVG3k/WkSLdFJslsXNmgtZhp
CDa6bKlnZkLYcL3PIoWmfyUGOE1O/IoXUEAv2Px3s4jbulcJDY3A0HMvcV9QP6WGUk3ceAsdYzuy
dFOI05naPByrgk5cZCxBMEETpkenwj8hx63cxtwymGjoLmrOfv4CsyJsyzokPg1PU5L99j1gjro9
3JVqUC2Y3vHdToPSBULA71rQcuDkveAyvUWqiqQR/AgSAgmUyUKYqRQvIIedeOXc/n/fytcU68Rr
GOECWA+FMUmzU/J8NJ7mNXIRgqAj5ojPhNaH89a9EIgU6k4P74wLijOFeqJwxHPIXWfGK//k3ire
eqW39Wn98GQ8607rVZUIaUlMzqQIm0woC0cgosSjHG5Djlokl472/1HPUc1C/+xmaDGRs/A5Dl4T
8iuWtcoik1jjdd3OlG/CBklxq0aktn4ZrR96VAMmXMf4u8oUEvPgeeMhDNNOqbETswWcTSHoUhDu
68hWnfBgPzczuzsv0Vioh/V5HKEtRoz41UGTA/QAAEWhvRrsNIvK9R+OXLLh5qYz2MeyHzohbwV5
tgz/THEPhT3DX/URxHStSBaygH/ZNpcrsjYSUsjXliFRO/BvZNEf1Sj71SkCa+QER3J4y1zpTG+N
BqCnQkyBVA+5miXCVdwBJD4WKqoSJ6SWMV0q2duedwlDhiyBfX8NPNY/K3beEbmwbtyFa3ei5PGu
1QUp0Sx3z05qMTjAdDzL989ytoJrgXrjHoFZ5GF+TlVf1OJFSKQdODb59whVtUz/kb/cgDthbHz3
qJI4kzYMhbsShiU2mcRnZD3g9IMfFKYBnJMTMfbNLAmBjm7GfOwbW/0Cw9Sl0W/PN1bZQY4P8TDf
dBBOI+z/wEk6P1Hfpk2pXy3vmvE8KBdxVhSig8ZvqSgfG2q0swbCR+9nx349R2dv2UBqHRxq1fwT
3J3IrW3O28QNkIMOzicpOs57cJkTB2c3sQRJ++ib6FWYU2CqsjU5blxZevuRZ1chahSOt/EuPUEB
k+ijtqOAK0Gw/7g2ZPN+9l8bgSadQE33z8x2VpDdxhSKAWOk0FWhLxvEEnIc5tcVckXLiq3byViB
4ymX0+WkYKNaOAbuaH05MoPqBPmivB8yoolaFO1TyOgHkKDCsiTRzMSPnSIfK1Xci5n1JKLWWwpO
1QuC9+WKS1TKp/frIANfzQhPMywi53YjlEhaOGldcFUBQ4yhF0RNUSY5xgbqfWfEMHnnYgBYsDP0
VM/9RYvymJzabBo8OJ3Jp45PHKRbzipIgPNSwT+6A4A7/TT6yrTrAGpAX12YCXczQC2r7WivDbTB
KzHC3KjjTUzW4BQwsp4AZtTv3La86bECNiNXPtJQsDlLQTmtNcigbzBAQlDMvwP9m/s+8TUFT3Gx
gmrXpY+IvyXjNd5keaKBm9EZT8tLxYqs90a+REN7wn1cwJfAkE9R6HKqNMaEjAwFoU9vWAbYcvOr
fNLGxFbnjxRJw5tsHVr6eoTWgjt7zjpYKGEGkbZiHZ3ZcrxHgzc2Zxf9URDMt1SFYw06Ua5XGmWM
b50yYN7yhg/tKXQBc66nuRfw/WJIGzv9CNfvIh5qpc/R6eRSTPJBLQp36KUxHOnIeXHVfsu+6V5N
e130FJHylsfRqfW/SyTz8WwCN1jMG7LeBubEPcH8gtAerKa3JnCsEi5fCcHOmTp0bs+068wwqPCk
Ls058xaAwBK2inX0p6f8DqRvRJV3hT2Nxo5Qy1RJzNN5VfgWAnZ/kYym8W4uvnQcz9NXFuIPHicc
ExVt/U9Vapb2k1HZBX2v+vjkmNdoyOuLu2GKZGTqv6m1g1wxgNCk1geY8H4GtHDrXYk7zVr1W1WV
YSuh9ZILlWRKtwF5ISrfcrSZ3h6CoFdnJG5QRH5tYZcTJ3ljyuw0pY+vXyEgPpmABMuAqH+eUtHs
RQHA+ugdGR8IVc1JkFaZaW+/3EHxIhVXRmXo+wfSRqdwRX2hOIHmOYBb3PPvlKfNwVl1lZmPnZ6U
KSyxIWIOHM5RGvyoVdTxncqYq8E5NPSEoaB498tVjiLQJVTgIKv0aDRtNxRG5kSSDCqgdTueh6EC
8sV2tK2FdElDFog7B/y+ZLCl7186xsHQ+6hhDLxNjp9mSpHjOrzg169AxoExdZTBgM2IYcV6/v7E
hSQeuabUQt8e4lRnDnhLoG8QdOknmVA3HYUL2sJwQoch6BvORKT9rE8fMS/HzLPNacMfmcr3+zBL
2p3GeDknDrfHNQpJC1g3lRddl0pJT+v6mUSqZisgeury7wEU9xLEjPXmG6F/XpMVCX1DgfZfPyGk
MFJ7mtNvKcUgjWMkadiVfqcmHtSgHoHo1Z4APtFiSSJ4Ly9PxPQtpZgAIzHK2+c1H/ocAj9VE6RC
FLImutS6ZYOlHhNJaGXXFppw0bNb7NNJFVqgykJmiY9mKMHddIrCXrnBUFCdKKQZX1m5tO3vYqCp
+IrmiRU1Jn/db+NJQYnROVHoSaF27CMn74WcnW6O+9JHG+kF+TZ2LG4qziR+jvNVKxLkmAbkZ+mA
fvFTNJa2i34GLUDW0WZH8YK0hXZV9+DBBTFje+Xoh7STzEmiCBVmRtZauq3Th+LoN9yy8e/cYoxV
nFxYi3fR84VC0bcUCw/izqWQITC8Vrg8+AUjaGEx10GfSCPsNIVp4eo8DThvUbaYFWiUNruouIR+
UKXst4PFO3vbOv2EujflSwh1h9ughDXLxxOY8jOGn6pVDBovoH244YIui2iGmrTYAa8isW1yTDiA
yoQQRqU8uUe6ATUGUagPRu/Lb34WGH+9g3kp3ZwCDRlVSSTkXQaK1p/P5P0EUHBlyetSfLzHQWMn
bx9XBaCLH5ZRT+BiusLbRAMPmwwX8QqwKS7i/sine62UQMPPuQGvaeoh9CKtP5Xl5VrLncDGvYrp
VTkPu3YQiFdJ9z1ZhaZON1IsEQAgdLLI37jPgYErAtB4rbyCBD1Oue80MtZ7qeRk9RR2hXx0eqOH
wLbWKT3xpe9iuPeU1mtEgP2YKQN14YCKY7LVd6I9pBaJlUy1GvJl8JiuHL8QEumC/NI9b/yUnTcI
bunIORQlD8iYSq8XdZotaUhO3chX/GSD1l3cKlLOB1s4EaPtu4vYHzGkA3EJlURp7RKGx5E4JtoN
Eky1iiQZY9dtTf/Dx/VrT33AHScbq7m5AToc9IDqHAbXEud06iCxo12ycfu0qPZ8fE/hWUZZ2M7e
Dz6vJsKWqcAzh2nBR+wIpj3AU6u41rGTMOuAhncnyPcFO2PsKp0ElJmKfn/UWpINPyW9xVFSTScm
WeF8urUFnzTUZjGEmnuPZAjsbM8sANDgrEwpZAvVBrhTA1Sfi7WVqlYFPWVWrAG2VENA4GZ1HXdu
HXNqLplrE9cKVvvqhHBk2ZRfp5fDc5yiSBf51lvI0fEmoWm7luPqZpujBTsWMwHDPUD9owB8Tr/n
YrbbfFvMRy8IFOH6Ptblq/iQUuMtL0ydrdjIe3qRfzZtuFXtV9ljwr+fc9LZzXjgolxZPANRZh2/
on/BO5Vh3eyBHQE2jumavybddE8MGl/UeLD0O35qql5DGv0s0tXfJaQ1GmfeorWBqgExxl5mhX33
9sCgqTbOAIBbOKTySIH/wD4uHp+xFdFTQydVBwRD1EDSG2r9GFEh8QB6LeDdrRu9ZNX+3/u1DCIM
2pnq+GzjOIGY9Bp4sXKlCXhoIJscG/KQz6qdKpSd+BR6kE3pUYtd2LynW+ZRJmNwdX6l+1PfXOv+
qo6SKnERADr9TQ2wr/35vyJaIiCgYz+G3p6PSlNpcQiqeXSLuht9PFmp7syKsqFQqC9DMq20dxMD
PKsYiAkOTvSA8o+XcTi1BfxLXeOlc69xw/6Rt0ETtQUh+3p1eyyRF5ByeVTFZ2W6GDfIhflBc2tg
Ipk9IwVDqMQbFl0w6QhbjeiXHP4PqArUsiZBglKZkP54mVZ5Ak+uiG2bBgYlZ3keItooZUFhXO/M
p1lvCW5SYFVT/bTOgJfFTFNQmZXq9KgQzFXlcnMpaO3vEFR2hOmi1NsAYQgcvtqy5oIqJi0qZoFq
P8u2sprnVIj3ySHseMO7ZuL0VCtW527oa+10buxVbbVmAhlSMRudsiW12sKUMdbp9+urFh3ZOs4H
Yu7HxWm5Tnyqko3coNcMgNbq/nE5YKXGEc+M6pBcq3NKtF+ehySCwiTGlifSkaExr2xeMrvEmMt7
v6r9e788OET8gBWAtNNaEaG/w2zISOQNAiIPJDJAkganRx75YalUuOLPmgfSRuvNZjyO1ekQJbEN
SB8TysFTY4hCKgtZnb6FhU45x+H12neQt6LCNT7sNZgTMLbEONKsTXBu0NQ0lrXesNTCVIQ7BQT7
bYgsoYx04FhC2vxsQ4/2vNJxJ96naYL1Wrdp0W/AiQX8Tmd0aWy/Vv+POnFJyYhIajGraS0wqqqF
ejThHnAawsh8wTyjp51/+9gCvtRHOB+2l2XJGznMbQkR6So8Umb3AaSH0uKC51IBgbrSnzwPxNE6
Of1zHJ6Ei7MRusH08mXPk2oC+ADWPsCcXtJ0Vk5hYo4XmVfcBnb6lW02T/af/Iy3DAaLK7oInSNA
gQNtTB8GKb199Z3isY00U4DPpTxUthlKkGLbo3uq5F5cALFkFqwgzMNMTujf4F3MZ/5Tfm3p1BAG
YGo0xpyFvqMDEE5cU1ujAFBiSnQJ08HMU0T9BHHWS+36LaawDDgut4OXx1Od7LSsFREuBgXDGgfm
kHP9ssJ5Sy8BVrUfSxqHEBN5yWSMb7TC+tj8t36815haS8RUJoNFXnFb+UcEj2AoyL3drLU3Q2Lc
fdKHnqyv1N1wINHUGl7l+diJz6O9lkBUIRCWKR2Q9TiK1fUxEkWbLh6qz2q9kiFv6GfLyRQzRiGQ
j7R70ZRihK/O5XXLkFEIqEeLwhnEJDJGrkVXzzgnNbIydiuojzH73GTW4p/vV5uJW12wF7Mb+rIT
HeQzwVFH5r0knNOaqujIRAJ67eyfsRnvGtQ3E42PsmQ8zjItg+AEegNpy2jGuB1AK4bFWecrw3AQ
9FgICuA6Ke/GIirEwHdzIAcWOW2Vybr8L2XI7yELlp56ZES4KYAPGjhLSh6y+maWc1W31VCIKDTr
FHDF5mlpuwt+gNBhsv8xiiSbu8zKIuPflj1OskzWPs0rRQpqS1aXyFqyu/xnk7He/dmay6iCs71v
iKH6MHbbVHIBS4DL6tEtIjDNhHBlhgjYQbMYGxmuL4FWSDRLcR8gRCIq2StCq5ka7TGUQNPtx42z
QR5EdK3EXjPYA9+GEP9C+O1ddLdG70G7EfB7sz7zA13v3qzecYC3IgqDW5oTh962POQpGoSnGMHN
fSm2N1QVR27HrsRblHGBTPw7mQCubxjxsXSgWU+oDUK+nb8ei6wkndOCXW0SWrztKuluAy33Q5Iu
YpGf9wn0R/DQd6hCPBP7HPS4KgP2+ofC1TT8uypMWylKlDhhPxBfyI7v9RBUUHTpeE2QfhM9j/w/
R93vNmWie+P+hogvCMVuh2nnakVyfpVVeTEBYFJZf/iFSGy6pgRBzLAxbpWNuNq/drXYpqIwgvxu
1VP1FtOsEJZUxBGE4RDT9HuW21s/Plvy0AqBfwxx8B7P84/eirsWyPKu6XN8G6OWAlz4GNk/yT45
dRx4vDH+mpaABbRiGecCgQHle1eKMxVKpXYBWeBGkcXYDoyjUWKGKCDH40pny6Nl4U9qRatJ7/Rl
+o7buKqXsBRw8N+nprkj3yZQKeB0jBmvfRw0TSMeBizAaxniq9GkMED23/WnBZjcCFVav5iIg52S
IQCbNA+4iPdOLALHqpw2T473lf0OkuBRW2YK3SMi0Hz6ASbUy/nBq+G3N83lABWf0G01J4mXk0g0
nxymAQmdnSJ+V/zcePNlF3uGeauVMXmdsz9+uS+9kPurJNEs3U6pgfY5AF4XzHr/M5w9xXGS/aCr
LvxWyt0BsSkXRaRGjAH+nTjLs4c26gTRj64VyLLR7WuLWHQDxdHrDh7O/LzU6mQbKPlF2YJ7cu9i
d80GChHELnQ5rDdxL/vUDneIneilQT+YrGweJeRfnAKT6zkaAQCQFgwo/NdCH1C7cWC8+HtgkboU
P7d1d7JaIe+iIgnb7mldRpzFmLjL3haRlOELHt+UTPdYkiCiN7A0sb3gQ+Cd8CmSTVQk5bfh5wvW
KJlDHIAZ+wx4/uoiEFsAgiVDUctjWq9Z+J4De+T/JzHVb8j0hw+B6HzTenF6zH+Z8iHWMh6gDrEe
uhuBt0FF+MNR/WbLIqTtPJ5M3RzWYY7oFZsEXiV0nexP47eD5CKtty90jmbm1WPko0jIqux6V116
FXZNnxMpP69xRYbs+zsuRMWjqA5oP6MOIPllHZcOvSLJP4XrlGdmmv7rwVdadZwx5lF1wVaaPqfB
JQ1SdyY57PACHJBOlc1Ke+hbgrDUZgbC3gVGwyFQKTGZDOv3mlm9ut572Dv9gkG59BEa7hU8bkta
oy90GxmR4DwvEcELGJ0viK/9MGbuVhHsUG/1b6JWGsTOdRQ7CVHIKfJqQ84CYjR6ZY0QZkBxsXiW
TGHhLHL5YEJ4po/V3Y8rk9oeYy9nIH2IEt0MT7kGQ2rkpxvSt6/p6Z/SUis48ZxbswIUiIE74PlE
2H9XzFDzXl2+In2uJdbU3ShXYHaNW/qmvkCY5b90OF7ghyHPU7j/sUeqYko6TGjPKymZSd/gDHPJ
CJqZkUDEAi/EaenUWQopse6hC62bJoyGgXeGDgP5XCNNVo5EXgGV3Nk4DnTbKEo3sD5BxaSvZ6sm
9/oWPnBWaPXntWy5hjNxJRPxRr/t5EXZ/Xv7IbWgTUmo5Dga3gYeWcrSeHncdku2du05/dTtYXTZ
R+VtJvdlDRCZexPhgZPIszEKY2WCB2QRuqmq4+ST9i7bs5yDX6iDPk+WX7El378h8qSV3VuuwPYd
+sJwPGFdTbVAA/3SREai7HODy8TEDZzyHiLnloaJVcv4HHRjaMPsoNyb7Fr5d+bLEihl8iMFdqrF
cxoetzsURIRidloydX1tlT6IARA4+kJQx8nRen/rrvh3/ke7AWlEHb2MR5BSKdGpOEFkHEMMVwgN
HqcxSNANZ1fmyN8gBwFRXoUC4oM7/LVF8V3Cub50jhkO/TWR+EHJPBjxkg1DxfxTn2nua2N8K/dK
sIOvMWu5Ak1FQqn93haabvv+72wXBe9xmKSSxOzJbgAlZ7kad3N/qDE6Xo2yYE3mrSSjVu3sL+CM
5CVsoSRv/wtxdWJoD9C/6sHoKC3OOXcG31gfMGencN75vzNSW4Qsimd+wnCW1Gcsa7oLA/zE6kfN
4sqAc1QYeDbv2MRojyKyVpF8foM1A/erOn9sfXiQzbOxWrRVeh+TXK0ZvK44HhNVBNWjFpYfsXqo
nx3XZaS7JlxIDGVngg1kdQ/wn8f6aAwJT8e7zxmPp3sqQ3YcMh+oz9wlafcbSlyoYiDZDYqxl91X
oYm+C+krszx1GKqekUGIgkdlLiZCwGL5tudiubbFb0gXH0MLAypiDFMxCzVKQ7SZjkTR430tdj8p
9IvG6lXweCBVDh7/7pwYoCepfQLFMs763Er5q1gtzIKEC1s+nUk91ldpILIOXZvyIclA2R3AJk15
bq1N81VxCmdwgVjaAhSBhIqAJm2wBcyRr45M0gd0NLEUUUK0LXNZD7sdI8m1v+GyPibR2sIDKSqJ
AyYZyg7rlRipPawG0x1H6N1Si7CR88U6smSazhmLC+ixF/FTVRD50iN1LYfCdwvUCKkh3H0I5W4n
/x+59bJVIg9D6YhGxAhliGbquF7jJC4vC+3FR5ebPX21/bAsg4Q0Sv3u0QlHvIE70A/F5I+1oHwW
U8QjBKuiVaDlieVBFDJ+IQnbCsMY7p1208O9HYIrp+q5SaKyqEUCI2j9FmMyx4XwMhUshVyu9+u+
ph9UJiq46Y5lp0c1pPpIWDqb4UVlwqmBiy7/BjJRNKMc4GDCjyPQap2tzNW+PZKkVRwvRf5L/gHb
loIYbWoyHyLgiTqQ/XpgK6Sg6347BtSmdYPE4ZLjBkeFQC/68wqKuTdupHh5jMOJ3EDONmLBCLyb
cbTXfkzaEt86SfUrPto4YIyHd6obdBO0/ovaueOVOaxWMZc9JQ51roN0soUABxP23WvSClJitrdF
w+Mb7l1GaHlq2nLtThZf4q5ephegThW4+uE83qbK4hGCl7SMtH++0QUI6+oNpge+cpRGZMDarxJw
1otXPZSHwCwCVe6AP3UkAVHOADc1o0LRPBgTiFud2wERpQRcjp1AdhgfMW0dNkGcuBHBq7//qNRi
Jh8+bMda9VnvPwZ+4Q/viyiXqATCxMO69xHCrLeDEpG9RnLVTjw2zQpsuJJqMfZ0pNb5/G3mdfpJ
VwTbozNJKuuLYBTym5HflmxP22sm2EKL1wICz2t105ZELFTF6a9MO8MhVQh55M4SQxvqeGAK300T
0AtVFmk601aduQqMFoaIlOcrOkKFFGddScXD3QroS1CQnKvicpVuSEqTQtgWm5wHa3ylW8bJ08bE
KwqPqVZDK4vGu3VcPzzFNzHL3Qz29xTHMqSHWfcudCjVV+xVvivNKysHNBpZf3Abm2lqyuXP/4mq
GRo0ZQ3HQNVFZiNO5c8ank7Di/D6S7pxfKwwuJRIRrxcWbL94JnoEZA8kKZfoVfFNFJBcWtQOY8h
nKtNBIvhoT4EjlsDTAor8uiJqVG2MAjc6WFzHmXUn8LZ0HVikaay8yiyHPqJy1zn8RRHJ9OA5V8z
Rqlp9vLVAxYd9lXLm7b9R7u+pqBB4lXXi3rubE4SjpKlNCT2Z9u82oshRDDvQ855soIgqY78gJxh
0YAyN/Kwq7/L3FMhUlA9fLHBbVSKGeXF3whwzSos72MAnFUvhnJjK5ILVPXHEUSJzW18aJfiFKft
m7gvvCoDWR/Ln3e+4H2aZHmJSD+KlvwOMp0LzqjdpZZBJlLWDiNjPUveeoVuGewyO6dXXgB+FfUI
aKGkx4+0jsZuzJqs+G8BYH7gmZNlJC3al1qpGvUc6dfaYR5ZzKvK/wtqnwjq4rtfCrOBA7LqiN62
0Zxs/KYJdlDSvMFlzvAFQunn+t4lT1Nz/7BPSbcZ8B0TmT6Phjx9RAP9OBzHgGXpIFsNqSQHZC07
nLTYJeP1xm0N+56X5WjXMVzgjKkCkzTSZUBq0mbByhupKc6ALKY6foeRG0PfWP5xp6zpTuRnoaY3
fT8YnY5PjHqsjvOywVm9nrgayiOfKw1xSURWibgEe6zBU8QXogy+tfkO4NHWNVomVOs+A9nqqIki
z6gI/aG74ZtFHuVB+351JtVAOM35ROAZaAQuIuSHXyRW3YwqgI/dFAlarKcdeoD6ZpWZK/czu9Sg
vdLn+M2a/4D+quBhpQvDvuSLnCgSjVl0zlVkpyJsFVAkWMfTBZHVOGfgjpuaDYlG8Rf0UFMw8us1
6y9MzloglrkKdWDJFjlOfZgogHoS5jk3LnLqMx3oihG2VfcgWxoxQJTEKud+N8tfJqMU29cHxqXS
8QlFKNnQ9WSRUeomoqVw8cRtpVrQDwPl7nOBETEw4qz5zC/yOTzoC3YP7GFpsndh9+sLBZMjb1VV
qqlncuhSp121tXvk9n7K4EwJUQ66ZHN4rgzvIBAGVYjG0CKIGUMgC7m0zYWjcrhc9pLg7CPzPz7F
+shEE5svimPSAcvjhYXostVuKW42uS5PKqkoCyFnlQaOd0La59j5Wfif/KUxR5RXZ34gr6wyTvxq
qt4/caHkHrPk2hEwvpnnPij1me3M7u6Dsp/xcD/24DgjnnOx2FxiTQXru/skhc6HwFfp5NPoUDD2
mCRrc9AkvnxalbySJV9oGJmP/fP37/3DfJNojPAKdoXtOWAinyFc+iTdAo3AvTVjAuGrECkcuay0
+UKQhliL6o0lsoUka216YWRup0li4gll/Iz0yCF8zof9a9Sg+1v6y+QKcED7RbQ+8P4hw0FtFsw9
tMY5FSsd6fh/UkjlhFqmkJYqlbkxs2+T6Mis9Y28RSrQPSrkkxmewHPjsMDpz+CLB0KAn9LG4Lx1
NiJTf8JrNwUVo2tlzvj+QSS1fM1EowkFfva+krV/HC52F+sKXpJPZGpOx0R7XMeKf8c3Mp4xMdP4
wh0PODkg6OKtqCfGi40yIapi2zfvFKrjlJldOwFis6Z8JdCM+kqhD39SkEHELTwUIX9FAU06Me0r
RZM+qw2oyr65jj+b/oT8S+1Gi/RCU2lkGMPKgMFUoxEsHKUZaa/4E+Qm6tNPFaRjTb8wFS/PJjI9
DJEDZYfdLGf4I7p9lvz8rwFzh9NaM937q/TM8INUeYPUkVOe1lmiV6R+6B7b3JgFCtIY3fFB6eDZ
S20WN5AGGjSindfYwNhCmdvRS9iAgYEpw4m51jjZMqOrBDUj0znc53Xyb6r10e9sS2I3vHg7rEvW
c+Zi0I1G2kaN7bFd6DtqM9ejwJiG9krDCPgYvp3d9OFIV4S73pMqANzaKC1uaX+tg/5QS2vfxsk1
n0KaFewVx5Cd55tp2yk7XvffqNbWUHY4X1ruo/zlBGojAC/nkTx8CV5IV8EDbYEoFmwhJnemPb9e
PyReq1q13YjBkAgXaZ2iMh1ChYZMtaIvWlXT4BauQ0DVTuvb1A186vaYgCm4cwfxjHb8gI17k3uJ
vzdQiaDdxfTkxoiaVRbWvg+hUCX3jXKPIH8Fms9Pg8pOqz624JnxOxfUWaO3WPlbs/7jt14VSNwF
gekRqCcRJCneXcxKpaZNehe/HskU21WJgBYTl17JxfSRO7dBR5XqSpLLTji3ubAwasK47PyVSVma
CD1xfj09eF+l+AfDKSkN06Rc2zCW6ji1JUO8RnLmiuA0xNFt8jrFvmNfwWydj5gCl/f4YJwaAiCW
ggIsBQT7GDFXopxVf0a2n3sHi0SWD6+hVfKidSl4FWXFLv1W0GSFTw4/EUTUkN+k6iULyIXovG9n
4uLnSw6IXlWCRzZuISPjAoDFATIr3hNYcRW3ADn4skRi+07lg3bAnTswV8HT4sQLE2mrFwKSABnn
n3eFidz+/sEOzrGr3VcCO92tiri2Gg7oeYTDlsa6pum88Q7bkAvRKZ9Lz63EE2FnedwdmJLpmLoP
/7AJMCVuxi+UHfkF6s2TJ5I4KmHcmQcHjSZM63+WkzpAbxWZDCTm3rP0nZj1IIKIUcFxsVT/SK26
LOg7yAi54O2Fu6czeU5ukORm+BJql6DSZ5iQTZRWnMM/gu0gB4/7yqUifFcSkBr8HK/PRII3WpLS
7zjqhYlUA0ioSeNy3RTXKRdH/xMc3yHGl8sUAPihnM7vPlw9bYcuUsHD2+x1Kp41EEYI0H61TDIv
M9g4jO0jm4gvq/Q5eJjPVDV2u0dw93SPKUyS5vGQEUTFU5FcI8YRZzWSeYgHAZ8rR1ob6aAbQ6a+
vucxU+dkROvsJ86+Dy229e5ZUV5RE09C4duoggbQKDFxU1PzA+Hcazhww/VK0//yghTRYvY5aUwt
4Gcl+6Ta3wHaO4Ji2t/SZ9tDzBr1JeU1cpFgBGvoUIE8J9G/ZfPCUVvBOgw1YHlJ3jnVRvNbtoRI
jTN5OrUJruL5Jz1CjxCc2HNPtz1TSToVCkUNFXrbTCY25MQ6r3OZ8wLQl/vRNCnOhT2u3rMDCPzY
4vjwxweA+xqhd0XubLZGaz/k+pO5enYSCM+MbVvucR7sunBzhzUxAkF59XI7yRuLbk4xQuSYz3xs
wMDoSPyNluJ99S2YpDj44KeebG4GS0eaZbeA395soQJ9v/MpMTqndbx6GXgdBt8L8uuctnxHz9ot
AQ9UrhSYnoy9hxGT/ZMvntMRiZGFDcw4U0mVfwgJoSxOkPPdkhpKyyiHylcWGA9lrScqB3B7iaO7
dDBMrNcEQcW9o2ZUvXsmOLva3vvugjuLgJ04I/K8d+wnwOmHMmSyBScUwrqiXuAHVEAXFKwVDu8Q
Dse7/1kCyNYqcaBS+XUzbYvBe/C7p6C49Ox4Mpr4tTppVVWSn/MjpMNEr0M+8dKilM6bRSyKhyKg
IO4WCZirghjP7+1JRIhy0uQuwk78XJysrLv+g6VmpTm9ZXJADfXVYImnq41nhqOQr5lY1AwfcyKK
nbFeI9A1UNne1K+lk0Df47lzfdLS+7SDwqMopOs7fAHwlUKajJkaelWSwRLdVQwwEIhhYszoqiLB
1WWpyQ5YJUHQDfd7KHpCnzqIeT3zmuRuET568uZB4O94rYQXcB+RS0F6O5/FaF9Gs45qLGbento8
HPjyPukNwHvN+mjpmsq7EZZMrvpSZMFP01I9Ejk5xeDGAB9wKfvgu9uz1w7XKeHTshExpPrRK3s+
Ng3E1vcZbP69Z9M+L7KVzpA5R17p+lX+6CutQjwIo1NxXxR9G/6mmV9Q1cHCv5NI8YbZG5VY5t/A
EeiUfqnqnJoTpdeMPPyThs6GKx7ynDVzBVYodLwIHrgqFmY4U6V8KxmvJPncvuPgyQUwd4d/VM+b
Epm9SN0LnyOeOLsXK9bIvMN8MosCSdjkFznbARao/rEkU+CUfqhikfyD5PsJdYvGjjCitvp2+AfR
Sq+vMIDIwnlvpTRYCQkyCHW8ydZ55onHkRLniSSsgWEvdJtec7H8NjNlHG7Q9Ew7/yPFAWaDnjbC
5IQt9IwoKYeNT43+r/WCrAtIpQoBRx3Qa2+daUKh7NGw880Z8IdW3qKxTrl23gMSuc0UZBM/TzG6
h4MhSm4xwJxEE7yjUxTEvuddQFIIgG2S6RyLoigWvW5Yp2HrIBJERCzRxQ/z5s4W3zdbCVAJWLXO
m+0gSnCBhCpacfCHOMDmI4PKC+xrvrc33KIYGcK0NP4lO0xPyu1s+s59UYiZi+VQY6SYJ4a9R2l4
6ae0dToqTUawv2A5aXAYp0t/xJQoWflbJA8G8r/+SLKJeidENNOnyb00RoBSxN/cGijaALUnvHIg
FImTOc2v4mFvN5s1+h8AC0S/r4iXR3kOLdU6LfL6pwP/sbdYd3uHBnUyY2CX+yrwNSOaseG3pBoQ
bepBDUkOc1PHq7CyGchbI5Vv6H77ail3YzIg/NI3hdSC/VvtMgCdL/R48MqEBPcNTCY3W6GypWc3
/RjdfJiYr0+t1lFymz4yZ0LPFUFox1ri1KIPJKnzfaKMTx7nJgPEDI/fm9/4PGGwiadEOpLiO0SL
UqBBvjxvFHgLrutcqOvFQeTqNsjTUwHf+706KZZ/HmSJ0OlC2nVqKKFVjFtKRcekr9zG2RftLucX
tdmA2G3ELXeFJ1u/cKcXNMlxd2PIcvl5KFuwiatJu1v8OIHaTxkZwboB8XKZfgxl9cy3iaMk3mUo
IKnjD8Tl33SAc6aV0vVBzg/pOBqiq4XtMlPZdSubQVtJrKGtwIKt/LvSH9OLgO2fuIv7UecfeyUS
cC4mjy8EY2VZUqdN35gbsvQVy54GJZUxLUvOdlcZcUi4INHf39XjxxDTwVz/zgbZbDJ0v+7w94Jf
M+BPfnXjXutHrGzMhN4lNm6bQ98tGN6NwgY5XLPCcfRv3h5yv83mYCKIQhYRPOnlVhL+WS7cz9PH
G/dlzeWv7E74dtdhVfWgTgv29MqNnLkHsJ6GFT575tNHlnaDStn0tmSe+bDoc9lpwRSDrQfKsL/u
r5MRmA1nTI9tgTg1hkm4PzrHACES0GwVq103y6dsaIACTG22imLIbdLA7iszC+52XS1cu99uSzj+
BaTbppRqo86OEjadYq/TBLipqGAwC2BTRmXm0h6buxee0IkONnDoQJFI72dIWCg9BzcYLZDdNprm
DI+7FmeKYmp4wmrm2m76W7lxGzPwJSuyFlXdFlbKknNtb/gJ6TkVQH+pocbWLnQFBo7cOEVpdtty
CoFMa6unROqwGcTbFGWas3HUPY7g/GKtdNrj4HLhCaCDcXuwOWy6wuXu1wUOgX8hD6luUbbFNBQL
L7iJXfacgXGYLs0m6dRVgBB7dbkf0B2gwZDH9svTe7auQbTjZJrJINxTi1LUUEoz+6Dw/xnoZkGa
LVFV4uHWj0JLjLjqrQMZWV81NrkUj7UXVRswziCPSrljRLwiydFGips6hJ5O1twneVPszrgqWyQd
LsLIZpULZFXq2h7wkTN3tqRRC5l0nE/8MTvC3X9X0qFE1IZAOldQljhcPVIvVXf3oO4fo6sBKVDJ
u59Ow5Eh1DSwwrUpoybK+877vPIVL4q1ctGtIxkbBcTtEp2w8tu02rIheU8eL3ABD68PgsMaDpKE
wQv3V3b6NcLJD9lfySUciwGpjhX4+tEhbmDjnZDQStVKsmJzmre10mhhUwmwb4CBWUNZqhARupNa
bRloRn4n1a98VjMOewIm/Q16tkuGnZiBbXAD1zJfnY34J/wuZg5wBBYupbdDK3c3fmQEzm0eOIcG
/rp39GBxT+zyeVgefzOhlgDHvl6yyhV6QLShLeqhFFHKK8U3N6S8+xRt/9COZPqYwT2E9WNUY/Vh
t0/K96EyEzQW3Ai2fA2/gi3Ij0N5uy3/io7rTioEM0ybIFPagYCMeKoSK4yo8caNokJ0XO5OQCFg
4+Z0KfDt0jKDYUmui7t/6xI7OCpcF9ipHGE78lA3ioPJFvPwsis+b7qXj/KD9AdrUYsHYxf+hVg6
ed+UAAFeWQVYP7NrOTR9zEA8BaOXcUftHPuKQfgXa/hwCUTp+7DAOCPl/kZlnb+LLTskbjA31L00
ljpnY7fCYzAhOBkvQ/DxenlNtFZUXoHvWgW1nLxErd0NTjKbp+PCAsvQ/oou/1/M5xLt6pD7Bzhw
fii4uo1nYUwcRYALgH4uDj237jVV6OSPpsiSlsCMMDM5KcTbPZZjmiI8DNPxwuNiEhMhmv9PFg9p
yeMItJTbl9ioQFZZ7VPvOYyALyHEO98xb1eB/qL+CBjdaZ3G9Ygw0XQFcxG03JMP3lnHVKDD4HRy
bHMpDD3hnSauOmfYnx2YJQXin/6bXRmq+dlrDHNkDnPA+HqNu2+lQSQhEkCcIS3mvw9rQ1aG01vE
nRTvF4sngtNZaAP7oaK0+6+rbv5/fwGoVoFltDNHrQmUnapHc/kyI+Jr6o13OHhlALXlb2TvD4Ht
Di2P3uDy5jg1romMb/rJmxtoQt70MP+GKsvlpE8B5hPhqt4PoARe2AlVyYoBmTzAbQMxwAkywHkQ
JcfMGVA/1vebpdqff0MQff02NF7OUTxtuSy+/VGzSIEHL9ByzXaI8WslesMAAVIEuc/eFYY0feJU
KMa4iO/Sr62/N1dPoDoc1fRCBT2t0X9Ygoi8CNnFv5bpgh2a02H6edFPdJJN3S/SytSJv/Bkiaic
p76LE+KH7f3itP96FODP+jnhuDfpEGw6bPk+lTuZXR8cCaZN1C3eS1uFQsyztHErFPsYBr4AyeJV
dYR+5sVDwr0FTWQbYH6LCIPjlFQUVMxplXeRxEFGtd1nbg6z6lq+KVz9oXy3+rRJOn5Wa18a1pOH
SkTLcadkAdojaMjgz+JVRi8VnHKPTDze0sj9EXRfKBSiDJZxJ8rTEoH+iB0O9ia5538swkwWPOFp
i0spLyfj8KTSVOt7y4lN/Y80VhHzO1/wvjkxwSsWN0IgIlKTCelHEU7eCVokIo0nfFnaQlkGMOx7
FqP1zw/Mt1Jteh4aeb5qCvTkxtE3HyzduyCvkSr0PUIw4GbpsVy+rnNHpYTLfoRDHWxuAs7OmqXH
F9q06Petq39EznxCw5p8CJb+n2UeFsVW/h55KGEW78/NmI9GuhFqFNU5o2DL3jlxhfDR/KdqIMpc
IP4wCpQRNeOn+dUhR7YakptUaqOY4srJ84ruA4sgfkmBbDOXBJyFdwVSh0Rm1jlW/+MvimaNGDvJ
AIIejiEoT2Wiy0NhRK4XzH/F3mxuopuj54pHqvmPV1ZgoS7Xi/mCeqwjwK2PYmniJJlV7/nCC1Fx
Db9C5O43m5hjReHBkS4zYEbLtihvgirVUF6DnSNl3if6wEd9abyYEb1QW7GS+SiWeRhGBSMlH0UD
KFYe88zAla32sYb6ze6GtGBCzQlJ4BfHphV7nwsl5AKxsnuQeqWubtbMzMKzHkSkT7g5Sd+bjdv+
KVc4WAfyOrlp2NvV9DmZWgDLS77G2P4PITViA3pSNcNiTZvCui2DTNUB0KRPJKYZqFzZxZ1Kfb0m
UPn8f7PqXDmKDWFrKjZH5pZsLWYmT12MSep5HIRBnITjEGS8chHriLFHU/exQblv+LI23hALBE7H
+wUG825OZJHEkVpNrxo3TIVrkcu+54BWVqoRocZuH99iYU/IyGJXV27f+pnwexPZo6uDuQTvqQYT
DvPyT2CBgCGRfnrATQxyiSICP9oz3Z/Uu5djzM1FIE2pON8Pe0dLhRrY00HCLp1R9Lv7OZImrAqL
cyXipPwEf4EF35wyryLlnuu52kbjDQyd4XSmtbHGiZAYZjfxtCHrH80G8Fk12gIIxqNPVkyhsd38
1Ip4JytP7snSA0dbzxA3NzA7cjs+qtKrimV4f8qni5KLpslAYfxNtQ8NA4992CaWpqTLV8N23VOa
Qb0CoV1hO+wKnsXAcKBgnd5Li3O/hVvm4oRQtzi/gx2h6cOGTMnaLG92hDs2FclXU8QsTlNXCr2l
uWvwUumNG9kuyFK6+4i6P5V53aMIZr/f1xwUhXQyO+suAtQsAm4fFa0jP0AWC1fmyPlhDuByeFwr
1zm2l5JFxIx6izFLHLOuTHf9zvcqXV7rsd/Hy5Lon9gLI9FjJgzxY+CZlttfdSGYm5ajBDbvS4F9
U0WoJy6fcC0Np5a13ihqXOnS+Z0ZxNS5+Ha3Cr7/6rbwDsHGr/psiHjr6ZvQBfUYJsWRO5/UJtR2
l+DHfaxbE+Y9AZGUrw0DTORRgNIgz6tB52vamFN5Cb8tzQd+p65BpgOnnJvnyo+jY6jDj9ADPQBo
J4HlaefFt6VlL1xj/IhZn+aHrJV6zlCWLIUhNl7yKNrUPK+fzkymwiDVbuK2WyGlSw5+yiQCBpKN
w4OMXyx83YjwYhqHaZMQvOk2sIRIjR5SrGyC0mceguhWEp/jwf3V7dhgI8jSnz9KV71mCLECzp/h
xqCbToJdOMwm2sR+pzhtZGPF2toZzUOZ4wowrDLAs8tFUeSFJBnNBxDKIOEaliuPhwZ8YWqUEfkr
AVRwty+T92WdSAH56wWsasuB1q8mQN6GAvJyxLv2wLKB8dGDecGPKzHFeYIzhsYc/lRqk7y+3Zwd
q5sZ/7cSgY1BvSpFg/e5D9PNv72Kb+vcP/Pjj1Owsd/15WHghkNK2lHud0ocJnZfGPjmI2aOde6n
vtrifel+ssd9bGkAEsckOwdQgcxHik9OpoDDVAfpVdo/dTrlk3ZxjDn5MZTrbkDn7wdjvLQYhtVQ
K30kFiNSoS1P45+ofwZStjTpqLU+hHZFgwEZc4ffKWEYB+sX8WeWGaLmDjrmz3ZxrWSW1mlIdoy6
nto2KGX/vP32aNfRSooaBWFQmREGzGISdXaZbvi3Ukk8Fj6sjQlq4yn8zy4EQ4FDhxto/wh3+d6J
lf1YP5LP/KyUiRkBL9n+euIgv8Ub+HFAIlSewCNBqstPLn1kC5Rd96JA5do4R6PNFhZM7cykT2yd
rZiXK29+ocf5ZDeU5SfR0Cx0wLurfaesr/kq36k8RzTitRyiga+RAEJa2lgK/aydrvi02e3XfPq+
iiIqCGTG8ChItFd6C2xK7RY4jOXTjKbBPvs2q/h8LYTaozRKcu4P1fpOcyucboUcjnc4HV4gJRdA
lLqqp4D7T14CqcNMvYjCXdd++kFlyu8HO5gl98ZBuUVVU8VJEAdhHISclfWt9PYQP8nAcv2zjod0
Fay4mtNoxnzRnj/9Aex4Fkkz8v8/CRi9EK2WA6AaBotfYi0uq/nQ7c6sOcnCALV/4kbrtD/tJHUf
1N8Zz7ZhFem+TIakeYW4crg/4yrIRAOg6xLLHwT1TTTIteWwmEV9SwB737zRwy9/SH5qP/ptXbzQ
Y0qqYc+tfECRnlkqXFGUdE6lTr8zKfwgWYf3HKf9AEfcHpfzMQNKw/3Z2ODWAAYlhQx92RrmGoZF
8JmnTHVVWQpgl6nD0sGVElIbs3e1jhYo5Bc/N+HYFJop61P12xo1BuVoOKBEL8r/wbcEJs9TYm+U
wBqsAB3pq6tBG43MYvqwr+soigkTYvzIy3u7cWdFbI57XzYn6x/xbmDNB+SKGiA364O1++Z6RqfB
+0HdSIFk3r5pFlQkcbka1zsu3o/OMhC/+woZ8t5htLc0S9xbKADr2ktq9C2czhU7m9ea2cvnqX70
k44eRfFSgpZYSC2SjAZNuoIGzJqvlodUVxyL4j5sTBLlT6qBzwm0dvmnpfjepEiVU1+/SUmCXHAU
fW2e4y9v9mvYUgjkcRBBKw9Qf1nRvlmlhAffZ0WU/16iPo+r2BvlMbOc7lwK6GCQ1XgkTrl61C6G
OL/z5FIihjTaW2L6O40V990jy0Hb81efkbiOExgrGAneEsH6XWz+8XRSTXCQWy019KXYxm3P9MX1
PpSudHNPuLw3HWMGjFVU6wxjP0lBhB1pdc6nV4KPbO9OFxFL0dz+r/Er42j2JewERtMNZySAwlSY
U7dwOkVY/HbwPlkydt26vKMZOw2y7Vf4VsPEln0S50ZYlFo+fJgBzKlP7OXMivc0EkrrwHNXjC73
J5kI+P7Z4/W2vNe52706v+YIfBqOA+PYVhi9XjwPFLvFcjeLuBzhzgVAK+g34bzTGChWOB8wPSnK
0OybxORZ9Bri2+5NnCYgBkS4/fQoVxq0aOIgfaQFRaOMZNDbVrJE42iI74mxPSPJTFnmVl6gzRgf
6p2VMJrJmg6ySb30LfJcWBsOqcbFV6zls9iz5q5u426gf0EzoUdcX+0MwTrqKOEdlJ3gMlpPh/Up
kIwWpO/ZHY8ueC7mbg5pQcfdW8p6poQbEcBtzjOEoGdWmC8Lbsf2Bl2Z17JeBUel057/NWJYWYis
X7miJyMajjwkWHjL7d8MwRw4Fi5h8EqPcE1p+cCICghKIIUlqQDqGlesylCdXptEL0qLFvXV9xMS
1LIOXnjKZtsymn9BtRUgdL0C1qMvbwr8b1p7IMwdqOunlQRFLvRGfYd/X5IDYqNaeYPXqLTvrZJx
VviytqgJZZLfXMs3cnGkePM1hKEEC5funilLIi75dG4+6bHjt3lI9p2SGDOtOyE2TDYNVIp8om1N
4JkFkCkdBnrOZFR4pkDT5lb0FxBhgEtRvtXyhrfjWkPzgoYzbNzsdLKxdhsdT8k7GV51+/u9ldle
UWwXY8iRcdqTaV8NmjO5a2QOIvW91XMVfkl0H/5r999nuvVFZXRsl5lgcRcmbwsi4KpwVcCyeLk2
u4u/JiLr5DJMQo0HbYMc5B6EGQLyeny+Lh78V7SnKmp8Fm6GlT2iY494zc3an4n3dHXtCmRM1Uxm
B42lVZ2+2dQu+5+216dyxlwaA25aFwYcNGl7WRreItbiFRIGoiWKTKnl7GHxwyfzUJoL82SgvllB
BUhw97i312pd7vVcfGMHgrW6sWsZD3Ifoj7Ea7OfS9gdBr5o0AJHUFl0QiJuj2tTStJrb3xMh+x9
wxi+vyu+i3f3MDJezKFlhFcht49oAFskGcN5CDFIUn3DLZ7KlDwgH+xAti+PB0qo5z1OcKRem8K8
AQH9HISLfG2fktxTsxLkMag6gR9A0tP3Qob5T8Adsa0JZNN9FCJWKRzDB09RFMnF500vH8lhGEmi
Xk74GNSnfBJJN5DJRP+9/j/Xxl2z4W2Sk6MzHAAofTQjkwjvTRG1imE6A8pySb7MHIRoGLOGZh61
d8M2xAfGIYdN12fqE8wKtdqrvRHvLb6Graad2q6BKLGmFtbRC8YC6+btcKNsSo0wm2Xt8rwyZhLu
DeVwwTYX7kd/q3J2HEiEl9IFdU3/YNleG0F2k+6AOKmk8uqbr9qK8N/zEoz8au6Ksd90ppqL4xz+
mgGwP3t3e0wvz9FNuvhnfmZsnGSHiYZ64m0uAtD99uFLDpDzY6MfI5dS8ZATI1SMpvXzJn1wjmLH
S0kf6m3q7d1V23wZQ9/vOkbGdk6PJclagO1NuqaoYAGfx49lsQELpuCyi1s1yrlM0doCzrG6Ya7g
lC8rsSVnOq6PmMK9BR1IQfrIsTtjvGOruj9KHoNDobktjrkL5odNydhFrY/9YpIrWqSlHTTJfbRT
1lB61TV5ea0PAWVXq8mBuhD6sumnlDoDK11MpyXn1YQQ6MSU5flRfp/wpZh+1WbOb4Rgd8w3liNn
5dCF67CHYNI469YnUFrPTtFTHsqPk3SWrT6iyZ87Nt2yMdlW64G8/UZFBeCpcAq/DRZxOk8iTGaz
In2ZQOnOt29GL8vh19u3Wnv55SYAk2iNQ+0Kznilqh/OMinOKdR+7kaZgE/JL1BARdy0Oi1Iefyj
jLkMozhe4SFAoQ9ogsIA1ofeOriP27wL3EE6g0V09Td44xvmfdG+m02gU+m9pwfCCAUuaI6OyAoC
WcANonXNAsE6QoRXPwAPC/uzVDVDmUPQThdbNiYkFJTwtR67FL/PzZtUKWagFyoxQeoThoEToyvd
TKxEGZfsN0+yANLoyCV0+mHRPrc4uz6Q9LcEfv0kL3iMajESVhz/7IoIk4ZHfDjTyUMuYsnpvHEm
l3sJVLhDvwYIQCtGv2kjYww139nWoRJhqwPaFQfMdk09bIXOxmw/X/iq4D9hIbWRl68RIpEQ4YRA
Xw3c0/bm6LNMoRvttUfQNkd+0Vq22OlNNYvnAJmZz9AEe/AJmNcTkyRCKjCU9LtfJXbtU7FEM14k
9LYLvEu6mQutc3o1I87V1yg7foXuZKUVkhUc0T8sW2ti4QIZ3SOX4njAqt16fe2/B4Rjf1HXV33R
GxtiCy0HITkMXWzCvhBEo5MW7gha3E/msR2R/WQxxKHyF55ZMHbtwIbZS09IVjmNPO6SFOQBW98X
1ziceXuynAruzbfxiDW1qRuCbu3lCCcyh2fpi4Du/Za7Eb1SYn3Dkv+gpWm6zAxcwMt9r2aAY159
IsjqehiGrmRT8QVTySwCmC7l767NmvuLIBOHye2wYQsem1OcDQ6rc5+jw8wWVu/rx13+poYMbHRy
77nGbjnZkxckHMe6P9y/JkVpOHUc4R4e5h7gLX5UF3X+XhbzvwaWiWdUCs8k0QlNNI5UUEn3sWuz
703lyikUq6dpWGTePvZzWCUXf7Bm+CeNR5EbKpqkbMXb9Io8bbjmcjXO5YDnUb0qHoSdwHigzPqE
fhDdAnZkDC8BMzhII4F+2OICrVL7Q6Sks/kkmdzS4NPeeQ/o3KVlHs3n6GJU5OxnnGfZN2uJoI4h
YbZI4ij8dkRYc2gV9MeyLCZfunikhMJaQEFYrLC0crgf6OUkXK0/rxS/1L3EY+UL8rYluczjaCmR
vsycqMJEiJKowLfpgT2n0hDT1Er57u2wS8YcYqh8QnveCKIVE2AlvkywOK/9tTyAyciNdUldbUhO
eIuvLX9d6NAVbVY1jDMC/Tt8U7DXe01/NkvwrBIl0CgaHSo2o56S6H/OAhnu1Xh8fPX8dGlyaEco
XNdb+YWYI/RYFE4dzluM6QQVfMZ0LUfHHmSK5nxhUUM1Kgb87BB4JlQ4o/bHIijDrw2MgW6aOlmm
tYiOckm9DPWqDqW3jMiy14USC0JCeJI96g/2P/UpYLHwoTmiJUBCN7rFel3ZyXyeToeNZg3ne7zw
iKLzPdujs7L1AALlPkijFHnKObm8MZ/Q14JWlrGGLWlybtcMX2pf9nCqJgOmFKJ2tf//Hb6iKLn9
+vhopVuEp4clnXIIfX8lbYxyZNFcNkQNDcbseLvzdXvHGS2rz+XOO0bqDDg251UFEiRPxAAne7Wd
gck61NFUegioUIjBNv1zpbYiuy+NBfYzLSrOs5WhFK6LPtLXPTuxAxqDT5/XLGqS/KlIX4DA/qod
7S4JiSnIa8s/tIpFJRpoRhjDGfjpkXREBR/0onZUHPuRRAqa87LQ0AU/m55dozucdP2owUKgSXxY
ugXlKpeHPXPKj6XGkxNNgwscpCAyh1eVq2zPMPNpRbkPbqwokKa8Q4KgLQ4g+rmczXnbJcTVoGWx
n5RL5iJP+mAVLl2ZC1XGfX8FCPoMeqPDW1bgoWaCTAZOpD1oPV3BKrY+BFSnw+YorUp0+q+gl+Yp
M43/oJ39Ux4EOZFZdzVRbJLO0CGw7m0XiFLaEPJoTBz+X0a9vih0OIj6xzES5VpSF2jiJHzD/uCz
yn9OmB6KyMv5KUyXyrO4QnEN8YDNCGyW6AqGw4h9UDHXqVjuoW3EOhrrwL3Ue9W7Q3mIRt9XUYVH
rUj+jbDpCvgfLwRKiz6iIeCS/6BfK6Kyd8WrcT+xLJmi5ATTPDNyIOAWZmyaJh5y7bJi/AUTmBQS
IMwBuHlNBPdTF0Poj7Ueu1CFj2zqRcfPI814xyOralUpnKyiodhTfIRnwinTcum5NHOonC63NmFd
vSOZPRG+IeVzG4SnXy4gp+1bLN0ov5yenuntIN868uNE7nzv6PXnwbHzhBFjBe1ZXiFQpGB41hYr
2JTkqCvRxvRTMVx/8ut5czwu7nlgkddqPl4jORH2q0c8BlrKqoIABvBmDP3IV0kM+WEh79ODzNaM
fO0kJGrmZf8wRjH3Bqp63hGV89+yjkplV55+RAQMwxQn58yJ1wSSFenoiiUTQqhmO7SbCPBCEQVY
As4vwqJhnDgZGuDaKort28c16IOETtCDUypCZ7aqF1I5yn4CKtEOZDP6sEIhaoSzXqE7c+Bv6cAf
Ma4vjeQeDTnaJWo20WTgj8u9EDKDPhZYUwNaTMpMr+BQQb4SiWU0JC0wSXxjPLCxSXIMm841jyeb
KYsezOu2gy3FgALZe4Cqt+uMuJ3etpwxGIg/w7dnAGa/2+IU2kcqEL0I8Dh2ub0QmRBF0/lkk7An
ezlirjtCM6k2J23Y4tLIgtA5ilBDcDpC4eD5TXgBuRmX1hfTHAOxFHyaF3ojjfwCqwEN6aj+aq3c
Sul6/2gsfYxf14A1V+hPhtfC+LXcg0nxrXvLWr83Lu08R8078wkVk+BSFvX/DeH3QxNYMYQQaqr9
SFsaOvdhxBrVUTgKMc5wf286n9TWfP5V9WCffUqXXv4suS9DLJPkYJg1een+z1sK+H63eEtQPfcW
yJljn7kcCkhVZdLqsoBhZUvllAZ2wODVZyWhMhOYBCxIt86AmQmvXYGRw7dSHPWJbWcz+IsOhLOJ
oZ/SlOIKYYAwN0hMZ1M60nj5e0TnkJ/wSRgMKm8rKWno0qlmsgj8+dYSh/DN4o8cAKnVosPTeFGm
zVyx1chFqN46XnfkKpD+IJYUCwEg7x+O+Ggn2Hr209teDFOvVdZXfbV3UYMiOy4yXqW5f6A9xF7W
5aLm1U6vEY3Idx+F/L+XeIhycGqsBEeGvOQleJ3RiCxdOWz/oJdavO5CK9NncpaZwQ4KOx/bF7Tw
Ey3G61stWEQX24umHzStCEdpGJ0s2rWRW9OVUfF2mrjWwJvyMbqINN8ysklC2UntrhlnurLNNo8H
bO43HRwsY7iKorzH2/oYGOX7oqMCWDvc7QC1DiJpgAwXJaeE1QolcDinFV251xzOeDaPcuhKepfY
7ZZkbdI+zAEStQ2bl6OjmiDbnaeHS9DSOvqJqi/0ouuKGkpVAF7n7xytXwehj3coyq0mtCOPL3Nl
SlxiHFvxK0MQYbezzICYRuNVMB4+HLkYnbiRkz4d5Pta7eGrF+5/Tc3CPkDNqz4YYxNXmOqpzi3z
NOLNXylrEpj7ut05QW0jRg1+xk8inZZ5qShx68qmRU+017lJFSNQroIsqld8VnjdGj5BgOB9QUeh
jsnolsqv1zlqVbkMO2Qv5q9hVf7tuAyHE/qFvr3hATTqwBkVwn4ZVTGLlBpADmRGki2e2KwFZ9br
2cjHFvAnrR7ftrF14T0cJydFHPf14oo22fKSDtYTPeNFg2TFVG2CyLtS9KM9Ptk4qOJy2z0ENR2K
nXyGJ6P4dc3vc7Gl5mBWvH9oa+6017Fh68MpVUaUHXtzRbV6HU8MCJKUzWAJHc8c2xK8f2QN4NxP
OqN8EF+WJsGOfxN2nFI/QXEb1WPXt/mUcJNJYm4RunoChGJ9SiKpRKkqvaNa44/7iEqy13bo2CUL
DfF+Ja7jvdHQmGPxHRslSBgNc3WCUhzgzWnjogVkF9ZP9mjpwhwy9kJC2NqRvhQSXxndlpX0sSXr
yKx8+uh2kSmLkLzq2x42SgKwxsNFurf45tvi0zMRSXju6vSKyAjaPogDB+gz+2ZzMSxSoyucw3wP
JizEJGAs7l9OVdfCwb9pfa24qSTtgrHKmu6fso6QOsoCDI3dZQ4CZqFkDtNdUF2nBlSdUvk6ASmi
PWM4iDeS8Lo0YHR/xtFfRq1oMEvrEJ7dwtf8J8rY1ZL3UySQfMU9nnF5ubN+IxnxJuAIIPpuwkgp
NBWuL9QMO2xdPmYJXtIVsZjbL0HhtFcevhxrbpKbLHv8srWE0RTV/dDMQRiNlhjdl/152GcnfIqV
lNCW7FqAJSZh1U4V65SMudcOqcNmg6oiKfcHqS/CVi42xgmKDl2L3s/NlSr78ZcvWbZJmmqUPCJ4
MrqQgo/+uVBmsrvdSGErsQpOGTUjUioLjyVXzxnui5hxZi1ig7kAuYN8gHXCm+xu4M0Nnrk1+XQz
T47gA7mCDLNYwypHcY5x9OXaEFdUSN9NkAWQliecW/GX+6ZzwGxgSgl3H3uLcdk44PKPYYZ65PHj
d2fXcoXM+YjgQdvwc+ZDdGLn8HzitB6yBBu6Vvkxmv2z/ZPooypD/9+OdrqlkdO0peKxtHXme/GI
QXbr1EYxaDXl6OApBKfPPI8dqlsmw3ij/Lbzxnw9aXNbBcxFQD/GEKk7jYOND2NA8sURY8uQQCep
eeR9EimEkjeyl7DV1ZUIMefMmD3bmy7ndczHDBuflpTnKcwB3q6vHCN2YrTcqkJlY7P+LgflkR62
aG+SEHkk+rDPH3finf956U5Airp3AJwQl33bR1wlSjeau9mw84+npdu67l3dwNgTX5Vu8cW7Ez40
697iLEelk6gwzps1zNJgdxnYgFJMCc9Q4xy46ZzYLOa7OWJ5izouueeiqalZl1WziSFUWHP022NW
ezyTUE3pIiMcIyT1yzh0pWp31g4JirXsu2ZCQpKfAUD9VMSWYEY4Fi/hU7JZryjQS1/z9LIpid7I
09B1ED2UCub9YA9d66stW9g+4UE1UTb8OmbFRQSXfEgr/okog1kiSKKK/4usaqeGCISJ8zvAvsfp
OnTSQmxD0BvMZd5Mqmv1LJGqqxNXvSvSef4fvDaR85CJAxyrSv5L/5AZiG1k3CpJSZoeBKVzjiBH
SBSIr8X+Egx8fN6EzgD/3Hhqq6Q6H75HaClO35q2oaM6BiupPzwbePmlvhGeKvM/LNPGmef7ceA3
SDQZWlsEP8YiUPE1OpVlq8XBOpXLHUaQTSa6z94rYQA01KrBFp3tLQXLqRFYRZ/puXwqG5lqSXbg
E0GFDMlLG3EPNvk1b59PF6n567vk5IvLTh9INJyAb3RWwAAg/83dkYhfoiPcBpexDfsBxH5d22Mc
UVJuyXG3F96St1SlE+YDrEIhkv+LjjjE1Q6tllE1xHEzV//JgPGtduojnr1SeSXmvWBUikrHyGGn
J1STZVfchhZQ7lT2aITJa6dZcOo6l3Rbxz2vyrhQL7o4hl0ZyWiBJlwlGRBQCy/lkD7nimGCoBe7
NSGai3sYvbCSNoKKrCnsycmnCfJ/eXJuUoYQiEOB5NkwZpwiSVCC8f/E2wurQ1K48wn8ZQksYSwy
c7dhyIci8kKn9c5pbicZhtEPVwdGFAniyHgSoAg6g/iCwiKqHpG38M6y/SqVkygSwDQNBWcysoQr
7S7FxULw/l6D6RMxyDCAUoopevbkxtYaydZxaCUxxRhHO4md43T4VXhXAVH4wk+tKmnF4mZgrNFD
/wFMWkb9W9un+C/m3B8xEbWbQS9UDWGfyAu9PW5XftxtAGegyXpuffBT8/ZKN0vBMnIemUY5o2vc
yPSV680fj2fU229z3E7/INry8xXqHHiJbDPjDgD1NT6XLBvzTZ0dACfbJrX2E/4ITkC0VNvWotXK
q6U0swnyjVsHfqMAIQoWd4GQYeeXLNpNBL5NY6/2777ddbYeATYL/+YQtnWQPQg26wpWnCKqzZvk
U2S0PcehjKDp5v7dsQCkdGorl9cIMZPCWtcjo/qXCokYxdqDGdcqAt289NmarR9J/kX4En6pl2Ev
O21VnQbgVGOV2oenP7V2Ud/c89FnOBbtyeJD3CCoMdfXNSsFbMN1f72u/ERc+27SDahEnSDiYx0o
JuVTrE77PJ01jgP0khk5ON8KZO68CL5JAhVCFGCX8U6/n1xFtQpB566NAPCK3GvQO8aOvbGT+tfr
hMNSBOexJtLPmMfM3l3SzMZK79/uqYfjNxU/QsbqZgNEGYXjtZEN36AYrJgThg7R6N/1PfNqNC9u
lRQk07dHiX3LO4lIDySqCxMzfUdsxOqMM1GTzxEfyqR0YzChBD7JOrV/PMOSmt3xiZWQ/bCjNecP
BgfdZZ6j2e8ZR3jm0IdrB4EfNTD57yTc2TacdtxCXYiUf32wPPCBQdl2RFhsAIxC/dch/uFM0qFr
3J5vHjvjzAGHV6CKUumT9amOE4lGrcPxn22595WN27Qh/TNzZ+pUBX97V+Ldllyc5J9Fk6PjCTsE
YGXtcJ+USi3+Nj0wizy4icLayBIJqsK0vGO0qrKNRBWKBUDmlmC2TogaQzSU9yb1rLneTWfSuVU1
RtxjHK7WjXzBMqRQNjsasS2/PJ7XsBr4ueygCAFuYc763oP0mkpt/oseK0TIQqWXX9SH/QMBfNug
o5MB/PdRSWr6josoyUhpCOcLY3yL+fJ1pfA9djhzsmQgOGUEnBW11N/hT32ejuprOl0njiQNaY1u
kWPsIzVfJFZTd7vnI916n4hseCnwglbe+qn2cNH1L7okpGcaq80YZFDC7CAxIcIBUxArAu6EZUcX
463/d2M+gWRrPbklungulX9welSAc4yoE5kbuRyIOjHm0smw3pqm7hMovMTXKFNKx+TLlmYVWP5j
Q9K/VO4epLI4yyr6cADK6/YmABAHxB2yEjvZ4AntBQvUBTbd80SVyh16yCXWnVHqKO3bqVAgtJTb
/IUsXzv4kACTHjIqDQgxMJSaZ+VK+cIZnUQks2B+EEHspu+nAd/n3ZZy4jBPf+ycfHyNi9xxiyFk
BTjNvySaenqLKS23bUQLVwcoslwu5h+msP9N32jLfMxWxJMnEY3W0JknxPvRq8UHJcnHNh553DTF
tF8G61KThaJbDfmX5fv/Y0XzQBhnPg2Sm126qomGpY2cBPJuqObGqvspxduHt9p75Sd8dAUYYXQe
bzb0lcXfyt3EAq0St5NBoW2rVttlTc2NmZo6Vmzlg1UCaCNaL4Vh5aBPuuxg9uz3mJbf1SHCG1Y9
7kd0flz9kw6s1mk6NO2KjTnIPgJniLXT8e188jTP0mOhHITMbetyLvBypHK+A0DxGpny+J0DzqTh
0gHGI+fFNZAKwr6eD+siLLhWq6pkYtVMPR3kYVmI3JJvbHv16ujt3LYzxiavRjdwbLZCVJCiYBqo
P6BoBzmPZRm7xKEQCqVFgdVz3tbvvoZnXN1spvDImBbBe2m1mO0tWL+oAS4ptFyjJxHCwwl/kGOz
S+tyb+K6Dls8viJCMyPHVnnfQUHl/bhvxltyVHBORMk8Yay9u4J8O46qgA3/AVUm5YIFXsyrLfix
57mplrVDjyLFFiKCewjtPtamMrL3Eys4VW46dNDjmYEuW6+9/iAl9NTTA8fH/A1h1BVxlR80L+UT
8M9ZRy9QDyfy/5V6SS9S+wKkReqYN8oJkbqWHftIKJRgZz3LFRcKMmbLe8pWUIdfrP9tPjv1MlYP
7WBI8/fZx/1gMKxzz6XQPS1hRLFlx1N1pkpIu/vGCaNpsMB6oIA/lQBAtWtB9Q5T1xM3lERwJbk0
kW6pntkFYI7bVeyMFGOStciPe/ARB/OBymWGm6vmqwokUJeroAaKo1yE/Nys+kMqW7HSL6VaU8lQ
hJDwUyIB7WwYmFfRJ5CMd823RHn9MgKCiYHESClmcze75XIjfLxe0kmdBT5pT0nHOUEbRO0R8pbV
0X9w7XS4I883T+2ABjGCTItEc0qU2aKFwDTGjscRHTLIRsN3prLpxprmYqad89IVNVpvuS+70tPU
BMLnPUDPYfjWFtLzGnj84S4utpIWGWWY/dw3iz1AScW+PS5oYcL8A9p1iL4u4AqRqdb/PjsG8nYY
xro/5rIqpkBD773g1MOFeymLS4u++m/xPKfyrv4wIHnEhaW6ytsGc1Wrt/7hoeIFysiKEzoEZ+ei
TtIBgM9vRzb44hO/zoUtau7RI4vnjAbueDJfc6S7lh7IMBXZhYuzE9+AVdTE7/4JvkBP2x4/+hSP
GpJVd12ur/zJ3sOFgThOxj1oiDh7SkNO9B60Gs0GdMSwtUQtiAwyOF2qyQiNV6yTOmYyLBOHyncm
GIPGNKPH4BbIEIphcdff2DiT2/yyWziQtPutvZVkJHZBHnMFO7Qs+3/pbqy892Dy1+EohK5UWUCK
wC2z3JIRPD4EtTdOEP8NnlkzaY1NjYuoZGHdI5GxzhM1zqoV7yrg6+tV/JVpE1uVUfW7buFTY+5r
3cYQva9wygzwFer+lMSYvqTGo6eEGe9xJx+RtYIiqcOIYB5XCRpk7kRXTDYB9CmKpl0Yeo7oB9TJ
fXesFeLODO74l3vHn9PpqwhR+h0FwxIUD1vTasox1xTWYF3RSHzpW+0J0wv1MezrQoLEG7Osm8cx
t+lrPyHNEhWZi9QFHp/PX4DG8UqsSLsnMLAOAX0cZ8Aeq/oOHj4EerIWlQ4R87oi3EzTEKVfs0vg
SFdM/SMkbhp/fzxTDrru7n6lnbESb73lchCg/OD08qQE2uP7f4wjBXjgeW/yixjGpmnufvgXtgXh
JLo88yZkJWE4GhWIQIz7jKb8fkhoIP7wvtDURee1ikWiDWL8bpthMwNiGLmuFuBmluqC4XZ1SqAO
Z3IESlIA6UCAPj1P3AGuSbp+x61INWyf0XL2fp5tE05Gxb3zxh2jY9qW1bkzP4ki+q2wNv0MQLQ2
dFrlAax8qC5chlrB+DiEZLpbnQxObu4xd0w0sgYUA/KKamCK7t5KQ37I2Fgkl0mRxVNAU7/XnuzL
MIQNyfesn2rcRkeGH1xoPk5a9RW2aDWl7lO06G/ZgMYBIH2+Pcwf2yXnMOXkzT22J99s7u7/7d/X
67VLXGKbJ67in747UyWTA3BQNuEeb3aXjLSeVR+XRogSZXkKIQ+1MmRs9PQY4LO8VIDGmZy0fZ5C
TQ05ULbBWNVrFMLewQowEgjbgkq6oixZT1RiFje/NocL0tcw/GqXfTxvG+3aT1AfwHYfBhf0HGxt
OR21K5waWDMMltZPQDTaLgDWlILhzaTkXPLoUAvxUJo1koxwz09GWhkfCtafX8cDOQB0Y4QoKJah
+8c4Nc0sm4e5tGiT2RTfetvK/7tvFiA2epLwgmQBhhczXbgMjLyMm+/Mgnxesh7+e15AH+3+1nnG
uBKF9BpIDWAfZSjeq033iyXOm924QUk4hfTSApuAo4FCdG0WCGGLZgOTbHI5K1A1IuuYih6F09Z1
8M5HyAsnXYWDmj8gHhIJJwkt5p7nLdOcMbNwcKmy32/8eMr88alwelXCV3Ex3jbXa2bPggn0C9aO
X1/sRtl0lKqTrKzqGTLVpec414hiWNFW9bksx75XRWd0UGAUJouAZ2PJ+RDyhn7pVWDv/NCCC3bm
pKcz31FWR8NSFBgXO2FJyrUjmz8nqdpcHMwkiJ22ATk/mZigUxFDzeZ+0ha5C9kja1h2R/Fz02kV
vmZp5EW2HLbgtxGnOaYbHgU8/e/yUf5r+uhDMXUVln8gaebg2gySCCJCoGCXQheI77bapbSAkmV5
FCEMKYtN0TgMMpH4Ipbyr4h5A0aNlg4cFbtdodqddTfFXsq3wB6gquSYrHJkWiI2ysFqIXIGT0KQ
ncKZ9pLU6zPn3kBlG04WrZSxJsRhIue+iKQKxDJjkT3gt7+YoFGjErHilSa3oZ5JUxx4R99ez1QQ
rxE6wQ2QByW8NHzfy3YYBn11SpeAHl6p6iA1ePl+IfprLw7QzdcEQH9V4eM8ih5FCGjwIvQtab/C
Ot2iV0xcdp15FEvRboCKVjH9k8xLNHUoLeXuinbeBXFwWlxZ3IEZ5ifrE/e3pgaYo9mI2mP3G8TR
njKCqMlofd7maQQGZGljlRGHxWYdlaUH/PbPAMen9i1yt+QJkb/4eg1RRyAuV3zAuH6CilXaP6Sp
9oseXff8NZnmZaEAvj7d+c7jLkQRRmLiY6Yqn191OGs2jwr0ROH6UZDG1YYRHSMA7yVviTR3yP5q
UuqhtbRtCcd3VvGTlD0eyt3PugfH1ymRFcmFBZrtYozeNphxVn+rGPEIFL4BVerObU/751MTfY8e
RxA1Odx45J1UbVYA/gexA9iHJjEgWFwkihXJlEGsrZEdd06/W88wX9EVZZH7Yqxe5LAKl117XPIt
lkLWcsxkHN10dc2w7FGaAneoXpxIDAVAVj2M2CONbVJfFCKlO6N/SRfPbjp9C0xbfnfARjblRB4O
k4DvIc2EtnBUkaSHfZyenKXDlvsJvOgOPs5OtaK72Z8DFkd/3186CQ6P/yU6x9z7S8wts6mLwrBZ
P9k8sDEK3mpC4NiVzQYfpwcX9dMJheYoWIbnk+E3p6lOQeHLBwWOkcnkjyD8vIJv0ameEFmc6atr
+xl5Dt+ZV60m5HblfCsjrCHz+UStEdtvyY2NWbfsrU380MYqpQAbyD5dBUcmooVereqq9SRcOH59
Gm6lSDQIdGTdpB1omvYvulv/Qtt1QElMpw6Giv50Vk9RVBWuBIp+okejkZdYpUuL1Htc3QzPOBs/
vdbrD0oKMWMJxCTRRqIG/1bQOcxnQxuVqie5c1SMlobnipsB5AGOQ9IQ22nvCYOiQ/bO+3s4hpQr
+hSM5PERjH1IGpV1G5QmOwZFpOppp7Y0vrR85z4Uuvwi9EZsWNaItryyxhfilDeMVMaGKRNKnx5W
5AF6EeACqWoZ6knkJFfxU2vVcHihIqLdgF0/lX9bVhLFNpY3etRWvlR0GspLLhPQ/EBffAj8nUsQ
JrdvTGD5cSUsxIdXtf9895I4sgIAhgjUuqC1Hvap2FU7qQ4tF6m03iswHBc96kdEEg6yeID3hey2
a2g9U12n+4L2TeHafKzW8ijp+cAYzfZxM/9EQ3cEMwbrQU5FZdfIYbONBVc8jDqwe1yIDfNxPX7C
0MNKaHUucJiZ0ck7nw5OS1fbtZBUSyNCXiPlQ4p4+22sUm2nOoNB/N430c+A1ivR7BbR+2JrV22b
NG2PmWB3uug5K6ZY7bj3m0eQtdEZhN0u8FnK5iouJMXL0srst1s9IFO40hZxqJByWYj7KhnCJUM/
BW03XNJnIceWFFyRwDLT7ZpWwz4g5AQrHZ+I/ffXGR5K1FUHN8mMI1m03WJ51dnPb0swIc+o6Eto
V8D9YOKdTKMdEuasEFXCT70+dbEMs2Poj511DTKuGoIlbMncKJm2C6t5s9VXLI3zwpfNYgVH+ZDc
dzyYFNE/zRxMZcCdlfMG7WPdv6HMpx+3AquQ4apxC9WP/uFs0PQaGKY6qKWqKyA542M78jEX+9dt
f+6mVOSe49vRLKNv1Ym4ov6qAfmYuSDmOXHaiGyjK0xOZtt0PE+LRch6zF1fWqjoJQntHeR1nPFg
5Hd7Aq9ZJpkqKMCsX674SrILWJTuRMYoJsqB2ZktXz2g+Xc3EPiINykqktslXnqnV4g2t1E2kDVO
8HvMCrfLLapGF+hQkMQRN973MsOWQGL5KDYpXvwcjV7LRQ17kYM/04avOd2MYMnsP50v3QJGxMwy
vq4XTZ4iBojAJX+dvqW8OnjFxhXkvoporWlhfRXTQWnp1WSl3Iag1scRkcyvM6ZDWggoCU1Z9SYO
i0Cw2SNJgMQKWN9e4ZJZe4Om3XldOHTa1CFZAHNQAkcNIsu4MDXhggd0pzjsyETGJ8FWNoXuzt6P
lL6GDaVCeswNhqEPLROHNQgEcrYJUMDdfZeuhf/KkFTwsPWo8YlmbRRxPQX2JRjxo2FrxwTWqufM
Z7C446hFboLK/6Uj8nvFMJYJQlMU/9FQlvNn/lwcp5OlNIPAKAOdlyCrGtBI6fF30RYSH8bGZ7cZ
pe72M3hky0GihftcsKF9djh4zV4BAyZCZSD/hLRHMVJEma5RHFh4x9KmwU1jKPmwkHpNCAprUylD
PyTsmWNqjKVXE0is6e440Npn6nfUDXQ8eX1WHt4Xis+Iz/eDJ71wyXgpLvw2IYhp0C7sWlKXlVEh
kOP2YG8aDZC7ep+MPnMrCPQEOXoO4dpafsUpf8II9yzA9AuI3g9oO+FQW6XPr5tqFcgfehN8r05L
xM/2Y85A+QZRs0mpY0BmrZtvB7AqbD/1XdCuA6AxQ4or7F6rd5FfZ035mR+mawf24RGV8w38andA
zAB18wxCkpP2jWveFy3dM8me1+znhrKBdIctGe5A22VwOfJT1uNKOoQjEuQpZ7PBcmTpzzLSk9b2
SMV6iBv4WvJO4dzr/5G5cNBb5YfA8Doh6l0siMjmJcaTs1C/T6m7Gc2QJLWuZqx0QGMQiGpf9BX6
iiIurplyfQ5DR3SOO8jGdlhTwkJr+QCQKNPQzOMi3jVLkleFl9V4teKcNcH3ub/7ZlixTh07UzF6
Y3Y/C3YgCimpb95qgucndOqLHwITX76g2NdOwXhnak/rAA80n8focoGVeA7XS6zDVYkzr7F7iCMK
AKPZuyuwXW+9/D0YlhPP6ATYasLjsyyk5fnv4IhviAYgiGTF5KeUqr2NWjjDrSEyCYim4HKCb6Tu
heTOEVvQsglroKCmaQnJf4gbkr4WUaSIGLy6AY0zoTGFy5GWELStvGaMrJCzUfidmEfu1rgZEozc
Pr18Zitjo6y8CPyF3IoFA05Ea0fsmuP1StDLn/9H9D/DEqB//SmbkyMIARLZeikvWrYG7C8Qm7Pn
X706voM8UChxgXFfus2K7Ink8pPHYss0pS0CSLtnaUE3QUNj7vuZb5CF2nvchIHFawtTi0+x8MpL
mbosAkdnHwjg3R0zERlVnPPlYwm0IjtVVKVbOwOH1ftdIfWgtaKrRzM4MCvtW9FijjQCoOEkKDrv
92f8G0d3Bdzwg1RZMbCN0Lj/GwtaG2ko4TEgB0D97vCDCE4w8D7E7X7fnNvcoJ3trec19gGXjS0Y
C3SttsgEnb200BFBaLXJVsPZriuvL56G89R1vjzWGVFDbmR//mzARgCnqJy5zcuaB9WBwMRLr1XV
RSYI6OWoDyW9nnWYeknAy5b+RMBMQnFItx/S6WvsIq6K5e6dvDPrW4Dhyr58rOXwbFfeZmS5Zk7d
idHFbnnvBcFxCzZOztOXowZUDd85HeQ8hUT9qa6WQNHfw48NmrOP9/HqDRkavYprCAO2/T33DpuF
3Sj0q/8da3/hVHh/HXT5a77hBGVlBaelcuCw8Uff05c1zShNH5TZ1GxR2cai9/l1MD00BBYjVFUA
HzHOjUTKSYM4CvFG8qdtLwT8/AE5RIFgypifbslXv0A2Dagu1rwvgiiH68M15cd6TWyTrsjijF8c
YHry+YtiKMf+Mea9B+hQPxmUTmPwhM1upaGjCTf2pEh6B3VVBcB9PupaaiGk3Z5TBbNeqOATAyYX
f7BDCXbNbultkMolZ5ztAzSyPnsIo5gMvAymYde/IxufPWhA+YvD0jL/V3wNTQqdrf4k/M8oQ+aV
qIEfbli7mkIqGB1NJ6jf/pffTvSF518UaYGyLEdVzJIxbFEmrRJ0X1SeYa3kolkkS6HsbSTg34Ez
QmikX7fOVmJ5xWCuFpqXNFIfzloA+Edg43LX1+Pv47CfKvKbfCmkSg7owEFFb5uLlak83wzwU5bQ
nkrRjgFugSz+SaxJcEe2ZjWmfgVMUqTqdgI1EFy78KDtyacfJNJdmmLf+XrGeih99tX2Nni+UxkP
t1SB5Fyx4njiyX/3BeIYApt1qRzXxuvKPH7umy4CCOtxwyEROfMJCq8mx7sRGOTJXnBuafDi6I3w
3ZJxZmAWvn9V1IEBBIvKLoc4zEs/piSNuECub5zoev5+zQCUaOdM4cKU3KsQNxZPazI89VrSDDAC
UIVTzEGwqRuXlGX0RbJxwhMpTUlCgb6o/Rdmkt0Irj+3mWyTz0aUhjFV2Oz7cyABG/nRpOFl3jKB
aIcTaeXsY8JfdpOGe7zft5WY07+7xZORiCLA64b6uDnDFzJ2CXxNx94xKwTYxP3a+CNq1+0oeRaB
9DKj+N/YBOtcl/NssgCzUdwDEFVjFgsJotwlD1bBTYsBl07+bozOFNo36O+cx43FC7blJLgvzjks
3sx4ewIxDwIhrSdQOYJmX2TY0pAdav7gSxJO8Wn76TrDa8efv1iR1JLl9dWMPFnL6y2J6YEvsyMo
wJlf3p/+bMArXb9jWqCNkrrRZqti6LWnMeyM9wgwJJBp7MXgZRN9u7xjmL/GwmE7fSSZNiIou9HR
pKKbRKN8ZZxGjTa1kCe9GB23gE/GejWwjaHiaP4wRAw9H3agKgAZEC9nz1X26BZUKnjxpWac3qwI
X8gweg++uFcTqrP+UIDwrnvQjYD5Js19LlP0X5kEgVOHQFVg8rYxFZ/N079e+35Ea4/5OArjwK4K
olcUwpgIpzZGF5eNBhNug+ad4i4KEN7dUPXAFB1zpis41xxy+NhmoFtwob9/MMeRMWI8qf7m89xr
dKutIgc4pS2oHuCW3SydbSifVWatUygb2AAnlUbhjJ7tvM8j4qSWmDiVcH4lIJEci1joe/xYYey6
0GjFCp+37BnTn+J6QJfjvT4oV9TrB9RgITaZ7gK3AGeeSAFin1WKW+8HbsoqWIxrBIoAtkVszVTT
ebHJp+c7qBn34zeaQRtEYJlUQ50VXQvdAmNTMXD6Rfhwgdsf3HGXJ27TbKGVjneRNLOIMxCQJ27I
T+MYwneg+IQ5p829UL7sfQBXfdBkjrc9c5GuSDppPQS737bnEvh9Eo0fEoBcgeuUZrjWZs81GqSi
c1270Lo8X34/AHNBbdlB3s6+1wU5NuywQszZLtRczBtut37n3cEAvd1qnj5fv/jbJwlqYQkXTt8M
ReqtS9svzogVr4AscPtOfkx3abtaiWIvhha3xajI1HYfktDJ6q9rLrnoDH0LyPS3Udy8DaXBUYa8
a7RA24z5fA/fAG/jjoKPfk3LfeqX4Tj0X7kOfjO7OHgwUFeXeoFAZnwH668KtZdz+1hGuiH2u4cX
ONhcpR2XswnUW/JgudnEU8KHt6swchF1bBx8zWv9PfCzUskCFK6wbLxCLUBtBDDmGrVZurvZx47V
7FUVnGHpSLj/uYmN23qqXAYQLC+35QxcfosMcMmxbiW1ZLb6a89gycqKY8DA/5QwIFUm8QnHNs2P
2ABsAKb9ROvyb5BAk+azBPnTxYM7COFqHR/t4XjU3hmwG9nb9hQ6fOCiIfXm3qNV8xj202SRaYVi
IZCNVc4T00ALfI6w4DLxVxyDIFTgjKokWjWZbwZigvgXHYxv0Cr2x+AQs8Ymh00T7xY6Qdl1pmOJ
vGpuARBnANnqhtxdu1AkIujsq68jWLu/JkJt8g8NQaPpaZFJw0GmD9975bd2KZuBuneG2JAjhNeZ
StXAICJOtQtOi/OwmZuxKPiaDb90fja1/Q5KutL+Eph+gK/9scqH18WQMhNomLPDTh6ZsymFMriQ
BNWw4s2Gq/wzZdk71740gGELFxZ+vLcT/YrKLMSegHjrvKx6bIdo+IL5hfy1nSplZKKa5zg4Z0SD
MEVvJ9Tq8hcBat5doE+QxfkJYjU6YrfnXOgsaVC+EX3k1V3ZGUUrUcCifkHVm40uQgBjcsmJprno
4BxG9XGcFEXtnWTMsWh+s6IsVIUWKr+bmMcW2ZhdsuRSDyKTz3FE2SysAl9rTw9vk1SIG7icqvEB
8PZBqrLXV3N8VDHnpbzypVxh/W00cW8vtuF5Xf/l1m597hJmYeJcaUBLDnb/xnHzA6/agyr3C4aw
0yN9HJ8mkJo8riz6zlGnsvqBrImp/7X1xXPH3qcM+z/+d/1rfJQptcrLQsRPfTlzBBQsJ1Bqt60E
BmzWlUZ3PycHTRT4LAy+QXLK84Mba4bZIwcpw1CZNZkLHPWIf5fNlz3NZI0IzfofxTlrE5vhnWBS
3NZGNbr5JhIw3dd/rIHL6V3jsZXah84hEGaGd+KFJEf/eYXJMPxL53C9wtFeJa3ksmWlUIoYP4E9
C3BZNH/8rnZxP+A8V7O0GxD9P5+AdXlAGEH5ZsATr2wwgloM8L9xtBTQ/CBWMsz/eMSnsI/OWEpT
nSbiaTkNgAKTFwidxjmkqbK1vHMxSK4uFE5pzUGEW83g7aqSxzlrRlGyMKw+yf11P9e6xQ/xzmnt
uDGQ8cY1r1sDlamCn0nU3ehQ7pHGaTB2cMpGCRSBYn2iqZZYBXmNSoKZTcqQYpVbOGg0WVaGKxsC
Ti3LJI35LpuZu6AYwcbasj4WU3tHonc33/iL8CpEXf+HMhlU4bw/WfoSN915PLYrxlQvGISx+9VU
oNi3dHNQQrdrSTh1BqPJuhjiQ50wkTH50E0zkRF5evBYMV92iQklUthDT2kxsm60f4ssjWIgx9GY
9NkHu6PbUkdAziDoIVzD6bwHLXgqQ7gLYAuABlwLjq6tO8mr87SrUyXXAKLWkPKo2GRPJCdewvv3
0T6r9qYsLgYcr/zaUhlJao9f4iFpIuvU1M2qpY37e1DNayJsSZ480qhzYekjEn7ihrh1Q/HT4Cqk
u4chMPojdT8PpCGPzP7KdCNl2x/LMMZ09T5Vshjxh4K8bavZp0Z7j8qZa1zJAGILNY56dssVYgLx
o1cOvwxKmYHMjGnV9VR77Ix5d4rHpCFsn7/a1foDM5BxYkEJw8RugVafHEVpQcbE158rTnz0ftI3
60DS03AB8Jl91JoslrmoJNmC2yoiBaKZFJL4Y7OEQjjYKRdouH2sjZMqm6XbwV7zcWgmhYNICvxD
O2/FkOQ3B/F/ZgGho7kki9qGW0e20a5gHANhMY5HtLbQYkvpNrJm2z5kKzOO1deoY6cXW/NP2ntT
RMK8BE4fZCYm4zsLt/sW/6utxFh6FkEzYl9dBl9W6gi5freXOdVbCFEdBGR46avp544k3HxZ74Io
WSw3mZhyQTc4oGwFg9Vzj0Vd+h7qOYIM+C95K0KRGhgdzNVJev94p0EXy/H5Oo+Ney46APmFep4C
40a3P69SgI4xLuOela9OJzzXSVI0PKE8dx0kXdO238LbixXtHYhDNWj8/ilXK8ZY/YIIPm+2vlF8
rZlfeM20ugU9BIGxBItEVFyBwCAKVDowR0avKFaxOC+/9br4+n39zlp/bZW5idCrYMhHYA9fYcFp
oOzcHhEtkBCJj2Q0jW2WGX24tKLdIwlQJlvfeUVbh1OZmhvmOmNMTH7bpANfBYNXkUk5nR7B7yYc
GQXM5xG1pzTNYkz/Jlhy/fYclMEWgEA9dtNXkAUbS8+HHpEqhT0496tZ/Yr+RTQ6iJlolOUbjSKN
Sh/m79slqmxpnhuDSD1Z0VdehLmXcUf1fFaJQ4+2EtI2ymto7xZRoxahvCB76mMXTWK6y4MOPyBt
MZaaIw+l4QkC77WjwwL860l8Dmwff0GWOhk3pXe4IbhwuKOaha72js64FvcsSORd6XjBXar7rdRu
WCKIk/EkR9zfWyJjUCz5w50CuyqA2PpKUyJQbyPr8WoqMLZ5qbWZUzEOclNVy2BicYfFjmdLRQyV
+j6K8P3Nsy4LBkeO27KuYd2P6GcuO3BlNUUxxBfqXIEVWqqOKA/mZnwkXwKoU0Xixnrpda/ucqat
E/jldWXiyzYJ/E6PmPqJU360zK0mmgK8dX7tal7fN3iT5m1eeV4KBC4wbGc3FwC2RaIRVAdXsUNz
UAo4StDNS0Irme2W3rYiKH868OvB0EWB4PSZJFbgOeJrIBpI/aK4R4TyhLuRpb9kb5wmJm5bXgvw
rkE4Ii06lEm9DbiXIDfSzDalAyps+DT/trIXpjaSym8tlxQTCsB08sAuodTUOmEkKAwzLY04ikkL
xugpraWLsjWbZHL/F2LSmjmgWogiP3vsLeZEbiETXihsEfFiVUIZMonXYmopvon+Yg3C1ccmrBBU
GMZrk9V0oEA24HBACYfaxW9Cl4tBl6A+RdQXnoIP0MTmpZL+nKMphslGRpkSp3H0zj7z7gpo1j23
P4Tu2tcR/n2XcJaBhyk791GjU9+H1B3AUOU9Ud4PEPKg/psfOnPmWQYuv661DIP8feoIfaAPhIlu
ilQZ8dXGK4PtrNHAJcbTRkSuisQZm0a/IZUXCN3+IvlveYUtErvjeGKeoJAHQjgSHE4/6JQ+JEw7
fW3axU7AorPlPUpv9EpitA8ftx3UOBPfdnOwYvIMwxUdCy9f+i5y1lS6SO3daEANwiYzai5qJOMA
EWtLotNg3N3nsdj0rHK4S7/aH2ZFqb02CzfQ9+x6Uw01+2p6q6rPLnZmE/f/YF6vRVTrhbP4IfzH
DRrzBLA24ZGnSRmKeiZT6GSY8utzUC/BpJIin23s1Metqgvrpja6yUQ915QAtCFTTo44L/r+chnD
YXqU047eFR96EHMHEOqlwCHMiCZMvJPFbpDm7yFwVAp1fISVzVqdZUdeDW7qk34wPRzTXGaVrrh8
aG18GSMZfP17rUNXx5HtJm6uehmnMF4bjSsG4VldHt3U0AdvN00usBwSwon8FxSVF3gPu6m/7GXw
t/cDhtA6kkprzFB5lwbZCDMzZVKH8Cmi9X3Ky5lFHuZwEYI1kRYPh/nM8bnvtX5s9yv2eBZmIVI3
Dxv9Xh7s32tHMaxN1OMc6syYT9Cg51E4imHSyY8qTodWNBCwafrpYofinta6sJijzjwFnWVgI2s+
/CS4kTnKbzjuVCYjJBD4snL6h4y33xQdzTIbVUMkxj086Dqa7zMxHKu7uW/i3/6ic3rVO7MrdEHA
SaeeAt9749rvE2y2LHgMG2j80VFeX5MFOiZhHaxq8901KRdj5pE9Z8yeCh0VqAAGJLSyqJxzy7LB
a2u2dxy/R5wHlOZe/8HmF4ZTlwkyJijHSeQPbI48/07obpSlgj25kRicWCxkkGH+rZvHJiyGrHai
kuWFBpRCFaerZPC/tNEleBudp+Yc73xV1579uGVo1kRVSR0CPBqOFiZXn0KFbKV7AVLj1X11xo1M
r3e64+9hz74XfPCVCkVBYe+PoLX6O5FF3Xr1zORxESWWkdG93E62ElEUjWQ8VrCa1lq5yN9x22QV
F1deYlW3JCNvB8UkQiWRKGmb15xtCg0G+5qCaGI4ZMBFyXmdRst/G2r9g41n9dl2mtZLy7IJXjVX
fAfa2OzZp0gPyEfYbBZa5u4UE4tbR7d/UPYI4i5oiTYlTFfhjYn9pZ+4r9sQacjTILUpnxpoavE/
OKyV/ltwkgzs27kT5Sw19fe+SMw+zdufLkctXqQ5Km4GP6gLrzfhEMcJf8U+iXjQGiiROD/2QPfn
+GKQKXPFXpBb1ywsqzCzDQr/6gXROHJrIZuG+9bTxetSXK/l0+XrtD3BgNEuskv0QfufUuquiAAW
yXZSsEs4zeUFYTO7v60F6OHcby/OgTpvxIKJ6QDbvQ9nEOW31K3Bpq6Bs1+fJ9Z+77te850QrcM8
LX9w67Wh9J3P3cA9Aed5JeP7n0KOaF2w8MPz1ykY52UtgE6cOCs+oDL3cbvwltNym/31VZgA95lR
RmDdwv178ftWRrEvvwdhd1NFuOJ5pRQtCR/Rjawpc4GXzee3VsrU6j2Sdu8HYBq/yyPUoH3QpyOZ
xEmw2Sb0RJuCafZMo+rPQwTNsXZUGd1DnnxBS1xNoJ52By33gUyiuBByunKlYvr9/d7SNdtbD7eJ
Lr8vj4a1GRMChCQyncvoFQduXxS6469Zbxj04Ifx+VbSUgL7ywn60EEXTOiFaHf1ixfH3aJiGGTb
6j1s2RFBSSgvWxnzS3gZbC93x8nzGKMorJTYgkWTUHVV1EwSPWgc0VNTFg30M9Bnhwr1PO6XbssA
DnBglE+sOISPApvdE3W4erlGLLQPXlo7ZVTFsogMLhuT9+NhsdqgEyqf840UV3nkl4EAzENJrC7M
S0/ARFzsdpd2/vHCO8qbCDrnkrG4VpFAjFv/GMqhpx20gL6NTuuVkl+3BIg42ywTO2FGAHsxd3eH
ViBfgLvMXG+gFtt8PY76lqLuDcFkbJL31piX6HzhPbUQgXkgP3+Q7XhG4P1qvq6bUYKwdTERJAC7
FxV31a+XbSOxku583HH0qzmrozWjoQ8U42LMK5wkJBA8VLob5QSVNc9v4lIZSx8NK50fDVI58PNi
UOphQV7AQ6JOPBsDaeO56mKreDjacwm8/rBWveW9LxdfUS1vWCAixnmZaKt9p4snKmKZWMJqFhNV
lEdAg96TVxOUUN2TqFWTY5ahtwYuHpT9BxUSWvQBIkiocN22FK9IriBU1OtDUNbCjJjFtWkDu116
GbqvphF6fkwvn9e+0v9hmelP3GZA50RZJXlIpytvh/RdJp9uA9dLMlqKebfoas31u3oYJNtyoV0G
1kMpQLDB/Wrg8NKGrj+p06buvFZBVrFEUZbS1THIwk+QEFxVYcHX9p9gXtZHYgQRYgT4eqreHU8H
6TMkT6Xo9pY8oeGseoEGGYOt4t6jjcwHjlv/NYTC8Bp/v84C7geQbTfr2AAjVzvpzVXn3bA4ejZl
ZJShaqMjnZ5DXeKXMAhv1aAr8tZ9+MVZtbUuV1BN4lV76KJpkckiXoJ1Y1P5zzMDoz6X5F62Rlq6
2UWt+9CuCItSMc4GVowj9pGyi+njPN1jVHbQzsPWhF69w5xjh6SSA0Qj1uBvKcqA19c6uQAWgX3R
a0k0ihV3QQL9BQVnZay7rCUACT/db5j08wiMU2hWW39ljCleI1kPDuuhqvXZRUi/44SU7QnV4yTa
jhJUWr0yAbRuag7WElMf20lksCaXJdzSDqtg2r2PZs3MQt9QHw7cI0og2ey/0WA5jC6kVcX7FF9t
PthXAT0m5XXMjnQpOzVuY+sPR/qYwsfW0z/g2jMNHOreBueDGwihtp4iBqwz9Kqh66QSzXizJfer
NUrX1yo9+pBZ210ginEYgVqesp/WHfE9jguViq9Ye1C62dSHt/y9JYERRPLGDMRd2bvjE2oMuJpp
nfeLWJ6bq/SA4wYmtbMXq3aUsIQgPrzyMTMvcEPq9fKk8BZqhrdAdEuRYLEoI9bi+cOp/gKcBC4o
jK0B2D93QR1BNaRJjxiqY6afLIQO1by8XLwwBBLUQiUU9t/kYvsa++vVJ3/y4/pwFd4gmhGVxXMw
KkbWBre36OV+U1iBUJWPYeK/ZhSUFLaxxXE/bHTVjQuUGDli8YLN9CNCETM26riDUqjUxaP4ozy/
tVMwCvI7/msSp4Jd+esJBhSqu0IXGdVYex1T+FlexMcmJ+1Qr0lnQjQ0r1eKi8vOdM1XQzkVMsaZ
FHlnqmSWqrsGzD3KmLAXtfMa/U0wZBm7Mt8GmLN0Oqdto+dTVP3IZOW9RKUvPaqzGTlZssqO/cq4
h1P8RahGTn+dd5krVYyubLik7f/BtPD5re/SAtIDlX4Q/0nyRgaE5CVQvAm6aOuRjsJRlnBLapSS
9ltUKYfWapJUQ8bAsXtAbL3FxKOLK4LdOapwFATq+zTCoo8mNKyD6wcox/+tMf+x/ujNYHvCdPCn
sQY5XhIcRkJfDBIIT2o1ljgI0JGWzNXLkXSKoSnP4R/WoQrlkw806T+iHVYRjOYHQLsa1TwyAx69
IoLB5tglj3Ki7dYcB22cl5Cr0zs+Su16OUIaON2pS2WukUo+WA3h6Le5fmFC5BxSesqi10xwTFUy
sgyws3R/0AKErbHeustKFAVtYjFsYguKS7mMQ/VF+QO3+8W5vUkMIdQRUl/knVrZIFYiyRxgg0Rn
hTbBzYpXBmzGZUu8hrIyIxhNSMelNcULREl3w7widucOiEYTjpt+YZKIk7pvdh4VIXdZAay9cJ7J
uR++/EHMYPfZuSLziDaOxURcvWcExzwGmGau6SkC1JOq6ZU0fVH2KQmxNktHCR0Q55uHwSUAzfT6
pj3mUIDpJy/yAJHAdL5QIi3oQIT/oSnq4dP3Ox2ry5XG7f0vfAoVhuRwZG66af88bn/7s/ubuTFW
Z9JvQlrRWi/g5SI0oYZZThuIzF0tisCGW2+FMHCwBmukbyB8oPZAINSJF2zljSY/sc2vpIhBq+d6
KW/nzFlbF64oyPVqvdm+4K3+qnq7/Hu6912EGW9MVeqE9N9/geu8Y8TZoXzUTjp78egplcgPSBK6
vp+LCZw2f2bbObC5Y0WZMSsaA8BL9w40U6WCJ5/PU5RvIeUDFAkELucAzdQu6iBli6LuPMEwCXv+
G+hH1cI07xSP4TldBR8CEsZFeBsf72ITshaBKlwCgXYDDL1yHzcoC7FQoK0cujfSJlxElqkQYHOX
YiW/HC7UT7+e5HgpXwHu5ftjJUpyUi21aKpe28bJDBeudq3F96N0DCoaL97QlmnNCvHKHW2qIL8l
yQ1h29aCRB1EA48YHFHszQfVqzAvzz5AAUsTEhKQNnQ+G4LoG3qROvnXkDRG9Nakzr+nCg6VEyW1
Enqunn1QTZyF7LxegPIwAx+9+TUR2AjmQQtniLIvtPGZU0Qv1p8V5YG5tAKp17elFBlfA31ekuaj
5qjFvoxCQfdQS7TbLDVK4dUkyRvIMgJ/czSfKPxUUrW8Hh5736p+gFjWgCtvmLXBZqNZKQCEbs7U
Koew933UbsIFGQCMYJ5X0CANmOjEn88pYkU1TCjUfwU5T7ujh0Pce5W5/c/sFGdHCVDbeKC9GUtX
4hRo1VqdTyX++Xkvaap2or+c5lIvXWrjZbTkRG+oGCSPbXVM1iHK3ybaxP9kpJLQ5+iOZmKAr2p8
fMROq9+FccYvVUyK3InlVOJ0r129bpU4613gqn2X5qfQvX8NoukeXj4TWn1nxubQuQWjdmRij9FQ
5QwX8bRMWDtqhhOBT08KFEN7N879l86i866kJ+n/yy6yn3ga96dRX3vCeRmeStiQnhAFEwDqNXin
yy2Z6DX+JLA/B4YhbOZjODJz4hmmiR7eRYquXs9GH/Xj2SZKm7o9+9vhGbS4yGmouDGQuu3ng7zv
HG4JPU8R/OchIcImPl+0PhWV42p9FLsNU2mvOzSpLJd5R6EWTobMuvhTjNxJbCg4P79I12y1TtNo
PH/RsRLo+qwtfyX18b/wNJ7TM7dwJ9NuAhiE5mtIMWsSnrE4IfbNv4eXUlZPAL0lzAV+ov3c9r0l
0uAubYmLJemtJaxEmTCkvyjvNFNmFCtm6Umksw0J229Qw1knL79hjTlEINY9oybuq6NTaB5QSaP8
Cg1TE5W6DCjDxeeTdASyEeNf4Kfj+9gskRLwwmapM941WEKA8p75khAIJvGYDPhp4rdLljKTnlZu
SCOMUAo0tgy1jANo5IbxcD6inooQYwLviAvO78qjhr88chiQA0u8jRF2Fv8y6FrTWCH+vSjpUjnU
7Ic4VlJ08Q7E1bM+qME3ff9Q2cmZAUGo2TPWgcMxWVMGvZXzH+cNQcx1nn4MJJYPxwI31Cj6nA3q
kT19MMhzzOaBQH7FEe5nZBp6ZG72YXk0R7A4jzADXpWN6SD++SUa7eyjSq3he+mR/hz5td/wGRGe
imSpH2scZTucd5WXNRWE8cb/zVqJx75782wN7TY4lEJ5htaPNuXkLplStfJBKhg5Sz2lN70hf3Ev
QClXDydfDxHj8Ah1QLqq+RM2Nrh98Dkf6PfSsS6lsB93M/ayiGBn629mOS0K7/len1PArQ3wI6Vo
as3q23xJ/P3ncD/EvvrZ/sqbtGOSA/qeg6ZCMtPA1Z/7VRuxjzumo+cCdVOFbCgzWrD4Z5wIuSXP
AqjcNWagkw+zbxb4PQw2p+OXfACBFGQUvRpn3AyuiIRHb1zyxlxiFhoMwUVXedc7GwzLUaDMqgfG
9GUkugtVS5tmynaIBKZVmbPYCe9vzTYRiE4lVoaVcFvbTOknHDPcwTg8ZuHzDTFeK1GrLdFu+8BF
tzVXcXGR9AijCXGuLDdTXz6LKtjn2sMC2PO5Wv0Zwvzm7lS4azhAPfHvp/pvAjKEyOw9mUIoHd+i
yE1g6YLrWWVMtdO8asmw6OBJsgTe0+MKHw+xzhig050lluoHbR3xc1HuXyesnyDgw/qEwupfyGGx
6Iz8SoBuEdkytKlbbY5fnvj1Pr1O3lucZxjq8pPHb4NtQY07QyTa5RWGoz70+/MsN7H+iBINo/AE
kFruNafOD6vvcIOuGdwEfgTRRlVUiiPPCAUeFx9TMGJlOQN65SVTRH3pEqZedbrJQ17FOKcWqCcX
TxNAln5efXdi5vAmOjlU3tiC4s0fHqHFJpjWlJSV8Lhqwyp3HuTYdUmXuxiqcGyf5KzG3xBlqDS+
RYfVVqXbdB6KmRyEUt3sJr0jsP3PlZBrwePNMry4WoH38Tu7aZPe+KtVxlnCRgJzpoqqM6J/5DHV
cUSRw0xhbxzF9qo6imstgDITSf9uCXXVJvBwfhIk0/mkSKFE3KbtgqConkNI0TZ7y1a90Z/xTUXf
zyofP7XEpgOdnSxbvTvt9kCOk6fo3gKhTuYB6NtZnpbiXBEbQSh9UNyn+4dXXEdUmGUnHKQzVlLN
ua/YoYl5LcVsVJ+1hLZPLix/8R2tTghJTBkDQaaRzfInG3RjCa6FD1eHOIOEqEw1RRruyBNaa2C1
RaAKYxLsulAjhdEOquu9pK6nURcW4+D+OLeaEJdEuS5ORUoJL7wtcykiQutiRW+0ETGuftJjqctz
P8qrlpaYF4AreszaNQ51ywgAmyzzMC3K1UkOnd3/vRAn9s2zVdP2cUGzg9S9LyEB2ABnUGy5rkuu
K9L38Mr6CI8+HQHlKaKS5fKwkf02dDBlrDoAh7oXzMF0yZm+yNukH561kzZstamx9ovrL14LuJtK
CNJZprsjQ65xdWBHjWZuVdfifJzwx6HiKp7S9DaG4i/zYSBu+XRUUA//c9H5/gdp6TKcQsVTtKi9
xlqaKEL5d4KUFiBeEvjili+jwxz84g1NcF3q5A8RGE45Mo7tSjnQB3NXaX4lGhOFXjXBapzClUgZ
NG1E7p2q++Weg0myXqk+ie4NYp7vynn18Gyab8vFoLhgs5zdQ377IvZ8AM2FWNsdYrqs2YtX054J
sFSI0/XJR/JW/OqMGMYa2DVmnl1K30+SLTSrvlkZKBn1NhoRN78npVEsKO2VMzDGRYsi4iyqNxSt
A/hGmYlN2GBdraSidEWVcP5FYxpwXCnDDv9UQJta3LqRBf/o0F71cx7WNDJ4m8REqaFsRw1xy43w
7AL042dZnDTVtHruKTu31i4XIUbZxBmdVtJ4b43Gwzo/t7p1wwlJN3avi68nK0HCS5Aqq4bFfJg+
/eG2rXpsd7cZI/Z/BAohiiBN8MWe4Vo02T54SLVPE7WvToYDJqW9c9xoO5XViWAJ3SwONLBxIvwO
u/SNI+vUK3YkiyxHlCzTbivsW/baHrus8GCazSeCGgFmoG9sT72eXrLteAaBCmO8yUXGH38pugcB
42074ME8P6z1FB8Yl+O7aZheYBnh2AEa8MTsbetN65lPPbo6srLYc4oc9n0/1wFsDXZ7iUMNx+GC
29pF/qPLLxp+A893Il20SGzE4qNgZLHveUP54O/320bsfAr9G+wMWZZQH/wSCzJK92zvw5C+cyyJ
MP16PZUxoJgNSVa76G0Bv/yno4xdrf2rPeWfvjYfqo7wlfUb42T4pZ0Pbly88jiBJ+qxOg9IbexU
04CoWHk7PIGTitTtVQtpDPTSOJyl77vYzjK2nQkCB6XRuGW0ZZl0fGL9n//Ur21Ud2SQLdcJjO11
R9kk2EB8tQarcZzgxz09eTMZ6c+8ogayXhzL7dqshp0fnaM2wxCwg2Zd0dsWwKoL6E0qlkT8Tr24
pJr2zHYUc45pj+Zw/cCTeIB7cdU/C0URMmLuja351YrZeuwIudcVTR2qiG9g36cVKvZFy8UWNTBK
TRNBYDHGFJlfV9HDPpRTAP7d4B1nnQWc5NmQ6LeL9OnY7rpcS8zWT7U/9IQVwvGrSUtYtoCZjlZ0
Li5NltST5o9gk5zojgWOc9dFSuJE7TAqNeGNnWEVTjuB7cSFVTaZQsCxn36AOWjJ9u4vO8yALZIt
U7sur9uTkYzOv5UWe4OtWXlM9Cx1ED0IMdTogDMtmZzMmovk+RktUUpNvChVNdH42za/XttzglA5
0k0ys0+CeZCod4gRzCcHwWObTlshRNpw32QXifxYyameyTTl9Y9tUAo656qV4hx7AJiZjXsOHsyJ
kqXLDdcV11tKM3oiGsZSqiaVKBRihlY/RATm74RMTk5fcpUkGnS5lRqlteHXdHSJ2VmGXHdIc1ef
9X3q8zyTo4yKtl2MdLdASbbilvIV9ekjGLKm2j6CGs++j0dMty/OXuMyDWqAQxLKs/NeFN/+oS7j
+xENoC0jVXLRliyK4Doljq6tHJq8qzQBIAMwbyk8cvsEjnFUkD6Ke3nS0SFOOINLK2HE57Go7enp
jABEKYo66uYyLJ9VYSfa0fXjlNZ/gEYh63aj969FxGiuqKoAoc/4u7NiuTZQ9fYq9cwag9tbt/jq
Ucx7vsVvCdGktn3Zgn6rhcaNgU6Y2UkVSqaR8tpeS54OVrvPJZWHvfPN20YpjmZKq5WdEDTaBKuG
Hnt9CcsSWAmD19CdlDU2tL6uIg7lDMwNNgw43Dr1t8bcR+9rrZLk/sNgBYte/e0r5SI8Y6akAI98
SLjWO6t4nG+hnBFMuA4ZnFmLxNKPF31okezd5w/qVFZLNAix3BomXpq69HY072mVZ34S+5vHLTFk
WMatW6i+O/8Rrynxp7HLfhssbV1KDLtgorWz/Lx1u0u52P+bfSCNQBBpF+O5BpJ7k0uTu7ht6Z3n
swggfvzFepsQQlEKzW2mSUpXeTTt0ZeO22fzqQAvT3+3IxzWL10nBCYD6rveV+apbLhoH7qDdhUa
CSZbm5cwMsZaChQJvgwqOEztEZRKuLQ1XeLCfdBXlQFBeeB4XV2zT9KqCrBCQtgcd8zCEKDloJ4t
ECVEQgoCJpoYsMfC/ZU0QiSiG2ELyuQ5z6BY5VVJ2nkoCKp1p4dxZl2mEkdQ/m1PKisQiWf/izYV
NNaXoU4fVU5Y60gri6j2Mn28LzDhn6qFH0A121D8lv4dxmApjhSkGgt39xXvU8rGfiZYhcUI5ilm
JUIX4Y9I+ftsNvWrqg0QXM61+hT2sHj4QWj9JhftfB4TKdp93YMccb3My4rGJh4XJDR7tjGpHM4p
qzs5Reht/FNbl5asBwga3wDrGoPKfA+JnQd2W0JPPqpdFnkL9dsdxltMegcXJ5QQnAUikKzLfleo
7aUsiY/vc0RFXf6mIB5ZeiXvQZvEiShHBJUEYHQhLcF+u41tj56081I5SWTULiOle2/tyMZrQKD+
N1WNEnlFTrqzP8fuKk0XOo1djMy1rNoSDCNpl723/gWmhw3I6X3dLeeBY1D8/2R9V7iWLlLIXgtP
XdglnbIj/TYEcxqXq/0mTL9BiDIiodpBs6ZDUfRPZFwZB3nEY+scsVWAREO1HalYWycEVFoHl13i
PITlddOXXeG5aNh/RalFKE1lZzzzRrYohYaMQL0Aeop/kWUh2CtOXqOnxBKbd4a8DoCEF280I2Dl
KseTimqhBLlrZoPk0qTT2XEU1dX1QnTG/eVjm1RBdaqMW0s43ktJ/CpFKCJ+e/+OiwCiEIZcfBFC
DfHAPB7YkdpGZ+0ZfAygNa4/UBzSqlQMwid3gcc2mFYY06Evck1Fo1xGlJh29r81i62jv3sI5Ykl
BedYzyrauxD6LiM7WgR5gKQTgdVm/dxFp0hinIVkrMXtjeN7rerunwiHAOPY81Ghrs9mYQ0YN0g9
iLgPvqpcqaaihaopoJDfDS0dm8iDe0FfURUIZTN36JodSOHF+m6F6LLnJlzh4rS6HXTHlXTXMrkO
qCOEqvRNQZfUK6QTG+yjvedgCR+YRZyAc7tTHqLe4Ie0OMxLPAxxI+BiL6htXIA57ADnBmp5TSzb
IK4QhqEeqbYmOUp4sW2NP3loA1SSFHaXmZgXDLncGuJNxln7pLLyNIw1JZGaMoW+CwiGrLgd52uX
HVT8CS+oK90cOu73NraDO+sYbNV92wa6s1b8BF4O5R1TNeFvdPccMkcHuVW6aT3j15DEHuidR+Rp
LWOz6P8RBnzzY3E9zuijvB3/tgqnxI3esIkRCoZnUK3npM5YrtW7zkwyF+mla5VRBYz6tLlrpQQu
TppehiyhAxHsuZonQp+2Hr04h9gC2quAu5r4VvdaIcF6Sv/UNV43bBZbanI6BicrfR3/KPvl/uLg
/d3qucWdzg7jJVcHs9oYujO6Fg/OwGNFISaVzdFq9Vcf5X1ziuyDcMNEBGFSP47VfDqW73Sqhy9L
SrsyzLQMr0p7Boko90aefXodR5mUzTJ3WTp0fGNUtAIyRjz3GvQWL0kVgC6mz50ZkZ7BvyTbysV9
17kU2fuAIaKNqeJdA48ZMEc6CyOu7cKbI6PLLMIw+Fo21JW5d90YODU39vLdFlsrqZQ/9SlRkzWb
Kg/XxsrXkVp5jh9MskOp5JY/v1YDD/KAI+QkezIQjvOVG7nsqvnCUGAQ+savyQg0UqGeDNdx08jE
s0O9rbzDa/2pw/OFXeR4IbzLza5B8IzrCnUdJ9144pcdcIRZmoA/BHt/HyPC90Ej1euB4QMpp+5l
3eGHjET1wp78gqcqqiLiRvr4qUDbRl/qtyrtkaMnNuQfq/zLd40QObe+SvUwCySVMvni7JTzp548
/X6vfnxKiM7k8EsmonAn6XfcO4WFo5Ir9K9ALT/bCqX2OzXd40FCAHJXIdr8feeHf0Np6FdRqjpV
syWuw8bf6kbrgwvtngKLZH8XrEMVZzZcJYRO9LzWQFIKHfcc/3XNg4E4dT+HnVIXSF676QUp55aa
ucNyMy3VHmzihUlfrSw1St7OTZ4RRc1cX6xMrrvr9/9psR0am/avTdtALULZKNtrVGjQn0d8swjQ
4F4O31WwHmD+/q7Yp7mh021yW3GtdXQ0b7weGmLP9fFyMfbVWeV9lJFzgNiWpDSHWzPdOCV4cXoD
Ov4u/HeaL8UHafgMt6OZw+jiDhH8OLRU3l00GweaknxCczA2zLjdtzbkgj9azfFHhSNdHt0MNmQV
pv7QVkQ2lp10isil44Ls+j148WCNFZS/kHjwFzDMWhcpSxglZQFo5gSrWliZsDhMj8I8hwisLI8E
aDBu+GFnyNQHf7ZyYVK1zPY9o5dEF+WlD+xqn10kA6V/3A9WidlUa/Q1ZuzniaPmOpOCWrN06Ioh
P8eVeEe1/+2yg9C/gf2WCx8GEvCYf+s8Mk6uAGP00/046srznzqVl1GPDmoJbOM6vH6Vhy3jNDgy
FBvplZAeVIfdyZKu5axJ/pzYv3NI6X8L/SREJJVhvf7Nhdg1uQwMzNGT8AzcI6sml56igdl/+dGg
lTAE7POVCo7qC6GHIKNa2d5s0k/bhei3MMFg68cyvxsyZ7mDDzSZpneQ5f8pJHc7VQg40BErdRtg
QohdG6uU+RBu9vEMUvSDUn7kZx5gmpuSXmED6w+Hvu5aKOHW9VlBZEeGxoHP7qr3tDEq9+huGjmt
hz5NXGucRdlT6L/7Ej8Cxage93OGiJcYsUf5UGd6115De0iWZdNBN4vkbxPoRHNEDOYvNaGJ1tv2
+AEkuDtghZn3YEzzPzP7KtPxGcaKNxi5mrM+WkQy1CQiRSehlPrq3rLQrJeAqFm+DVzxqXSQzzy4
dbXbQV3BteVv2F8r7PXxnwDOATp6bdTeQJEQ+IUhP9/LFiST5bRZS+hYgjVEtLp8aXwhz+6jPB49
MtU6mVz+FeSzE8hfJNxaT35Cg7Y+e8/ml4TBPudOidgE3Ing7KCOAyeApGVbM/QHeSs2CivjEjcl
plU/DRJA3MNFgN3WnVh8IdfhPqrWqVaZHLh0mOxlSHJ/X1Xoqju00e/5z9ZBth+XYT3R8alXZyVe
pgS0huzXCo+spDN0mgYKJWSUS/2DXCbkkx7QbI8pbr/HSXdc42J8Kvi9ircGRgwccGuHSE09JOXt
QxOst9z/JLyyntVRc8/VU6TGjJYBQFiJ/8swV5wcM+bKI8VqGHW/EQSozkHsLBp9PDWjZz4FkuT3
VAKGXOzaWcGUA7tU67SMtdH+MCNDJhYSOYeS6GET77x0ZM2nQtVZFskVCG5gdtgoW8LqjgY0XOWu
/cuOhZBxktrmNJtPbP/69l5XpzMu6Pum7tHJ8qXbTpEgK3mr2GjF9F5xWyjPlxV8qWRyHTbt9Qav
4QgqdT7Hyzvsf5lqMOWtZZb+LhK9qFfYjJij0F7W7n1/RrRXeBf5HvVMJse1LW7N3gYGWJnRuEQP
gK9pH658T/2e2VDrm8WPaXmr3VjPPusQ2J1CrMTiixhbYLRJwbxelySEQ41A6nP1RLaosQzTNGrz
zPHz7ruUUYqFPyidXPSlFYeCV7DkqciA88e4ZZZl7tBcWIJAmRKNdR0bIgekKHsPVlAsNMxtahKB
5SKTb8u/dNBfxqZNJ5MtLPcNMoq/JnVIRgTcfwq42y7zKw3a/cdsWv4ldZdfRuSCM5GYZW8c0J3p
uSf1uNy0+2cLBTSEhVNSBDU4tis7l9xyb8MinKx48IVl3ETecBW0P0j5cvlGrlmypCKGiqYHHmM7
ZNaoj0roqgu8kw7w+m7NI25QK75X18pP337AiI9uBu+7WWxGrDK/cQitWnKxtT+bjH/JY8pm3h6D
w0hbWmECP6W5EQC5UipD8uDfiRkdyWk0qwe4Vi9kaaTWBxuU/jYRIJ5CfWDv4QFrrppdd4GfjLCs
KTfwHpDdZeAsnbAvfRNecnjWg2etuVjFKRxFNsdI5RwTOXpCd8Wxme4ku2yqPYjft1aKDDq0i4Q4
wzpfMVfQO6orBtV4s/vMQrfq0Lno8bNtfDYgVILDgSCb70HjDOYEe6ympmkkE87b20iUirGMMIeb
1mRuBel89arKRx1x18SLiLyKKUwuiUe5f5bmOH8Ben5CugxseBIhwbaC2IBt/euSy98MqdstWuht
V8yfEvsxOEGligHm0VARNJEy6KxiMdXcm4kzFxxUwwkmGl/XO7EVXC8gyPHz0fvnefX5gAnlZFkZ
0K1MvmAXcps6JPbH36Bm309k34oGwHxVH4hQpOLtVXshhCcbClg7psPVobrmqDbmqo4uckqibUbx
Yp4yw302+JIdmdPJMPy0MFlQZjk/wB13sesLilTH1WuriHOU4/8V8tFZipSaPXrESO6iPtWuBNS0
eeQuchvkjDwgP765LX+vUD0UhYotziR4d/gmoBsh/+eXVGwDjnDcC0OZz8nc/wOMUNuKhmuN3Fu6
jrDUGi1bR26NlAZIGrdHOCgL+mejLolgzNot9CRwuPMkD/LHYVl41EZS7Dm7jTd8W00zFxSqKeh4
FcUxli92YCSZ+c0oXF6cc/D0KFJuN05ooNsRyBLd7XBfbIfRy/AI2OHtKQoaBgi/lmpZsTHDWXYB
73R9H1sZTiTBUoV+TlUoX3lMJSWz7d+NsjtCbn9h/drVOeSiepJPmWPdqXQ9/vohb5R8JdNHyL4S
U1n7zW92LGkDgpX+aOP93b6gGY1xUz0Vym38+sCeo4eRR4u/cDEdg4Y5VAbx42LA/tuIwkUg9n7q
13sao8RxYPvW3sx001KW+Q2mFTwZ74vL2jIdQF+BDuV7i0cq1JI+cSPNDMTXA6EtkF4DhOzAOekk
lK/5ht7twkf/d8TEX8TWJVKPVp6y1dHnTvsXw1Rq/G1IWyo1yTRV2jENbEVIJ3fYQBS1ADESEWdc
F6MfrNWKvwkurMvElbD6lJEV8UiSFbYLq+MheeSZhB9Tgta5nFfLEtOj441BK7/dZqDqsmBTUCau
1/Ukp24DdV+gIIU0WL7xgnA92IE2Z8OZ6HD1aQ4eZgFaHx/dimvlyjnZz0duwr+xulcs6hPnK41T
o8tv3T0ZfwQje8MD7x7vW0Ey5aafFhpOMRa9CwD453jesflBh0ALgU9M01fALdephQHAlwhzfRsY
ZucopDEQHaXY+Kr4H+7hpNkd1XTzyH028p6PAeFZ9EARaKCvachE7GBADjaCK4NrJawJis+GcH3W
qPn2S2DATaUhGxqAq6tnpAYqccuMyBcdAJmSpKk6zF32dr2BpO5/AnF4SJfm/sPQgjbwiasgimA9
sBg8y7vNnH9jQlXcVSdqSCj28vRykRwviShQwIp2FPnnI22bdyFDLxcRh7u7AL9W/B7QV+1lV3hw
+naNyvLPs8EUgRRKIpHggIJYLdEkODiEzYCnPZlPara/cRj4apyFAk/mSDuPFsqbU2qrgQtUNtAg
X2LNOgAJie6BDrMhCoG2A8mxA77zfMNCHoMXfhBMo3Oi/g4tb1rbEo8Mmh/erB5lI1dzcq0DKK8q
WduYuiRtam3oXmasFVQ7FnVv0LCRB0ZdDegUXGR9CSI7NAyomczd8bBmfrk+rWY/dk96xUqzY9aA
jS83NSJEEmNj/IS/3KRdcG74lU91LOTwfYqqdCs9ZUVTT9Nu1HKzzGenKd+4bNcUA4osDOPRVd9v
LSeDoqRu+UvXhGSNRkN/u0umZ6e442nfzmygj9SOI7HgHQznECB+HijbHayKl0gx4AX+QWeR2Aq3
lZb9VuEdQK1x5p8c3vZhw4WgZIQhFcVzM+K8itAFepsfPlQ+/vtdGhZWEnkUF0hM0r4WqzTHEZ3z
Srey4vnWA/X3cuSwcppxdpvMCyY09tU5X+z0YGNwoKqYWpptpL9zsWJIlQTI2Rce+0Iivsghr5qk
Mo0SNlGLmZALMibB0akS2sc9Kk/omXTANvOQtM027VGwpZYKypHakXdNWRE3linlm0Lcc6V5uZSy
cy4zOorIvrVJhoaXBbFptASEoweFH7f1DVqZpJJjyYqoOynsTjo7wtxnl/VgryueuxcNQ7k6n4lS
j6Me6SPajF+huH7O2AV9Js/reKl5BAxzj1784JNPuocrlx79gGYY1njRzuVLgtHOkdAe4lNqPrQO
RK5RMKyHHQY5P+Q8JEzhX6EDNiKDzdnKNkgY3hpk7GnoXKCR9Ia9X3ZZoOR3vrzgLk/cw5f11X76
qXngyfzD+atiHV/0b3+9zEPmBn5w0HFNhYF0Qxd/sK67EIPu+2T+xHHTvRs1gv8zQwBDFwKUakxF
UFUn65aY64vycFOyi9RR3QM9umSph/r5/emhoRCurSuqXdcvrPFP88xk02EqfecyMwE0GmZe9s94
rlUWKd/rwxDv51zPptB3mrrzMLXCsKhHvqcL330H2dA6f8uzGcIWCWYricUhBprg+hJfoLISwXDX
y6qEyO6PL/f3h0RLSFuWVaS+BHYrb1UPA9dpmHENpAIj9LZhxDiUlgg3/NDjBQuaFiWKYNwDncOG
TDHYZCWHiLOGkxV17XQiIyEup/M79Puo0Ek+MrVeo2MdSaAmEblTVVK9HgpLM22KzMwnwuKjOxZh
y+A3/+lr1FVuGHjgtubpvQcDk+04fvwPKqObVKBNEu+644L0ulZDGlRyalUzHXrUJ/bWMAUhmgaD
lnsupgy63MkAzQ/mp39/pQHnOX224yDVfgR1dB3YpRg/Voet368XCuyic7YUnHsyupmfiz7ZTteW
jW7vYi9AMHqThVNlouRABo83O+GjC/+RCbkYPGyxiXgfaQV7TwkudJBpvnmKF6YmHf77V6sjG/wZ
0akOFRyDVVd9wZ+IFCNnjeNmKIMbLBPyUmTUS4di5BtNCepjKCbyBcKAfjlezp4iEHepl+QshM+k
cf7EmqYPQUtI19OR+ARjCXqSkRfhRqDdKnvzsiUGzFoaxjCcKP+poc+X9M4DXnFzuBXgmLdNluhs
ZTpzB5iJ7LOHnW28z+jXyFB8D5a4wJAhheBFFpgfe5fK4ECfLdrW7/l2ufPXW8lf0dx+G2Doo6+7
l1ZsvnuPnym89Lf0rGFuJXFHlkby4t73AVDLT4xK6urEkqipaYaBwFrch3m/e9nfEbAckUat1+q+
a77X3NuattCPn+JiJ/26Wd3rCjEALeismhGq6l5IbD98fMAlQ95veZvX1zSgt/CHEHAT8xSzkyJk
0JKUXQsZGYOrppkxE81STlqFpGm1UcyrjlJ74Bnkab4ven1PFHXboFG0/2+fMlsBpRVeVrjiDCrE
wKeua4pJqAd79yx5+U85SXfjhUdY6XCI3uK1dnJU2o6JkrlR03pL3eo8y63xoFaOY2NbL0I3uvKu
2PXPaOTIwDPasxtw1srZoy7YYp39/+cPQW7VmQGMKl5giRgy1U4dvJsWubSiO3Tglt80rSR6pyYp
sa2D+LF2A7DtYEUY+yXyQ19kLUXyDtzQzGkWQ/dGW2RXZwiMtTyLOdfFMVtyFqzz/A3EQw4a9f7/
3H8aTwcUEK0nMPHK4TQRzaNQNIJNheEcOQR9tMU7QTcAuvv7aMdvNxCQUT36kfhgTcxS3jAj22gT
/BJrjtSNzCqEm6H+/Hkn+77d3LG8VL9Xf9HFttHUP8QA2XSIUqaIAosLIztqVB5t9Rw6jCg2rgkJ
1fklgzyPXPhM59vvLZ83RUhx4bRnQpyRBb8IUFPiKp/xxSz8clEmHDrD/A97fVIDcg7hCzK9KuX3
DReN8oqaFNaCFnP8GIq8BJeyX2jyRhQIXCPGnRE8o+t2TkcCUTitD6LvSNUrYxFhJxITk4Nx3C33
sr7JMWGsTsctmfDDV6NulGC8/Ypi11QjbpOdJF4OCnpyJbRDQdSgNHUddU8gWWQ8/Y6+0CAZ+vkm
ToGFjlq0tsT4RDxqGFNQYFm2aOSiQba2ddkWzSsriv5r66oOtHKBOT+YE7voRyT8DCjt0XLNPw5P
V9/ie6bEIg4X4lxVxv/OpZwTaCzCWeQIQ6VoLcQX030+bExrzjnkksYj0AdCXC6wA8VqDtMisW0v
m0UAaQRPjd6EYXFawxv7Zg53rOLp6h08333EC9RuCX6Jxcm99QL1Ysqh9UWMwgYAyTbutF/7MPaK
nfWVfaXcGBO1f0Y0Ht3+hyDsd+NOXxD7Z7lr49SRbixoEBVELK/4t51OkOHXJ8CPJyYsxAmSz23b
B9sFI6zbB4GK3WELs9+k2SEkpys+h4EJKDY1DfFsYTI4CziATjbMROHmEsw2GI1dDK5Z9p6ht1nf
0xKSCVzYlcxHd//B8nN81LsV+aeU50s2TrKXKNyyAcaT04fkBf3N8LC5Qn83chuWeNk96tNH6jGG
JJd9Sa8zyC5z30JDhPX2KkbUmimpIG3RP9orHvIg6osePs4J5tzBYHh7x9rUEwK8idwpQYg2rkI4
1FxFhSq2ciQsBZEpARtl76Zs8AmXmi3/i+jMNgHVplqEDo9FdDrASRbNk4V7kvcQdriVi/juhG08
4HM1x0dFO4BUI8Aa/+G1rbPqTVLJ/0fU+EyRUk1O7nQjg4OSBog6pgByx1H8VDc3qivvdiIHnnzy
nzZgS0Z6zNQYxUDT24pAx5+oYCZHbmPdm8/AA7PmVs542JTul3HydzMW9sS6k78C27Lcwx7ioDWh
wn1HYRegRrCDXd/rwTyJno6vgK4mT+2CxbMj0R9nD9B5J23WpMDVuDjYsrHvMKWCmAC0+j5sRLtJ
HmkcY6Key+NMC3r9hG9SabqMDs52xzCgO5FmVR45UWKyOD/w4auzSQ20vXt/gLUp6Dr0tRRZuS4g
ihiH/t0XKNLKBtAmWCEyI/QhzyhfekxRJl5PGTfM/kpU/KMtz1jIeYPTCPqWWHXp3clASzyQCpSz
GYgaku20c5q/F8xBOxufaZetc7m+oL/XD/kr2JS05qor7HdmmZ549YRSSTVYKLQyY+NOh8yhJxGl
D6F/y2G6Sj54RDe2xa+E+kd41h0+ZIRk4GyZPKB4ly384aW/8km6uTx/FpYbRhTSEBJU+HaFlJzh
J/VWgHuBNh7b13txZ1EswLUiwSpelJ8agjHtkWajGRk24NKou6CgjhJWgELJKAIzRmnBb+nskgIe
hDR0CDxYCNI8AZX1qMOaBAXiQy5zjR3gJddnJqrdG5JC55h/Wqoj0mDFQ8scQVkDEQBgmvUjnMou
ip4YZ9OU/rcT8knJ2OPpkUmR0NSZT41cW0OmheQ7uvCSGcnY9O8ElzgNgraBy6o5rtC+/hSp/8ia
/KTeeunZliN0eWGETP3Pb1WDJSZ0MCtkM0zdoq0OV72WOMq+3KvAze/7xrW7HBQVjOhYHtusAzC8
VQB0ciI9mMaewuou0mdXM2BGB26Xmw8lIrFoft1WFAJSH68DjgSEGWImGr8YtoTs+YVqOSIRvygJ
iDQVVSdi5w6By5rY1v/Y4Rnl7A3CZ1nVCjo7Ie+OnXX9rvTXeUF2GENSJK+mdAPCdBpKNvMYRsR0
n6mdTnlWVj0BQIgyFZAOhoYjgvd5UFQPbIa3fCKukDmoF7R3Y0popNoLxuOTTDjj3CMMVKQ3NA3A
rE8kgOXya53KTq+WTXBhcq+F6SNt3OW3sNzz8367zdNwViCOFO50AUVzPT07zjVr4C1KLVxHwfJE
je4T+rN04LNsfzyE6EbKrV4W2ejBWHwTryEtJU3T7Otl+j0ydPCwS7GHrmnri5k6TPov2Xg3uZMd
nTxx+AtZWDobDYDT8aSH/wSXbPdRwIl6EiyGBWFSnNxE1/z+8hSQKyiXV0iroFyJ1q6+lU/Re30c
HD8JV//ohvCI5OlUsJNLRp2vr7QuUjerqeO9fov7nYXSRYdnEZVstf7P+jQ9b84VC2HsMINnqZVX
x6r/93F9gh0CejYDxVZdLfd7bTKpN7yLXwlZG/RQ8BY+d5T/EOmtE9rWj6RK3cs6wUbxdxKyEKWc
wbFagqzPEq2CneDC2FCeoMeXfLj5fPunPkR403ewEDgWaUFvxCB3sn2ptOASP7CzwNkDGpb8ntOg
l2DgkesOj4bZEIFyUhnvtg/L4ZHXQwtkqZ5FUIaeTLe0bdkHSzuMvt12c8Ay44m44ldySo8y7dLP
1J/zww7FHw/ZZ7O5aMgFEBM8NIMiXLFKMhYAiKwlzY9fzcPleZUNA1r1P2+SEtynp1MWnYofEiFH
0qiUNGeqK2YkHjy6QnJJWJZZTQd2PhAxZZo3vUP21Cku4PlSvvY/3C3wkim7AWbOsGlbjLjc8281
j6837w7d1EtaPcn/cA3HymuGmIfnFr76pRaU2PptUHRu3bJ6avU7Mh0zskPl74tJl/UGjetPgd18
Dc0oRI3gWLroTvC04UM05NCRnLZaZrtMx8mX7tLwUoRafJ1M9RfIAdQw7AavLKSq2jcdQP3+7b88
QWXnfjQrlgkVC8AcXCBqZmk5XoVPppmafGvxFQAb0PC98JsMGgBVuvv/gbrz9DVrMINbrpkHv6GG
RLpPJAhBtCG1SNG+tM7m0LyxSugdn2A9B5j2k5itwBwUbQoK61Z/prZXz3xOGWKec4oViV0trC97
kR4AliXzzKK0f70ueycT8VzOGg7/UgcbShkiTJJszCSrygtSUdzKbZ81RmouBxQrIpKigOeS4t17
1uGMJaF2hqo1ntjoR3rQ2aNcSFijjbADdQjLWI6eDa2s6njz03OvXJKvplVPthKA2rgyw8DL5UCV
kInjc3ui5OuMDrpdX0UciDkmoI6iLbI/dqDQXMWJG3AgZhy/SeydLBianU5vUS8ioLkXNAAXMJ7J
9zc4/SSHRKiJNHfJNmfDIn9Az6oyQmyBzRGOx1PIk/ic+Hqw9pFJtorpd8RRGnse04IubB5I4Hxc
PyUByd7R71ENGefCz9GMtjGkYv1G6/qsk83KbRDLDlHyRVFqBt/0lkyGskSe8/GNBSaFhzE4SMBX
YdwAW9SExSfPAqygAwjk8D3veFBae4q6En0SkdtOJFceons16VDQaHWPfeGb1YeDBVNKB9aI9TNB
3XcoLyB+ixsNWTh1HfXTe7Og/RjOgO07T6uZqkAsmBX1GS9LbRx6bMtj8aEGGuiTttTyCbDWz2tJ
2pAeL4C8bGJy3LtngV5SsCmjz+8DeUqueLYo3/h5baJX4yz6fWYb5fpE1e6Gg5pISaQ6sMeMAvnA
NdvHr6sPugKrd8jJ4yPO3ACfWPHkPBCXVEAIRR/zC56iYDiWlU9Nzs/KDq0BLkneiGN6F5+DTHq5
4nEQYSc2wdOMSsy+ibukhN4togBtSXyanUknZkbtWoOwjrHiGY8kmqfejsW5Gbo/pMiXytcBGDmA
KY7YU1VGxPQFE1zZ7c+KlLOqHsu4w+I4Ssh0Cyxd+5A3QOVvDCADYLQBI3HKrcGy9MXfiG8nxVIp
VjAg0N0qnjfoiQO5P4b/U585OP4Gaabh3eW1HZmGOcfxPRFIUtvkLlsRh5iilmdLgg7F75vSBlEQ
grBqb1ts1rVXmc5jnnygeH+9wIqQffEDMXcdgiX/Jym6KrY+WEAbu1My5rnraEz7hzqwkau6fI5L
x/8scJdL4UDGZgoldiCplQwp9NL0DeJaadwOPCOb6BUOL0snDSGYPRR2WgLHvUClYNDRPr7AvDc9
Kavqx43FY9f5czapuKooEhpFtInwE9b8TcbExnQJua54tqWN/1KAD5MLCaWJVYKQtycb8CFxC9i0
UD4R06axDy3v9VwHLBYzbCmpnPxJdro8akgQkihRjq2HIxeT65xaXe/VP9AXYh22m9Ztf+rF7Bl/
Pn+y84LuWNsK+3jq1AhoMnxucSJL/Ix1X+BJUi/axumiBxE89WswwZhOgdLLsvLyOH7gL2zS6OSI
fQK8SEQIZ/5mzFjH3BdOKnFrCWie/xPGlqy7yUo33LqP6ETwu7lWxpzJCEPiAVeEklW/6rStK9IA
CEwfwusRuMx484lozqIiWtvpsVxZR5TIaP14gGWloi2WjiPTfHaW2asPEgAX/cnGXq+6BzIrwCVA
emSiCB79IhybESs6r2XalMqyNuHDUMI6OuzBqu/03fUyHNrRCFCKS7QvHEs+byrBUkiNyt68XrAN
rH6rEyRn6nzD/KAxjOy5p3v7jcsNWzadaEKHKErTICItvTYZIwvADNiTLgOFmJ+Wncd9qaRW6ncY
8cp2A7LjsW5Cwk6ZVh49IsaDDhMrBzyosdIvwSCLQ8p6O3948e4ZhtBEweM2tMZENz9TyPqgBCeS
WgXLNE+SSmD+EXHP9B3+1gRGp8mDdNrwLeyTZE/JPITd/tOTxi+JrR2VdQJZoswCadleWxhndQv9
UgVAVtvhj1BBAkcIzsHqmPs2c2I8pXvut9euw/7NgfawGSJ0dTv+Op+v1oWirrvuqeGjNTH2vthS
Za6NsRfvrWbq14+wFOK7TIsLPAoIga7WGsFTANWt7LyfF6ggUD0KS22Wsjq6sw1XBZJ+gGXEX31h
nI+MfwBYq+BUSXHt37GRPl2JB/tdLHK5Rz1mcAumYO4AzJkkT3VYZspfCqE1dxCdnFPoA6h0FO/t
who8mKGsBlC7zFH4qtmMXrpcpt9KBi1qkLyGN1MXxvVqtUCnfNDz63ilXnZH1oDRmMgSSyT0v/fs
Y9Rhwxhjj6uIShB2nYFQ3RPJoH85kZHtFiLzoUlusTCEmiuID7dFCNxnBtHOIVR0Bh3omiXUedSF
9TXVh7HLrpNEVCkAcJtYGJj6qgcz4LfHzMKGzBFiz1CxCv6aI6+G/LqPMk4SoVzPyCaAoaTQMrB+
fFm6VigVs6HqvQ5xVegRSlAMsbjy0P2mdSKzMLDFQ5gxFJYhDxb1fyc3ElY/3Lhl7gpRKogK1ThM
0DU4IXEmEp4ZiOBCu+3I4QnGltsjgBLvnkSU2Bn+N4KHL9nWdvFkk2y2gjXxQX1bcoMu+ep+JHtn
pMesEEr+LlxivCISc3VMteAzYvVmn0bYbWRhpca9qY4wsOYRxV4WuHK7qI89JDo8vvfwXEdwPCey
FDwIBLync46tobBU/H5BcBQ7apKczRYtqK+lAws724P9JB05U3BKn0QgQ6+izEYSZDXaEVqDbRV6
u90kcbCPvXa5iY0fr0B3VtjYgn+VxRvm1PpCjvfGVZZNK5mhZpw7IE/raYIkvcW4njdS0cATdJxY
gB3OANuDRuHtomy3RpF7KWdcxA0S7jyMXUiSzEdERLQgnDqa/6CknaBZUyv/cp8bdPIKYbkH1fCL
qS/2FNFjfElKRUiDZnThuBM/rQAo5jqbOJp600Bzz1FegXwj7fgPv0s+FIcDQQDtlCoDNCBk4oLQ
xTS+oXKhE3IuZDTVQWKFSQQR14cvBd1uCjaJv28g/zmPt7JdIVE7i041Vzk4W9JbddCWOZ0rFXWc
qlgxNGBDRLSlpetuiQXZgVjuTJ1aNBHRT2TFXQ7w37TmPAN+9ZjYDT0yXHI3LzYCw9wMvpuM6Y+G
JkEgRsd9kIfPNhMR8kJs4lKDUCk39AQb9mqMTeSLUvbEVYfsOMOjF1ksXidhHGE7fKD6ay+OKHCE
2EhiTgWP/V3nHgxln1KvP7/PJv1O3cwl0D1AveJQ3vHw2CE4Gss1jct+X35NFC9SUTJ5P3YhgUxz
nJGK4mV9iZdKEA/JYejJQnGWwVMiP+Ak7W+jKXuxVGzWZCkjc6hGvbaXVAiHQrpQV7AsHVwX6FrB
YVzNkNqcNQGbGgYhTrmVNFdWAAIx45fKANJw5O5mrB3RzsQez+mqAfb1+2IFpXHpLyuP3AVWBRIK
qEavVRs4jwHEdmRJNO4L09JXdqgNyCxgtI5cxbmSdCew43zbCe+2eBFQSvhS1SxeIZj3lRPmN6f2
0BXVO/Hv2HINb0LOE9yMXYKYrb9N/AwGXSsT33yh7ncnafyyAwp0EpKIPiKeBpCIUN9hUH6awX6H
SokvhZieYiGrIoExiDr27VUsmuK6h5uj8j1s8PyuMTVvXRRtUJS/Bs+vZdJeRkKzCfUXmxWQWFu1
tJzDx85Acq3gq9e8x0+TI2AHXsiuYP792gvKaPc8QHXbP6ggj6YobFUqGMKZ6NE3m9AiRADdCx6M
jPtn4ng469c4JW8AvvIGT+Y1WzSjSJfbh9WSgPsOfVy3KtW7isLBXdJnhVI6fu0UROWSXHdYFHEl
o/IC3mlwSD/af1ohsqg1KpCJvCftbJ9XxmH7gF68FTHIx31/qxSDGG4WW4iFqNqs+eL6DCxE7GCy
n+02dz+oJVy3zFxlYioZdsR7s2AxHyNgihya5xsx9haK4hyVG5j3nJZo7Ucf5x4QxVk8sCzyFKSN
61Tx8mm2ZnZqVP0N58HyjftzQpe0RLJid4IduKklwAsnd6v3g+jfPA97d181XMtW7pJwganrufQp
BGHOz/ognNxsf6zfAjisp8j2xmqT++KUQ0YDIloFTipGSZfJ61IEigyRfWoMvPWcrrF4bdmy9745
oHqVP5m7Yr9uic5t943o2uajs9NHNuChOaL5v/edCjcOLe00a+/qJa0OcbaULVGnjTIFOnJMYBVm
bShwNoLwMUP22XdOOGoKHdGiBGTX/X1YN5wOFXwM/saBB9gu5Ut3exS0mC9ddYtnvCyiVadPHOzI
0nE5Oaakln8CqaR4hDgzrbD3s5/nKeVLH8m4PeIa8ByPg/e+xQqRN1fRNaIVPBxd9GqCjB98SEBc
wZO1wTs9q7MTgyhFn/dGrg1hWw8UnNnrDfKXERBa4jvtiic02gyU55xd3b0v1sncJY5tHd5yLfFq
iyl0IaZRFRr9oJxX20l3dxNMWUMsH3dmUuTzpgnnXv34K9oTKUoyp8GXuu0x67jgI3a+KhUmQ2oT
mPpsRLeBK9escydl1k5CActxJNQtj61eQCBo5y1tip9l+jBS70B+O7B9rCfHzTA4z/S3xcLB/iiz
vT1x2eMDhbkpd0RvIVugIMMbKRQBxKZntSkw1GY/86tH2Z56OFabw6c5ln0lhY0ml49ReFYZcfnL
xVrcErt2w+TxRH1u3YPKV+bIDjjJLATDh79mb/GGPVG7aAyH+fxO6EzMRqSevHILhsxq/bzjkJ3p
15JouEu3Y+sWKDGLPq5VlaoDCE+nj2NGhlgDm/x3uJtk5OM2BTX8N12w2MUr3eopT8cpXZCaWBzm
F1W2UEIagRIxVKzd/eOPX7OgPFvjjkqDVzxlaDgdlk5qBDNL6uXcbzR6M0d264m+2DjsNyKJlpSd
pGGa1XarYDDUaqmF7+cbuB+01wwdKRmE6WTmLyVYi6JECeG6O3jR2tewCOUA+ci2LFwvUbeHk2wC
/uB8LdPUO6LX/6ebdfFDREAoHyBYSC+FiWdX0otkL5+bszCdL15uL4TfRyrMf7C69QQa2VGDSD8x
Ozsny7Sk4LmaaJiQqrRpuG1ltCu8m/txmfZM/MDBgymiGcgXtggbE1FROAYf5srW/sC5Z4xmAt4S
75KL4IBjCpOK9aqAJjOvYHlCNPvPq0an8YLGnzGcQPZ2qgCbLKprqIAsai3LZC6k5Uy+vOgnpZfR
ENFcepOhVJd2JFDyZqaNzFN2wiq9o2QSRLGY8oKedjBd1bx4jIKBBOHejgbTJQYAfrJ3qTo9V+M2
xHtXpm3X4KlfRo2JGkqARpvMdaA4Ap110VO2K2MBlaWqHhfnr84CU315bG9jFe5byAKpwBuNeBJc
RTEYatIWcOQsfVK9/cKEw7rCY07NCa7hpA0fa+NhU8rE1R6yD689Eb6KXyzqPLe8yuntlybnnF5k
d2X8oyYFnZONnqFSDIXO+NCCPOwT6C3ldbxuUAefoUvITixqy0xgE1c9pBhaH8meU08hURxjLXTE
moMNSTn9pFGSMNPqCyDM8zDVO7OIODeFj0UOx90itFYbPY3jh/QHu5V+X0SHRTYCyeFj+8Wf6l6F
OpkuFCVzdWcX+5fFddc8lMEU0n7p/xpBug7mjxhAep2GI7DSucOkrJGrQEI01Y/IrmF+8gDAO3Pp
B2ngQLq929oyG1pN3POD7wHCXguj0i5fmZ2Kug3vjwBlJzcmlDROUqOUGK4G6y0ft+Ewe4nMk37S
OmSuCiSxfQ412X9U75ZtVoVSnnsFrhcIi2TonERue9z0Vwa1PrJhM45ShB39rWm5Pba0AeZekJ8l
yWCZVlbLCAyVLoXG7B7MQjg/afv1HvNerCNryUs9V4zW2Ukp+OJM1qRzb+XhZKaQqKMLJdjVM25r
/id3CPIWGOH3YigSxB0jMFaOU0kTXPzHlBDeY5WCPpYbMzeDd7dikGl+A8fsjIVLmxpjpPySOgKh
NN0NB0QckSmEherA2HqTTBsEM2BlEU5UQyEKVX6X7BC7+E1z0J/J+hyW4pDVapvQpBGL4EE92DCD
EuazSXB5ypHKx1Q/hWuDbzN12qDmp85VLe2L1WiJHzntAyaIe6vzFAfRTEy3AHJFIKgtyrJF14MY
Z8qHmLUu+PaUUhm1VwwXeIXB5dgjirVivh9SlRvSgHgN36OKtaXDfSrGJlOWPvjALAy6bBEK0dq/
GDCcJmP58ODXDMyGYBCpT4/Dc5nmZpJ52P0I/mJyeL69u4WZIxxYOHEREwtccQry3AMo5O9AON+d
zoCfiW8WI7HM94yLhnOvYrUDgmcCz9VYE1eLCoh1IM+9jRZ0HQxyAnXxlrfAQLsRo7EPlsiZvjhz
6XBodgGG00ogGqjJnh0WzIj/MSPo90Apky3g4fY+VKg3I8qR5795sBsYcYvLgzx983EHEJY2lYfx
SvuiXoGZTkqqPgOFAQv3uql6RvmyzMj2JZZRNV9g+Xmwp56zn87N0m/xeencrTsiXNzzwv4bm83t
hsGRKUKzmi/LhGOQKU7ap/INzLY8eN/IbrbRAzkvwz1kb2U1xbA350t6zHPBxt5fEIh7FH/jMp4Q
K1wllXtPiKiUZsLy/xDhgXuwdiQoMRtWAIbevLNPe21o1SUjCZwsTnkEbK1DsN46Rbvs4jtTaEys
JCvrK7LRNnCdMzms1rWKWAlllDPiIYhaYaTmJyUAyRtQ5gYRLpgUMIRCTLvkWimbrOryN03n6hVO
UzHLs1WtHcP/d/8L5Po2meXZReIZ9mt7+uP+/ML/HKplnxVcjtdM+KGHOEPfBzPtQdpeNc27SPym
e/z2GDSAnj/8tnqHgSy2T8WCAzDeUOwgQ58piIjheAskBZxL2w4anDX9EX0894D3uu703MwLwFEc
V94WIAybGhf8ICCePvMiIIgSudhaH4Q5eQQJolcxOKXGkNCnKiQjEAWsf1jIzeT5EdlYAoXNizZ/
3rxBktOD/U2BOmdUOkfICYHMgEKuvqmY2oTjBWdUcCaczvEvlK7OCvYLrwAc50bjqJCdBy9U3f+0
54nTyPb4O+A8e7aln3wHzsI/lvExlao6YcNrwO3PGuR4pWaOFxfN7O40ImwgsGJ9emjkYAPlD8UJ
oxwF9JeLnip1SO7n896iIp0l1Ixu+8XY5wr835CPqemSGsZeYQNj5+NtpTOpR43Pw49RDDAtezEr
AbL1SSuyJi6XEwmuIqYUGfjYOW+4rODRa+sEZNDc3wLdfXK6rgO/jzOrjmpA221sc3Gnfd7Ev5Ep
QH4VIpf4umeEP323VXh/zkypfdmusoCr0FFTGjFAbsLwtn4RYpkwbF29QQfh4myUkq8l61CGm6b0
J9KTwFiJPAaz02aCTLU/mC3J8J0A8stG7dn1Mb1Uj7O3TRm4g+H287AoEfOyB10yvR8HRErevfdB
oYv1jN6+f9bAFQ5hqblOkSskgBRbXDJc9FXYrIPw/aWubaXehsagE1HzVmu6rW711PFvgSdBAsn7
y9XkVFkdxskwkeSmTXPXiWiSKMnyr2R85IvsNktvJnCpu/EGHQ0gBPlpe2YfYpE+DqApkvK11stP
5P2Rl+jvG+swpxh7YV8gUKuk2AWLXBbnrA4Na7zuoxOiJUEtufV2Cam9TMakiXBJdIax+VXBpRb4
4MXya5IuIA3mnjJy468fp0u7QZLXI4I3t0ZDWZDhQXpm8S6jt8W+eyoO6c6KkJsUf4QFMdFHz+id
LmgEKlW/NEV7wl6sF0605/mSovG4Su+OEUp/3iIQIqzamKgXGsOWVq/ngnTzGMiNShMsGW26mtF1
GbViFG9CKOcSjSq15H65WJE1x8k7/xZ/hkdmbdlVrXaJzVQJDkpaD1xJ/avJiSRkrbQATj4FVZWQ
Ew3RKevWBZhq5IRc99f2JCX7apfM9qUAqrevmqADEg2M0WJXCGXKoVIQ21giRNiOmUHRR47H3CZW
Tj8hiWgdkgnj9TnsYLZ+k492dbY5NE8cWeMe+7GNePt5lKvfEaZ0EQFMJpEebqpPOfazlw4bcEk0
WZsk+UEh7tye0h/UuHsTr/JzF73idlc2OkE0AOfdzveVKe0qhnu88m8vW3eRbBV0d0HIdorQlhax
y7fb0hXuPB6EPid3NgOU3iDWIC/Bs5ysw/GTPpN2IVopTJ+HGqXDthu58BI9d4eUgXup9DoAC5v2
FPabpWWwkm9WPR4xr1E1BwvUXe605nhmKCXgCoSjvA9oB8q0OeO8vLAuuk6VRIjaYJDMWboCD4Up
J1SgZyz+15gJdvkWk2zKfAVwFraPgQmJ3xN/17PoVaR+8pTFGkF6zR0B8zoL13rLaghbfuOej2fe
9IRrlnaStHZevuX9qFNNcFlcKQlXVsxURR5FdiMjN86bejDduQQ26J/NNmXQyN5tdU95MAStqGp0
E7dAiD109vnbtOhcE7BI8iiwYbOxYs/E968cclih7OVN2GfszFNCji3iWf3RxKtyXd/Fxj/dw+RK
X/DxhKHI9I4VimLcEiC3BeCdOdQYOxwlIOUo/g1oLzl/HJS20pOwc02L2qMpJh2DQNxVj53C6YqF
xbVazOrxFkTdprFaG3/Zun2MkfKgJExjpv144Hlxtrb13ycjzUNInNAcFGEoTEliTMeCsIQJsVzq
NhsdaVarDWFj+lwqtJMpsx/E+41EYocJE3cSHy1d6ABb4VmAxIK8eIy9SpU+n9VC06d5m3eUuCGa
7UwIXnIWu63e6EhcG4d/lyqdsFQVRD66GShoK955y+g0HjnHX/ds+MqgFpIi+Uxg28rJlZDUPq+y
3r0CEcXu4cCkATcv6Ix1rC1BJPoLk5Ev30qBhuis3LwzTH5R0JcySGjTRKm2698MvaxXIBSKVLPt
0hkLSilFWwBm89uo5X+ph7NQGTGKssz5Ncp/qlA4kd604i/Ps/ELDgvssB8MM0gk13MyZFFAxh9R
zXHD8xfVyDqmamVElLNQMk15a9i/0cRVjofvpVvnbCjNaowIffOjLvW883ivlo3QhF+rT5rFAeKK
M8j1bahZKMn65mEO+4z/1zuoM3kS9DaQ4dkOJdEboqgW20YLK3IttIb+GB46acOKdFAFGUYWu8Sp
GXAveupEkuxfILXa9R4Fxh42koH2UROXpJKr1elKa2T/ZpDrybQQw5MKOAhdsKDeX8CDZYGFRcqg
k44m0JPZToAES0fbbha8md5Yj3nxanxbUURqwPE66tlsSKxPDsPDGJa6b0sotpFXBbMxd68fUbWx
NTQY2Fx4PM6w5E4WFLh7eilBOTIDqZDGifqHj19q/WQ1gc0p2HfUBoPBzLBBkTqzcGuLuPrvY2Qc
snopIL02c/TAfF5aurGvdYKR4xNkHhf62+9e2jvZmSzEa2as3kqEFbgoGD9TySkSQjiKpfNQMBl+
pcsGSlkJy5edJkSqgs8lee1Pq8vAZR+tj02lgpv0Wyety0g/qTnVo0vP6IZZuuSSzrgf0Md12zPE
oNwGwXvGcPOmiEaKqSF1ku1/ooG71/K0Oxm3ZMstcwIbO/ZgZWagG6CzmAgc+F9LMAzyVPisdxsw
VHUG/ECSC84K7onrqeUd6SS7unJKex+rLvEkJOE6px5SNkJaPT3RbMJzmx2X9XNaLRwkscRhdPtD
0eUOqi1AAiE6GIBIeGSFy+8ipk4O8vNgknfIWQfXgQbyZNdpHPA33MWThJdEsa6UBoVy4bZyDo5e
KEMK2NFhcwuk6nMi1gh10iIn1joNgRILyheWJxU0O0GHsfLiynLJJ4sy2f2g3LLxYikOQO6Zwy6L
MMN161sRKORfkpe5m/OlJQyEgUdnvRxN4PuHJfzQgP2e3OMlcwsBu0Y0Um6UEaHx/oPluW/HggRs
YUpfhogzeYH2cDcg0YLl5g838uTDZZccoahS5SNneQbXGP5PRuy5789bTZ4YCBC9cPvB2IqXJbXc
drvGRxOuu0fkKxhVRGMWDZcbHw/TqBFKgpfqg/LKhjVfNqMm5K46GFiUHee0gDE1uUg32Zav21jG
HMN2zTTf0K2I82Cp8b7WeHui1iIrsi/pLCbNb2bhlcsCHPadN8vy15jdunmfKLb5xr0a/4OMprwz
lK58nQBynWF3lK0YT0EbsEw/7+TBfG1NLPz1tpcYhXPUkcWy/4stjM+39prZBKQ5f486a/nFgpAr
WFjnL8HZPIpXTZgIFy3zPpXx7HalAuxrr1hTlYBag1vviwdzupGTk2oQMH6onYEOqdILwOMWEI0I
dDHKeSGHhcMeDoYKiIcglqDwgkFsQs/8AeEKBV9B1AdN9wXx9VVH2fgRsn8wU5iJLYZDy3gMsBLg
va7vxKcmOE0yKqpPdjHSBmFcVAOtyWuh6GFSgYsAM3RChSebKiB0BlW3MOVq1GS6gqLTYwftczGN
EfibQ8pGMbhFz1BK1HW0VspYExM4ZUWRgHZz8Wmhw3/nS0ug65dgC/Jo4LAlBYWTjroNHrbjH+Cl
ewFpzXjadcChjxltiaSKtG8tkExH3dGdh7K7eYFDVAUTnPS3nQCHWgoWDAl79KnnP0aPMd4S0URW
3SGmPcLqvXfWBBVHKaj2sX+ACAN48UMUUxfnvScU9nDovWKtNSkqFbXXaT9k3Kj+4BNE7DchH2IN
jn6QDcg4OQQtWxp6nskjEsVgQut7AriqUk2Jc++kZiq982rkVlz0MCquNVUJnJIA2QLHI0Q8UE8Y
QVd+fTa0hoIyioG2vXYmVToHeoqZ3fk88yCiLncL75rY3rJbOgDDNQx5LL4A1uwFZsjJgqYX6dxm
C2dfK3X9XqylSVkj3MA/tSBgOJiLTLX/3yYBlT4ecxMGYwDIIwPq0kwblyNf2e2pF+kJ1fpBoK5P
ltWPJ9f9lFcXBiH+uMWAuKXMjfvcg78tA11AFeQFeh3it8AUzoQio9OwmItyDCqd/0f+d1NqaLS7
+xDsS11aEnzPbE4C5eZnaBAZjbpj1f/V8qrVn/AeXOIKQ/kgWdb1gLL4HSa5yk5qeKCDZ+Fu57JF
+Wotuwde5W1qk6aseP0VkJ01i3aTP2seU0iw2A/U4P9Hbz9S3mEfDjIu6ayrB6UxTk9eWMk/iCX1
KnI4R4+BeuKUYOtNB2OzT3E4qMQZlhcvD7iLvZ7DjCMcgFsyAzm1yz6cl0SIBrjRvPDcYqYnwu60
TqGJ+lCF5ouFVgB4gCuSaHDtfGWjoyP0recXmj8tCl0zl8HUxl96Fmfkoke772ckD7rtW3BHqkY1
yeRUngbjHnnMaLXTp15tzfSYYePtlSxTZe2HTVQ9zqzgMGHJTvvzX18M3q3DOLXcel5ijHWImNye
4mCymbg65dcd98EL2okxu7E4XXrPC7lXUcmRSdYs4Mvtzb5t8oos8OyZNphQcEXv71Fbkw6cOHNe
97izPqPwQom56vuHorslUIy2hXsPGM6H2zn3OtPOFiYTFPY/hcZsnvFZzZUEDBlE2Qj9k1o1F19c
6aDRcTxnabSJw2brv8HGTlT63SkdrfVCi5KlbZz9eIyaEXqRqfz874YlTV3uzi+ib/ftcdXZ0OF+
ungrOdzoZxUHoOiopnJawZhz0bFxzX+iyKNUyXVtm7EEZ/x2pqSHiw2Avb67Mh4Ro8c9jaB84KPn
86qwl2vwc6Jscjci7R0yrJUqV/vZkXaoWW3XY2QXNBgq9VvtKX9lGm51V/ztKe61kIsvEHqVyIlq
3YXVcE+JYtVUeLBGkG8kNtg/kiCWt3fP/UmrtV4j2Tw2qEn34n+45RPKI18BvB5pzJZBij2kaHpd
GGpTj63RAOxpDps/wx6KRm6kTtR16fzqAzQFCfU8MCyrS9N9NLF9/k1sxIJQdZ7dqvNPAbDXALa/
ywRpKnA9POGEVwj8DCD31ph1zlFH37URciwFkoM/NTes/rqnvJsGQlBcuYtVtdxg9CBACqXFbu5K
8K7Ajvxf3ez0VbblVbmjl7hbdf5WOsw0SHr0gr8Ab0mUKhfyQp2Q8Y3fF6iXZgmld2zOuV960OMF
HdLbwIcVsfSrJxC1CEOIKUpv5HZmnB+qaF6JNGvCTx5/9hKwaQekap9Kga0Msu55f5SulZg6GDTx
B614aTz16Ugimtpk4piHqfxkQs/QfLah6o717Zkknn3x9HQ5uxl/+4m3YzOY0AMhs7Kw6zkLtAWd
LqZJqLjZMs4oar4DZIOiluMT9lM2AdRwrPU8hw5xT9Aj0/UXQwICR2sEApCm8ZFN0gD+FwVRyuNB
TcNibSLj+sue6LdT0K6LSCEvGwWfcsccHa2Vb14eLoQtiKt3LKttwGtGbGCF1W+vqBt41eNSvtHY
hnMvwTqgesSLZe/ECO7+RxNnXBPW0NAci6jgU/4lJadwr+VAcL7eEhMbYf1QKYiwUn5jZTACfzbo
pzNXL0p7wDGLWsUa7siP1Yig6gzXjKyUGAww16FXzvtz7uziOA0DwJeHaXy8fJCx+pxx3FHNb461
8HHhOcD1c7OJHGjeygg/xZC8gJKHL8TS2wZ4p3QXyj3ZMpZDuMw5MpNXtMKON8eEMCiMTPRVbcRC
j3muernp07ApCCCsnaoKYmk3gz1/iX9qxUmkc+JTqmXT+NpGIgoktD3hiT1vc4jdRpoSXyX9Jxb6
b9kU3X7qN3SN2s2wh0H5wNZWpgwwlzO/ONKfAAgVWuuAX22IDq5KFWwBU5xqru3TOOfulOfUwly2
lbObHSmz6A91bmtraNrOTQEj7Zpl1L2LIVwACkyk2w89qf2vLiApyJYD/jF2mv2efX7bRNhnUURb
eVQ2P0TCxOvwSKZfqq39RlJVbrxk7He3JqFvTLO5JeLnOq1FxOdOurJBuRRSxsQ41+jUbNMGuQ69
WkUFSKCj/hEgR5ikiXIE0BS8VB2CIg5ideYZgWRBmIRCHbgiJHvrEBSFe+473ySMUZJLpkuZ/Y0v
rrxJDzA48q0l0PwifbDPQUhADt8obR/sEoJL9Uxfh09nK/hTAKQRgKEYHt7fGHmtgcBzCP0a5FWs
rX8l2DrzTDtDoR2gDTrLN3oxnMQyfYqzndJg+nKTFK2aRUJIzTo7homnxGcWemajCcfq6f3NbahR
W6gjJik2qYApgZNoMkOew7HEIoTlWwMPadrhfxuAZ6iFZT3o2rk6JPu7irMgmsLp/+UROUiF4NSw
Tx8HIUUqmZcAvPC0CL1hvEORxK7ok5cUS0e2H9XVGpOJpgCHM4ibONkCPAC7k6MUv3YgL3MTluJi
HX25U6yyVogcu0X7a9AKPDi7eRzW+swEBTtZ5PX3JosB4sQT3V0//cr+3CWCwsoIA7xE4kRoB+Kp
UjCF7149zLMi5NGvuHoug3EunvKoh54T1Zbt1geNbLAghL3BZxTwmsFiwsdbIn4BRHU6ZZSl0DSj
qhqeEq5LHkKMpFHFhJSe2u5Hm41E9iF58x2jvS8JFwn6QE01hxTdKyUloFNRx/LkQ7L5TcjTqNI6
UENpC5AuYnpCzh1Ps6PIMqoPo72dahZoT9npNtMs1u1FVPFXJqXTVfu5UFrGINDp3T+Rf5fn3rHP
Aav6W5ye+fREDejmg8y+pwmfOOj/gVCmCwHF9ubhv2hoCziUCHlIt/oufxmgvqew740hVWugaQ+n
Xm1zJob9H8Qy5y8obhbmLPnqBpIv3lUOA98OzYnl/fQRV7+xdUoqRo0E2UgMGGHFXEiwKtewowmp
5SbLtQLjVFzImfNOyU05+Li5fSIJ1ih5ffyGBZlBV1PG3M2hDMpfh92HlapwHmFh88BtCZXnfokJ
cAgnP57DQ9yNYLQcIef9rYRXbfhYGQ3Xkf2rAo/MGaY0xv3ziQT97ADKFr3axqTnzhha2oClsmQE
Ju8A72zMFC3j3LXt/gVrZz7TKdZGKxkSHdWNF4PYOtV+NipaQSYH7idKI/lwLRKYkxxSvGGKY2MD
buT38vJuBAn/G8W2qsTVmR+Vt2CFbSta+wL+tXl4QCwV5JQjEXWVwV6K3q9Ub1fC4XquevI/m4US
Ou+HDh9xmXOZMbae2jrWiX8WjPcc0jcinwJEb7vZu9yaqhcbFJunawUaPgcgDZkcaLU54qytv380
51x/YLpfExv7KOZ+rwnvAl3ULohlUVfSm9Swo3zckIeoAX5kaGnBYYGbTppnUaygpLyw5gDXAC/i
mDBEwHJuhl40HNMGptUGN3Op+0Ex28SC8+KoXXyUCuHrtLXTU7yoUeCbUC9KZLehCJrlk0BDV+e1
56ZzVbMmWbFPGSTI9wv/u4il1zL3dpG8/hrz0MjpoiaSNtdBUwG3B5+d/J5H05O6tfsvCqbX6NU7
SCl7Z24lChNypVZ9n0IdY8WHIf2++xD7gyAtqz/I1UEMw9/7r1K695GY9mxvyRE4Baq6ughL9kuk
L576P+SiAm+ccA9sLFiGfgv0kMwAd7VG1BG8HIpHqaDXjg/oX8CsX+oWFcAca1iZO89eyIAJo6FT
fcjAzWtkqozDJnIxnq0v6jgVAu+ee1hkr0in5tNu5Cgilt6S0ysrPtFTlqeIP+j6aiSFxySP507h
MRs/KkVHcdPqHfSWkd9DPVYWHNeUUQ4wd2oa+LQ764JSvh0f+6TO9khiBELsnh7fgxk2rx3UCIge
J7utamDWzpL3ORjKcycNhrpCkI056zcVnX6Fmx5OEL/Va1w3l2XusE93dK1agKooI9i+4qwdNFZL
tkTFJ7nxDts93egL7t18U7jw9ylPzBBc2dELpV6AQVyQ363llezLnfGZvlbI4OjHzDAYqk0Bu4Ix
3MM8bskytN1P4W8odcFozODDOmmyuxcg3wAdIJ6FmRI9r3HdZ1bftiMUzYvddj1zrLmnGwzjFka7
FV8ROP0aRzO5EPvjdR401hGTR5iMkye+Saaw/wpjPIRBNtWkNWNqDxc8wDTD10mLfRTPp5aPbmVw
wmEan5B/bth0rFEeDd0m6F4UfR3+rgOLpzK29fw79MVinL7cd7+Xs09lmThbLYqAv3ydvt1vrzHQ
EDxbGNtBgNtQB1zobJe2esSBX5sFsOnDCi5VLBd9eO+MblfUFBgKzBUXifSPUUWHGLlTNfgD1jyw
8IsMHC3iYR9q63W8lxaJrsmYg/Arq8e/4NYxJWoJhA3fBfSrt2R7G8Wkz7eGojf0jdDj5V8Ue/cm
IUAdyX9MpER4rI7cDpJ3B/4hsWjoPsYfkzzf+XjlCNqGrLRxfX5M35/ChHbIsdho4ZX9sAKuoLqV
OlUrQPpjX4USA0V3tRYD4NUWJVAR/Qva8DhheTnuyJ1DWYfrS3XUCG/St/YBjeGD3Llrf2325R0B
+rYcw2WGxkcX7h7VQBJIwajpGOc69l+BD4XcNO/35WWDbAnRCS3+CdKQ+iQyfmr37NHUaF85TJak
G/zLQq6yZyBOkJ58FyNumVORbtXgLCZtg7yUZfeHuPNucwLGhVuTO1J30chwg43vg9o0Qle/864g
RZ9zxqcaiyPSdVmtlTlDnuOKHKcpVuYg0arF8dC4Yh1ZkbwuPbwmBkNBimkn6Yqub54DYM8/51b+
S1Z8fmyP/qay9nQeEOehnSNKmUsNyW+Y6pVV2O5YQlqYeymYFKLp73YLpIa9CkK+BpHUDMEsDCQI
tdDvbzAErB4OL0AYBbizO8eQek/DT8krtjeQeJlBI3I2+BwyOli6VyH5BTOiwCwG2LcaR/L+eJJb
oia44MsCZmbMaON51LvqeedCbuG5qqvNiyP2Q7qFUFGXaV/WfK+L1CI/az7WExowf+TeHxxaialb
UU+pP6lSRXcMU9RlGYUql94mU8BD2L/Ki/LO+3kyxQwgvGPbOdWEAmnIQaCuAVw9JNxfFv4oTfDe
erQz5GXna6kvYBkUO7Wg8F5HN11FaIGdBI+3dnjftBti2Neh/hjkkL5mN9jrqITkYMajXeWVvEwo
pE17o+V2GYq3p66RaS0t4RbbxMd/VM4lgLl5QTfOM0BrazU+hkziXYP7xmRMK/UbzLMGZ4sl564m
gTJOaWyxrCYSilIOfl7UNfiJCZwJnKhaSeChuzdvxxyAZPszjZwoRP6dV7OLOJnc099+FmXAR52c
oybw1rDDOCrY/D5fwWq4OOE9EGqC/a2Up6qOIeHedN5PGVCaLFWYY/AsMBSnCtjzVvNuRqFCX9qg
/krikfjw9g1qbijTMLl/hgdtSYSTk9ZkDvM8q5M2xVLZhUViniPq3e+ce0RC+7N4uVgsLTqNn33Z
bpA7zrkl5vRRcI5PTXU7l/ZB3f9Tqf1Mp0IA5VHJV7ao2NTtQYz5q4TcFTlgjKVOpus/Fy66yt78
o7kMdLdlLxn2rpTRDdf+rHeEWyt+eX/JvhQ4GqcniUpU0fD1Rl0ZOeTdDjObnYGO9nLZ3ogPyR5v
iut6h6x5QKTuVsPuWXtM97JixG/QbfdPqn+9b46nrZUeVLoc8qVyQariI6DFwN5TDwqhI0by2E8U
7ltBASQUPSSAwuMimPoFSnf4USIbK14XAf6zNH1SpTOIeE4olmLhwEfmBrBoGxF3BAv0T9zHeQUg
/OtAdFYXcJ2nCB4MO4O+Z/4yTYfRD88ZjjLJV0dBRALXaSbBeE+vHK1h8erk6Qth06OU7TF0Fjcn
Ht8C7WESg6SfObrwL9X58+r3RB0xEIJB6KBoQa2mWpYT1R1P3/9JmP+WWa682r+1UjZwbQn/J9dM
S8wR4N7nyLCoTbrEMG+f8bMEowIdcRX2eEiJBeee5s2Re7sd6sqaDVCrMGaLXe5lzIBk9KsxBiyI
yUeRyVXSKUK65yKoxCcEAPhcoEGAIqXdlaDATewYcAfPa8s/g9XjTG0uPhPkZWik8LXue3TNwh38
Cw3p0ObGvpqf7WX1HTMds2dPeqm4hfDOuDIzKNXcgDJdzAN8DqVIDqeb50OJGNOm6KzSNRoF6ACv
ppTBVUJI/YPLGxmjYiLnQ+KYoTTicj4IB2jo3b/QpHJvL8bngxt57O7T/TS2OLBaupNFAQIzew0p
KE+alPvE/XUxU++ZXHKhkjrdJX4944ZR/93We1ml9IbbGdrCiNpwMP18VQPvxE0tNA6E9Si201Hb
5hMeL1nO2Uy1BmMQucECOfh3nHuZXKYiwhqrywpNUOAb9/2l1tYS9B3DZMieR54s3O1wGqZILitC
YZan/k04S7RUflb1BwUHjKZBjShBx4+D4mhC1Mg6YP03pb+YIdgnpG+23wKRb5HMHs7iOYGOEg6a
Ek0BflRQxdN0swuKcoywesR6WtRUidPxfQODxKJaccCxM9YVCgoKit+mUAV+n8Cdug9HoQU94i6T
pbOCH9w1Iw9CRnbd5DwpWMPeI5Fr9G+CwE4LPU/xC8gB/2uLimYLkJr71IElfIRM8Yo3hQI7N5pk
Dc/jzIMvyYbZ0x+tfpubbCNJJ9+C8LEnePFRLgjKznU64e5Ard4UR1sD7k+iR4c9aLjpSXWDtsUW
ibwZRBkP9g6QtwGBhLf7e2XyA2SISoJr1QOYquDfi+UTgq4Vba5D3RLptMUOK8uQaNy8E+HZy6af
IsArBnEs8HYgyiktnUi3WborAkwSjmX4nrrWA3LfqHiO57pYXcIzTWBLbVDtQ7MhFbvNS//5Cc3N
tkR0VvLY5l1Lf6f4ijJIw9EZDf+020Ts1EhvDENrMgcpMk4bOuU/y83kgIFSuZxf5LKZas0w0V9G
tJv/VeK5eH+3mMM3dL/5KCWOZRbHIhp+EPJlujiIwQ8lmwUUK5POCYh4LbAmVqXg8GlAgtSx5xd7
aP4OKnh9AT4AuAmHGpL7zT3SGUYUafmqOcgEYEZhJa9y/F+svxt1C/qqYLW8aUYm8PAk/+svhtpy
I3HJa+FeGjxGfVGvgMMZYVGFg+rS9wXFY8ZmeBICTjVEG0VUhfxoCHics4Tv5hJjZooTFcRcCYE5
iRLJP02R14dD+HlkhNyOAYpUppuwF/bjn9oiwT5n1WyD6bcG/zyAejDzewQt+YaL+7DOfJHBExFF
1I1fZYIDpe6CaTVEfonGnMGIZmAWwp10F1wkJMs/ggc6Q9hcEfTAQo02RDQL3429GdB6FJmTi6Ub
i0lKZw+LjZygvNlaB4uKj9q/ctONhtA/Arn1hJCFVGsGBdHyGPFQdOK87jxsH6HHL/PQqq2bhmt7
p2XYtrJ8AntGzqtPdXuklMWaca5h1i73kITv5tcnJZDC9HlCizMb2k5oigIQBSZpiErgIwIArBTq
YBlc4jaM1FSiHl21O5c+C03jzpq1dcuhm4HAr3dnFsZ00BronmDu4oqeIIjZae1UkszFXyRnv0tc
8XxzqoszPaVb9p9RvOr9yVgAeMCzfYnaOknfwq7CXKxs3SgC8z5hGPHKEQvC2R5ezJBFySWPjdzk
OSo9UjKoFsGa+4+a4iP01uJ89cWN8OoUsTvgOkcJU0cAIUzWdAIuJG6tYNWlWHph+RoMWLrxNsbC
+XUDRiPHd5MgKI4rXOzaUZxwIWpHribqZK/89GcQqMzV3J3cA/+tI3EhNIk8us92e9JSNMZnB9OV
2k9fCz08LYHHuGCmnwoTr9p1GKpEiml/tfBQtmvM07Hz0a8UpIc4rqCS/IP7i/ns4Az0qzr1ePXa
ZdFGNqaYH6LVa4VEdVk/OD182rm5IV/+SCL429zym3egwnbhcMGOsi3jYNwi4fp3W1FnluKeTX9y
u0rc0cWUvtXYLUvPXCHcx4ftCt5fhKK1QwzcHLQoZ8cWkVkQopMpYv6mPDxxUCDUak1PuSgcbgTr
W69OZjIx5ZRtuG/g7HokSeT+ulN9I+Tq7AN0jXfSfrH+zm0PG292L2QQqgIAnYXOv1+M5VHEM2qo
ZpzALwQO6+xKXBvVNqbnkgGpKXI3iYGyOznp5WJOv1O3TIWzKK3tqHZ42OVZRgWEG0qeW7nhqvVA
h0f0xGlRE3T8zjFxOfU7R0JjUUrNpmHl6uJnWLaP9TW2TnKHUdvNGv9rsYWYeVR0K9laYGCOeGzu
iSSWS6IZmKfabVWe/3qcUntJWInfQ31mVjJVUvTEOJx9KJjnAwVG9TZtE6AWaHV3XhF9EeW9k7sN
ba0rYCBERGDhaL9/h3e799sTzl19fyA4iRp6ODIrzObS3kwt9J2R0fkLsza+Q5tj86ZqDxblKD31
wDUN9PRvp46zB4TavKSIW+k8kW8mZDLpV95V8Ry031zuBUQa1o/YiDh08Q7ZObKg0XAiO509VicI
1f59+UYOIOmWuhBdiojlkucyebMXAGDwWWDPAHE39U5Xh+qdDlliNK5zDc44YP+C/isYfbTQPvHM
5/nQLn1zjMcld/xIWWAfzUZwDmL+yWYdXaQQFGZtmaO74Zc/1SZLJgd8LCwF9uP3VrhU/bR4LFQy
QRf3QIG8xYKnbQBv0R+m7eupr+WMaIpjvud/LMDmqfm0C0/FpBaBM/lznKyNjXHSwuVse9w2pVDE
rwccFoHPxegkDf2SMa1cyEWUOqs4RN1p4kSXxt9wCUietBd3hDREUdb1L6Ud537j2i6ovJYo3bNt
GXvH+FH6E6Knf456vY3s/c4Sww+4G+TM2XxZhx8q8B16aFkhl78JbRpME65KAqI+iVbl7bDkLdEl
NYgJ9F1AeK3aN5tHmxDKniUPX4azCb1AKi2Y6HoTu7yEvZJm1/4t6n0jhUsUBo0neufm0tr9vuNy
sTFgUW9Z0dMmriZDWrk+4keqv4u082MLLjUuO40eNRY6oT9cC5kmy27DvLjsJIR8Z3nrY2hjszrV
Kqb3QfALdGHM9tE6sZFkNs4iQ1A24ZQ2ky0vFudvotLB4U/K1DFPHJWQsS/NVzDLk54S/wT8zSPa
Xx3VJkbiEpNTUmGkEYP+RTmXMgZ17NFFwQSgkpAQOvuBjnElQ2QUPi7ca0Rhadb8aomfm0VxnhC3
NtXTE/mKR3GOVXN9oQld/dpGK20FTc3HSshNwcio+kIbtYSHAH0GhcBuuOA/HYA7H5J7UpFfcKSw
Ev9G0sM2tUl0JUnVwRi9p4BXrxnluIJz8N4yQ9mY2EMDHelXT92BCRHFZq82oW3IOUiBjhp4TE5q
8mixGDyY9xbsaQ0nYWUD0HfzT5rHa88OEnLsasBMMJ95hTi28Lz5TMUnGIqwx31zAA9ilN9KO+kk
+BLSAlsZzGMFF63KBaet/rT1WBQ51pYWlmFSnsmzFCyORPqfww84eqdqAiDMbTyY00GGU4r7w2LD
NJt73KbKTPNtFEQqDF0cfueYd3vgTTaIabQf1Ga6rfdIb98mZ1DPBbjO+BpCBdaKUq6gUti3+F1G
g2DESB5zeQ99ON1jAn75pR0Y2e3RbyoiRxXS2QL6/Kl8ZlKTlsOhn4mt1LydamA9RfbGXSQwB8rs
HrJxQndn/2sx25tUYCMoZYevu0p4xrauHhRCZRiVkQZkm9Ff2h/F4W+saOlnQinNkZ8FpAFlUqdP
QOSHjjbl0w82mJcpvmyj5wUEYS9G24xTVI/oYmgaM2rxHALnAim9wjt02M2ckXpjxku8jMSRp9WE
ozlsoWnRxf5vTpILaw0u5XpGpw8gcAHiT8OXleAoJwIWUaeRzwE/CsJE1HPAML2Z9B1MlQNx61Ga
B+Rh1RdCgFpXJo3ho+R/zbY47AYJlys//WTu0/EPuNtJvdH5WQJXJ9dgb0VFGN0gpce/bQ8dekXy
VAMxW1ysPA1FhkwVrO/Ba56pi9Am8EkCHIJokoME1/F7YHOxDYwCfnbpQv8sPGd5gg6tl6MYOyG0
orqxCZw2ko1zEcsCuoiZG5MofxpCgYNwmxFiiRs9lrtuZW3K1A2vLRH0HfMz4I+Mh/hMuZJNktFh
+WerbgRZLemfaZLeEA6rgGDpvUUGTdd1BKT84/VXZgnfGi+eO1HIG4zoqFj1B5/0LA//vSF5jlAP
Qqewd6gCSnDGn+cEI9h+UjVzx+eEk/rTaXIxoUR5w9ZZot4WjSnAe/JcAMo2Lerfjat8quYibQsp
1K3z3t140uxLCPhgZdYC6drE+bqMXSfbZyVcj7HayI/Gg+buZZzQ0YvBDUELoF+ClFTvVb5SDLzV
hjYA+AwlS5prLF7/UayAmeQji8bDfg+DOsEw4EnYkXZ9bO3UImUuWmB+VLrCA6fZwhv2qBHePsxR
jAahdJ8YBaS3NxAwLM8LwjJzqQhUfkS+AESHebMZmODaJeqv8+4Bh+UJwuYLFAX5F686Lqw4ZRDA
6d8o4wbihNOdaG8FxmvucJgY0evF+gU+q6VBaBOC5kxrrqkcS5HX8kV/EpK9tO2hV9YbPmiX0BbD
3k8vik5hMvUbKXPNiGF9lRhXGBdLagMLd1ZV9EdTbcuQVUfI+xg1vNNxguNwLmrC727UqgxfMxXG
cTvB/U9/xzOuvREnHJxsZSWff6TA0we0wcNRR1sGnsBZN3/9TNNtp8KBUWW1l6TYPZ55wAwyWp/7
azax8rdyAKp+mFcUxfK9oWMbN5zmubgknpPsQ7Qhc4Q75z1GUIF/jfo7uE5tTdYE+6psNsk4dNWa
+fQBX3D2xLPYrSDLfJHFXS2Ooq04QmjzQ24SeKu3GiLeLteSZ6P+KjIawdeOR6KvK3Y9j5Q6k1Rz
t7MEm37XCrNWhPZPg11Jde1avdizDiTORqvE7/ed/yW6blQ+057PbSdcmmudhbpvn/N4u2jljNVq
Whz3vLoBH3Xck5hZhlAI2hrCsgeqWo3kjj5SU4IjaH5w8VxQQtN4ek/tDhGGWoHwlzUUWSDW7n4I
FxY3CvzR5ryMSpgkOcrCqfKUnEgoOBEcL7WJLODOF63YIHwpFdKBgkliDiryNtlMt9R5FhKRtrwe
BTJElAEQA22Dnym9u8RnNL3uyXq/I7r8zH/N04B9TrDoGl2mzwYLJFIdWgaPh9hACWTJ5Ef/iiDD
2SEDwx/hp+pXJk64aJACpMjRZWl9I0VDaxdiLBVcfVQuLF4MwSQAJ76FsZmUy025o1NaNtlvURA+
N+uZ3QVl/gMrUUkrHVq2xxksq6MKUMGzWB6eoLrKQVKZGgP4k3yFc/FbxIahScZ0JTHgAUHf+w6h
bu4+M7vIXzI4xclT7NgGP1r7lIDQYUqToJKLXE/J0PDrkpV3ufAC56FrKXYcr0RBw30h6+G/Zljr
l9bhUwkfzbUan9HpQ8aHhpHbtVJOKx/tO2dHIUg28bgqS1KrBj6Npqzz0uveFZB53KZbB2XWvv23
hKF4Jr8nkvUBPuLB5pAAPF7wHD+kUW88mPt1JcRGow7OT4GeWOZvRUOJmDpFTVGgEAQ2sDm0pw8f
sIZeFxYrv3aklHIHTHXXhPGmA0KXdZKxrUbDk4nN8HBnydwxcK08UoXBmYFI09QjqoQzD9BDE7kr
pBAYZ2xoumA2mn7q3w5lUeYLTLmDCXpIWvdiXo09wFqsBeUxt0dT9DhRrPGapTy6BLQlPXVrXHGV
PoINB0436cEsDER8PDB80tj6AZoLfawE1a+0FWbIUR/DwmET5CgT3YdtlV6OTfbL0u7QlIjHgenX
8/yz6KIu3FGFXGFGWf7T+A8Xzc6yeXkcXDE+hhjoteV8nxvh6SSfFT4gVvD8X+JrbJKrI3VRby3a
v2WmvVw4c17tHtmlRIDccdXnSweMbt6LL6tFUFKa1JsK4hXMRexK6rt+u+n6JDSCVQFNfpDzKnck
s83xrbhKeq8Q4HA/6kppB7ZsiNGmR/8fPuPEHfjZlxUJGCRn8lFWGT7hn/ajP4cIKH28BYVu2PXA
OUueGam156JSv8jpVxR8ai/hQYLW08DQKTXnUj/kK+DWxoKfabkDmpixfW8HzNYDWZQxAGckWcWk
lBR4T/JbiLW4JfVGtN14vcaYaKvJ8jIVTIQ11F4TCsfVJHyVvu99ABzKF/zARRjvrWMIhe57/g9u
my5NDtIHvPKscTBxR914Qnmau/S2qY448iKtbvFWd+SQ7vrP/rdd102lQkx1PFqojGuccIFlJyWt
uUuL68PHOAEZhVEVlXfPlJjJkCXInGRC79wb3XfOhkIFve2tNrVOyF1IKLH1xqsPf8WMdtiGMKm9
YrEx8CsAIjSSvmhc5KRcPzxCoTd3fkquYWleSyNrinvgzWAR1N1NoarzyBp/2seMxjD4ZSS2Jb5L
iD/ut9NGFFK47RbJjrBH0F9vgMl+QwxZk4pWaJr4IGiI/35YMGYg2pFf3iDGCrxzImmEmRDGnx9c
1dp8qQGHIzge7fUg+d+ub26Hb7b0OppeDCgxIX0N8w56czyuZGwB1WDOvZcsMSUIFuibva3GBEhn
gUkwkN5eG8QPq51qvwsBtgO59fYjgsdkfL0bWY5zBDw5JNvzI/3MFD2KpIaj/c9n3XQEcse9AGEp
8VPfHCMnKIxJQfsPhTUDDexOUlSJz1CmgPnUFyCR8cNBv5wVYmAmdJBhAD/G6H4JRBqCskojokFq
XRnvJoguJyGz+4Hbr7MqkyMk2rsykxvq0QhH7U6Zk4TuxBwvLVINLhQfmoc3qy2E760e1KwBeAF9
uEnBf32Q2UvCnojmCCuKK8LLQnHnwScFmAmng/NfV20wfyH0F+S87GhOaCv8mLQaItW43W84q6YO
pLEst2uSpmNNUJC/ojYKIpxxUJf9ery/vhw1VAPAZ6Q2Qe7KtrLtA08rjJGQP1UVl59CC7XQvPZZ
DvwPeElCsgxwftyLRKLLRQ/s044IkVH3pF4TeVMF9kePkP3o5VSGbXev+euCACKnZeSOXhQrM2NB
rJsOA17TCbrZWhpI42KkswihwzG/s6zX04f8T+OOyxvfeSuRQXlnfIu7slREhOsZGglkY54lBgyB
/7hs6PHxVYuZ3m9n/+3rAb9+MO8y23yEkneW+wKGfEyB0cijqCHfPZmtcnkITaNxqinxGyVUlxox
1TuG16WQPoIXM7SXv11fl8sLWYf+3iCbCk7KlyaHpUbHhY4KMbY5drpFWuwfR57khlrpkOs97B6J
5wOHmipaUI2De5tsBTiXPwe2Kmpt7gBtoNKOM34PO8y/oQjn0LGTomtPbOTfp5A8RdIWL0PNXTrp
UHJ2J1qYzkuqVwrbr06CovxR7+Qf/BAQkoXQuJ1/qZ7yG8hh1rf1yBxXTzyl7j7ozNPJv+J5B603
fyEaq5p4nnt1Jdz8q7Lm8bVu5R0tNk7U6nwE1tFPXS5XtC1aJ0tIth4nlO6zKERgMvuZ+zu48Lyy
jErrUborAuFL4FJCVCfJPY+xk9cbKE3HgSThqYmKGH0czYZTAGMYGtUmFzKi1pFB/em2QmOyh5nS
r/laBvHXiJ2I3IfNBK2t06SDeV9+9hlZ7HVgH1TH8tY2c4sqXuWzJeUiN3J7fqWnEgQEdFW4k+bR
DnOVuK871oXQ6whO9kPd6+zVfThJ/AwmSRa6KEsakGcRQtCCNupn0IWgG5U/IU0oCgqIGXbSa3Cw
0EhGzRP1VZaolU5DPyeedXl7E3tlxGvjBpJUN4L0p2TD/FoHdqfEkccZ5m4GGQt+2X42JFzIpOnC
Hc2t7sjx15NcQCWcTbz9rodGfHt2nfx4g8xfxxrWViIEBoi7MZeRHGPNyiWjbETZRcH4OPH2Nkd8
Wve2JtBpO3o5pZj4FgO0yYP+U7MCgDS/QNgkij3eGjryWryyNH8tiobmrYJ5nvc/I/uatB9q+OoS
IWZ9YOXIp+RP+142V7skpKsLBttmAg8rQ+Tp3CXTc7ZNjCeTd3F8IlDJhEvV5KtWUo7YjFQ1H5+G
+faNCZBRELtjWwP/MMs8gWnCUc/5KCmGYwjWbqC3VIdotLlPsF0dGchId6n43rwlCGE6uPL8Bks9
tkZsKOactmr4cbmi5IJ74smh7W/SQrsSDdXkK12878DcIrDQQ4jRZMTKmCJrU17mGnRRMjb7AbX1
K5N97hyUifG6LL4wXMf+r1hoDCdK1EsrLzuHqR38Gc4OGS0UwQdk7vnNpCG13p6fFcJx7cPCt33T
DOpcwBPxTRrc6xz9b3CDFyPLSe1YmfhOrNBJkGW+ZfBnPjAEq5juRN2E0TyHmfRuy78+yNm8v32r
cYfA9kVZ36BwGdbMUsmaiPUrbLk35zXuq0WFjeFCtgxzEJNn/uOPEDc0I3cLUu3rqf8FEkA66iVl
FFPwqGZMpoXBcwMGPK0JB1MGw8QJiU9yyeTBw5bog606wOBS9MDb6C4L/uS0KXi6WBIH5e3dILRB
99wPqXk7bopnfb2xeVWkhaQ7tSNQCS+gIDgFxxfvBvGll+dvmYBajezQyzpdRo83EujHTqOmSFh6
2VAzLDV0hOSAuNHxgWyc4s1O7XgtbbFifYWH5zzvtTC5oBbZSyRcZOHszWf8KH8ZoHe+K6XMgZe9
zE4fhSTertcTfJXj6soNWGsMvAiDHlmiEyXg7QzwuKFfDC5WJGlCduH7dzO/iCcKaLwMBkVYP332
2xG+QL99bwiZrHpDTj94XHC+/BhH/+p3kwifGOqStbU8pO7Rwtadz8o+w5bYAbCRRguNeIvBh3iS
swS7adK+0XcrlIia1S4EV2rMfsbCUGx/SpfsoYIbGjLXtKvn5JaywZeIS3O2tLR/ckHPhGFPLKwo
hk2wmL3AC9oZdByxMLadhURFx9lnGvqLriQqyM7OWwL7AhAnc7fnEVVzxxID2dO2WhVuVza1VAhv
3RPScSWGCj/IMbiBjSbCTaZtv0bQp3AZa4LSKzWTjRNrcORwhj7LlU5gAybckPQ0nZ/E/BBG7QiN
C1qZypklDqFpevUbpm0TJoKatCJf8DLuzn+3qIvjENHM6kjwb3I493vaJpRdLLqisnVYpTQKwGU6
e7gHGtX9OAGXeRdiYqlLRixV3b0ts5TULJdc70uMjeHbaA0vXEzfJ/q5X896JjPzYeTt0a+a/kZW
tseI9bfGV9ndD/PKgJl5NJ33wsgTVmS8GKUcPQuVO4W7IzOh20+w10gEobQMd90kWE81rlY6j+18
q7FSL4c/ifVdEywaxSlX0nBH4VgKrejuAvIdgVBB9mkU/T2QWdw6QV3kNsQTPeVHYn4Mq/X2yTNf
2gSmYV2Ie1tS6MSSB+4Wfy4+zqPczbJBUeC8KZrZ9Kt/JyA62zAxrNbImdJbVhmmKrCA+LIIoLgK
W+HZFTIzE49oVYigTU9R/XW5TSRExNhvu/SFw7RwAnP50N+H8eLXEpXfZ6JWXZm32QsaUoWulKKi
xmJfe17ACkqvC0yTZ1NVXhzJ+abrSZY37DCzhexXZir6wWbXJa9bMelmKKRaQ7WOOjKEvO8fTtVb
0Oo4i3f1Bhy2MZSlEAgnq+3m5R8l1v+mX7I/7vNIpU2hqlDvKdLzpE7qKKPXVgg3gi31o172n1BU
B18eVOGaudxfNe8JcTsFZyRIpblR7elfWYnJyR8ure0jPUX9xxbpUo37Qdw8HqOSzOujw95KazoQ
XOluLS9bVCzToQw6EYy24GqWKMlVN0ZrD3qRYRVQXlTcze0zzBLMaxcB/4h/22iM71Q6XkGP7jYb
Tak3H+6A8WbXgtAVjsJdkUpBCDrLPXplygNhOvsUwro4fkqUeAR3ClOg8Z0oU5foZ+cY62/uOd4Z
yeA4Ip/5tbVbGjX+9hbzpjG7sHZPgVqNoQdnJwYkHU6ZIsSB2Oz03ghMcoKvJNGm/S05rqrZBvQF
WtZtk8e3CJQhj2SDcB6OFIa5/3XKf1Wlc+6xNpeHZ8awOOXIlJsgsV0ihLHXHrBwAkapP2i/Df9x
7dbEMa8ZetxZZc8Fp10mwLzxUZmCBQM71VBYVTxE5fJ+yCeQ4xWgUJk0ia3FZdVtRYbfVKjKddR5
l3w+ru1XAyo0rLlPP2eKEPGW/8KEAv1bIf1GvfV/KkiwCG/5ZvQEOpny8PrC+QADLQOEct1bavIA
ISGFz83o36zME5XPcDBInqfNlLIC7vTWsrToKelmu3DyVDFGZHtc9qE1J4ew2oDdB+GJ3YqbJFZs
WGdXYStaDoVlRvQ0v7aOAWjljeRVpP3HuDFsHpYixpbVuXVR/tP2kEvv5SUkxpX6+yysXt/80zM4
6DeTlHySEat/XVvuSC9IAsY2UWYv8roSsy5lswy7umjluDxSQTdAFXG74+npgSiqrSE4pDrfPk80
lltIFuI8rx4ICLP5Xlrzvt1K8oTQKjHGnwHjbtKP3PThQ5zMyLRxCeNcd9vrAUvD87J3DNxmUn+n
9vzAoWowBWZj9BwUP6cuCIan+a6rHfDkca0oJErtRPSuEHgOxozjAGQ2mQ2KVK0l+0ymw4WEMfrE
XeiRG93IBDO9Y9/EpFMYTCbWn/3ymX6NDkAl5/uhkJxXQatSwa0dpqlK5qVDgPZk7nEL3uRnILVE
0m9k1Qnaf/V2gO4mf5oV64RgaCqEj4sFszs6HrOc84GBp3A2b5R3B+a0qpJ7MVRTvIKX6bqnHdZ3
HiTX4mK9vjWn0JeSMCzWUHJScMbASc2weNFXMsjZINVEEUmAQLq9VkahOXKbyrFs9GKJADp6IYrY
ZUohkhMbVs/Az4F13oQ/O0atNPKxuW8A7dXdakBe9qvjIuFPBrB5q+hKIpf5xZJ8RovozEMIJcbS
sK4Mp889drWO/zGV/hBiDN/GbHwgoqLk7WG2zE/i6mdh2DUunoUaFyn3tIB/Qa100XOwZBD5GUwm
i4AJz6fagmk/BVfHsyVLjn568Z3eNbmskpoGjrUONQZsXB6ZAxCVE6V4PZX9NjYuYIcrKdG18iyB
pbqtfI5eeaBwRkNo4fB3cKknucu1QUT6WkjmScR5VZ/GUsq3oExkc6iXR21vkxsoAPN5b/s8xqZc
7Uq6llFnBHacjtCrlUMziNQ7i3sxBSk9nS6IaPHYFWuuI+NEDhGWWhEeFJhI48cSAysxqxRpRxU2
NsSvavLA+E0TQ/JsYewUKOSGtw4RAuA7v+Qutms9FDmE+D2fAmatpElMuh129ea+RD9KRagqJGz5
N2BL6/inpw8ZCerclmdNKWRF+7tKZA1hDMfG9ZttMgRq/TYlDA6MDmN1gwmn0vjyEVXN5c0KGPmQ
9KSDknQfbP8r/kO/lLZr7hJXfJ8kS/pzmEVT2YqClgTdMGz2TKs/jIWBfBuq3RwGczUpquXLdrol
GJ/hmj1siA2YB7GjjWljkNkmtIITMDbBTwyeZXYdVzO7HSpitwBbswsAaPlDudFNkZB/lXEQKlGD
/ls4vTZBYlDYaLi6GvBZae9i+1lARS7PkOguvUPE7WCSv6qzhhMCEkr7dpYXxSAOsGA0iorJGh18
NVIjZKYGjyllIL/Xixd5VdfoPqvn0gq1UoMgR3ZREPiTTZ3305aULpzXpiuPoFYgwPFjxDzEk0b2
zntOcYtlsd0J1HpKOwU+PQ/1wiKcTPi2nv2g9ip+x8WMW35L8oUtID7I0S8yfKgnjb/8WLfFnUCG
n9T7t4vx+RgPbnv9qIm8Ewjuimglxcg39H6imbiJH6ydbTH6WYlnNfT5dX8FxVftd/MaB0ayN1w/
Dqj9FJ7G4zrvDtSWheE2NAFsNCdh5kxNzEaE947XEJd/u4/9+HeT4pbvGICpQoGOctiE8T4o4pom
5ac0E8yEuX3+B2VB1OZI0Zq+l54J73ZbTEcy5kF5tE1QfxcfYlSAOVXxzkALiro7KhRl4pZ7iDTB
Hlh1yjIq8gTCJlxRk8KgjOKZQ7GX8nxjSX88ZVRzM2jPtYQTauuowuzRiuLHGXmBk3aVCUFWtr2r
kqiNr47NjBLgXtPKvGluLHZoRfQuRtXHpJhHZA9ESgHWmk1fHiXG5c/AWbuuopIIpXonyMMz+Wr6
WUyqPyWMHBpbkeoxI8Tt3SR/4JzVCZP9uhh/Ceo1bRGsrAZv4GjpSa/F1vs+pbL1gImiq5y1fcXg
NjLBpJLmxQ1sKKf3yTDFmREboWwR9ZF/47vs9O12/e3Dh60sSjtcjnGEZFhueLC61Kb2bN/aFdE/
7airAAIwZ/IsSU3GDsYgPbAYrUIil3I5XPcY3uv9DPZRraX9vRaX6fbW6NwQ5s4bXzd92DcnBafk
R8eLLZbl/B9nqb72tAqDw+LK/90R97VyiwcYXxkfihIMRHyKCl46zVQRxPGR7ZKfA022m7UufkxD
VtHYrDH+UcyEpUgjwvrl+CpfcXvYOa8nXbmCOtCYbOfWIO3tfOCQxN+JhCX6CFk1EbOocpJeQ6yH
CCdu1plpyH3n04ZXVucRpDZq3c2si4z16AGo7ZBL9STWHgSukBqwJEDBW9LHtFfT8E1ZWWaaVGe5
/yRW9stXfnou1Z7AwAUncenFUqVmpKE1gxulOg+Kbbv2kkCDw9mUsrfaJgjpXgQkix8GkHRomUO+
53/9kIun8AFY8HE3R3WhRaZsFh6rX1Sph4E6+ewbQ2sII2IJHVjcETl5kXGhRvE4rHmFGG9vNaW7
3ICfabDvaHDrkyJ48RmiDe/HHkuFzOI/FI9+McrWyZZVb9M/BAbzWoqE3rirOQDIggE5yqhHPYe6
R0bSM2t8YB5oYiIsYPv6DaSRnoOz0HP1ucOmDQrr1WgMw5H0QdYVpF0fO363huBBeuPT3mRuwp2H
gjAbt8/CQhzUv/JfH/UmHCBZQotBgbhvbI+lZ5TaodJP+Bwd+VnuJnCP8tFjXQzJCyNpg8WRSvrX
HvJS9bG5ySJrfng6f8dr3iVAuBtwiQcRvw3oUz6gjBy4M3O1gCXkj7+Vy6k18woB/+9A9VUivB2R
2ZHIII0mAIJo9YWt6XlD+QM48r4eExxRDHUAqNWfTnwqrhDD+LWKvdeMX7WFO9UFdCOvfB/P9tGq
mkPnLSbMhP2Y3I/fTuXAAnzpBoSP04j8xIGyTvmnv+pCuBVUAoWY7vgrMoMn3zxIuPLm9sZuo/NG
+kKhWutEMYthMBaIL8Cfd1xeV0sTglpnQItEAS+rSSf12icaSRPTpwGTEpdaEI3rqv2ICn7urdX4
GGqEdMNOHfu0loV4hkGoWNubnV13r8G3PSea2WBKMzgu2uP0xr8Ua18V+zSd6hBWqKBW80iTzHzD
LCyVpTudctnGd0NANTKUlMslUwfTD53x0xKO6O0JHB7Y4gwpAx2DNZlpX7mfblESUzyuZyl+6qkp
gd7HFdUdhcjk7UMdD3Rz3ramh9EKEdhp6qKvZjPlUufafGPHTD7oSNdwbzGQ8GIijf6uPMaqSnw7
1FlXfgEQ/FMN8JFVIAd97E9f+o+I4NlkewoGUqOzgAFu5gPMQYOr/k7WhNUZMYXQ+U0oYxDO3/DW
DSMM0hAj9OnjhjmJ1yG3lgv9LBnULgqQbaTtVc3bXxIYXhJbncNu7EkuKWYI/LbkvCd+raFdJ9qt
IRSbQOLGOIQ+GrjaGFYjeslb78RouxFaJNTKz61HfmJdeM9EmRul5zhTihqOFO2M4D9JGkTIZ7s9
WS891NijJdGf6YjU4UABj67A5f9asinCxLbMCN3JYxFkRZU8Tqo7uvFgKZuhSE91Rnf8e6H6jZ5P
QqKhV9SalAi+svPBpse1RkqzAR1yxPiglSthUvM7fe2O5RsV8znWQwPqPEvnQdSS4bBVRjTdZHd8
98T+k/7CKWfYtEy1rTWQH1nytJW+G8zHapQKzKYt/7XCfaKss+Ti87cUsjVOd74qzhrsO3snBf8M
HboPZWp2SdDhfkvqo4M30avsKuhJLZOttUrAWNQUVnXk5EFj1R8QSlaxbyVroidlpMWn7+PGvfLs
DlINGzSoJhK7sHWk4gMqq4ouBl/y8iZ+pLjIX4neSlnLCDlGENnlMK7TRAxv9Tp6BkdLG6rS+wce
nZaHUIHMmkDQ9rbmUUnf0C1dEdhpDY/SFVlJ9w7nxqIOnq2aOihcH6Chi6U1xZ0mFd0+OsbGU6WP
yKrqU2LCNXU91yqNU+dIuCDwUOtB9H0f+opIgQ3PMlerAfOL2azxUZYdyaQFU0DzhslSSljVJpov
vk1vWgKpIDyPfFJBwuQxtgEhmpNkz9ZRWdhwPrt7+tPcf5jZr0B2mAkA/HpB1kn5RSGziG/ODB0Q
5xR1rVaUO+pwv/iq65q3Jo9N8BWMZCgSj4n+V7HojPq3ynVTYYoxEAQTltCZTYlPY0xz0oHERz4+
NsH5GtlIlCIWsmgDd9ZneYj1xRH5xZxcdHNEqJDxMEEJNluUaarNIx+bNBNPKiKlavptJaHiPSA9
6dhd7PRUretNeVONDNADf4+FSM0kxs04Z3zGoZks0T9YM0zZIHVB5/gzo9wqmOIvXuPcuZ1vN/oR
7kUixMBIr4CJIS23OeIXFMJJciZXcXEEusz+GqqXBlP0Ef3tPa0eCWNi/hBS2AS0NLtwYRdeB1jR
oN4SoS1kls0L4j6GBAoK/ixJxn0Y2CMcVo6hnaQKLeV5q+3ndL8K5Gz4iZ7u/1LEXCMQZWIXp3tX
HAJ7ZPLcRFQWGWWHzgqJH0mvh+DWi1kV+/sAmt2qZMVVjYGlMQHHf6H2wr9MP/78wqYkjMOeBrPb
rCCd/jhou8Y4jzvgBxEb30ycJ2pmGwTot4bf1N6EyPBCQNjVmuJ2jhaOLGko1XhGjG1HR8raCtF6
z7dg9BmkuhiqMybkiohy5APuszc6BBOT635pA7vTtDM2WvN2K7Adcip3/b2wMGaFL6j5w19WwJbz
VkotLvhOlb2kNtNhuzut57Uga73e3dnKT9Phwx8deXUHNRLSt8jlUQ0uqErmt59fFWtpEK+TQ1aV
oxDhSKInN65LAngK/ODTbfp3RxgfgByQKfY+Wd5YFUescIS6Lkea1/KKUmeXCD5EsaF2/lNVO4JD
v9aiCnHoKgieLGRkG6R0gN5krQNOpLpAFxwkVdwx1UsMvINvqN+dhm3UK8xZcRSbLONBYyvgiZIT
HHmFS2IC4nhWLGTstDy5YoohKBA3PPQC59HY6uNcqtiEC+Zez02Ch3cbRb9/Q1mOydjuqO6pH6hD
bupKKyFHYhzCEedzlgucBY4idR5sQ0Y2pPJNr2d+aijiTa0leJ8qLQvNFZll3FNu7DbgNoj+aKYM
SqssJwBKl/kuDFoENoOeMb6ymT+g/PRN80uui6gRQ0XqyyV0krByfJPLjQKQmRri2ENMbwCtn6Ht
lmo3KPUaqfllQJztC6CMcLbmVCRbJaMCCLVCMBPbVGKrYWDJI/9huHT/G0f7eCgDCzqhQZD+Kyqf
mM372V8suRWDCUuKv/Mrr8yCCpdNUz4TthWE7hyV8GPwGIfZXGAcQcjoJng9PjLGidghuBLE/CXW
v6Hy4KM+2mWt7Dr0GO63WZZIlOJKFO86Ey5Mw1chLcGWqlbGZ+JUDQ7zKq04wjw1iQKZjU3XhgZ0
d5mg5MhVLDAJzQjt5iYdjr+kEopGLObNY+S0wxfivD67Iay3pjp8tmp+5JUtUAuVAkQ5ZsYcMLjD
LXv6YytGpl6hgtq8Ro2DtMRGjq/c2RkV+X1JuRPgEN0EuvvhRTpvlOIaZ+uAgYbbZNxglVKlKAyc
B1YistaVEor7DxsE8DkqkE4Jwes3wWqAyMkGHhJPSjq4mPOxOjhr2ewM2ACmuP8NYElIjpANH7g0
/2KPjlvauUeozR9hwf9A+y4S/Wp+Km/SCEQISEHrxj4seYpBnsMxh6X0X5rC36yyGrQ5gKpmfOSD
TZ0tw7oZb8gFipRvf8OADayU3B3+ObXh9+LObf/knBAV5p/SmhfEpVjDTQA8taljyRdnjIzeQIOl
g0KwWlypMmmvn/yG1sznHfJ9uzhmyF0HstNToLQAI3ZgvM3ACSjEVdbrLV+tOFz1Ke9jJOEuxYxS
jT97D4C8tIDLoHM0Kg6eqO7jir3jTEP8fOf6Mctcf//RnOaHTx8+f4fNcR7kDCg+G74dUD64HPH2
u1Z/GX5YaPT2GDv1Z3Fd+1uv8zr6kIPPEHpub1S9JJwZDJKLc5a9JHhT6rDah2rkM4ZNKuvr4I+b
wFlUfuplwzsn7p5xKI7EUF+KvNvoE9IHsKeFIuhILbczhX+syx0kiaA6rXteTHOx7nv5+zPX8Ufk
QJHKTu8CMyWNA5uRmGQvcCbJkWZc+MVnuBE/dgeJ6IdjjzHTGK1j1dJ8x1e0FelDeJa+JYRsGSZQ
EpN4B574ELN/l7VX+uyf8HFTuuqQsnMgJ4ELy6aRnS7KhD8yG9eKcbBhnK8sN6KgZzrkBjNdRbL7
IRCeUD+hqLXZqWUXBVXkj50saJ78om4ih1NsMnngnrHIsfqcpbA4WlqsbnZo/YwKxzwW1UeQSHLF
vSaS0B7EQxRtqin8Ifg2DcF5dZ6SDdwrynN6yAuo/H9fn5d1SPZiHIxC794VuBuKfHOWq/tTOgor
vZ++4gCZz+Kbn0yQTJlNWF/o3UFTCibB081/Vap3j78qifupBB5CbmnR8r+iw2BtDhccS4zTB8q6
r33iIfiwOk1wTV4sTKPurc4UTrfi8lhd/wbtVYGU1c4KYFuFZEEyFJgRa+WX/FAEqrgme7jSChkF
HjH4Q/ulboAQsxvMekozGXQiUZe0FS5L/r34XDwE5IGMTSGA8OYvZslOq5FvQoWW1GOvyiLFidwg
aEgMlx8O9iNd+uJIU9EYIjfLuF+r1z04fDzpKdIwhWqoRzzjcpLDjwbZ+vo2ybkF1naPpLciNVxs
ntC4nidfHLq5MSmvgxNF/N3mxPdfthVgY6jNWun/i9s7Bgi0ffcjIwRGNCsTUqEEjApRBwvRMw2K
GSx+4bX5fv15b0mEZi4DSAIKzd9EbYpWbQjXMOPX+5jtg0u1bFny7/jyO2qNF4AO3USL3SZARVPZ
aootIL5lyu9jOmXCHLC38AscQgCx1wsSSx7+FGLXpOd3aAMYNZ+iPPWWooVib5jdi37sNMD6hF1L
/7x8FNkD+teEMIJt2d9LppTjPpa4N/+nOcb0kqH65bZInECiz2RXRDJvNQdcBgI8CYlIvZ0Fl4RP
p/06TCPquzwkOxWdL7RLk9WgN8yuvX2XfhqvYXGBF8T9UjWKyy8Ef6OxWiXJ/9RHnKdXztr7uP68
jB4Ds/C20EdYzmnWVg/tCmxgwCWostjy8118bdtPNHGAOfrnrn2Bg6c1sPT7bV8LeXbsYu7tJ3h3
3aVBfM/Mwr/ixjdSMawkox4aIQFbcfwP1Nre0q1ZyELVf9OBdt6QuyrTemmhyav1vpuTMJYVxxNF
bcNbeYpNDHgrvK/m5LT4MQ0u/XbvRsLliQys6t296TtqJXMnlUygOmF6QgIbOwP4Uizt0cWBNs4K
WKDv/xvaSdGBfVDHtbGG3iNZ8QqJVRTaD/cUNU29kzOamlGFK93+iWhkzTUK5gqcJxoN28/aH8Oq
rEAYGo5grWGPjp4z266KEAbryCEVFH4QvCGzVTAwAjP+VmI5GW9ikZA5kVEDqHFm6xb7MUzKlYx7
tK9omhBqxsDMDiJSjsRinTeYMlaj/fyFddCkTAXIaXi1rRzqio8QU8cp7oObvpP/6blyPXQssF/8
9qXE4xSUuQSC96n7+YKh1jTtJJI2VA1fdqfwX6bL/UXaYAtC1re0GDWXLzclt8DIlbompIabSwLk
/rJ8oOasRmYVbsOKlysA3BTw+iD0H46QsmKrhKocoUUOPioQp3vDwjv4cqzF2VbTzoop0qjprVtn
jch9n1SFj5A+hV2oTwBnG2MU33ZhimmiH1MXh1K+K2vHu6gkVdttu0JCoC4dpPnhHdAR88uUoyqc
Lp0JTL1V9mIwDLAxrqlK1jUTyU5q8sM/9gBV0j+YiEJDyG0EjHRW0uEnTt5tdoW6ceMdouY3pmla
Wq+cVwCVFD6GbjgWxyjooW5OIdXskDVMg1sJAU3CvO+Gbf2J0wvVenwF0CprwQq1IhanuGS/6vNO
pCQmAPnqPj5uagiZ0u4OC8A1LzGlmgGpVH8tWRs4r6/9ZCIWMWE54oQvhhVqJuLej6oZhlZ7jHBc
RAWhGrlnCXGyO6igXYl50hHicMScCDde2cKs7zbDQ4bx6dBhfpipzZExb05trVI8bvCLXscaDJph
HdJ1xHUT1GWmFf+YCrBuYgoU9rfnqYegXblAlko+zMbhZwiTnZMuQ2sTUgXcCj4NQTdNL8PVUbQ8
LQsx35uM5rJMehBnak1fZaw90/seFuVzn15IJKexoudGvnFSeF7ZWvvpelIQDTKuALuL4ZWOPnkU
vGtwdTQNf8h90s76XmVXwew3SyAqkAnxSuZOPit8Vg30ZtHXNw2IlntUqFftechCfFNqMvNLCSTM
3CR31/9Slh6/c9OTaaBy/JwO1A3XIJoqdhZeBqq5V5NZpAqd8YuYv1prsYc1LZi3xaKQXXQA74S6
geMfrmPhW6ua+0HvRNbRUIZH9QS1ovLIRDUeiYEbrxR777Qirf3GeKMccGp5TO7WMtVTYH0R+mxQ
fAVT4opHCYkjgKzhq14acuz4EnwNQjySo99Gl91dYCpvy6lBI8hBsNoj00p6A49bFTcSOTZ+Raes
BpIdHQR7Vh4vFe56ZYrt7KmgMHYtBEoaDmv6XfELJvu5v83z8pS32A0uY4CM526PEjET0xfwiFYu
kkXgPGa5bARCcZFZynFn1NEQ5r8Jn3S6EI2lrzTlrwaTTtbXxcXVySCD79bnVKf1LfLHCzE3g7BN
A/anwRJpA4kV6Vi2jgYJ5j4sK6PrqnIQt+NiI8TwFBAt2XQFB6wgnVV4KY0Xc1ZVqUBsn5B2kewg
b3jpeTY1kCbA4pR4bVSujoaNVdSsaytH6TCZNCvRWwx95JixGg7TCmdkDCKWZlcL3gvi8ohnRBC1
MyS5E0P4u0EycRDe52zzU7KPsIIXn9MX/1P1c/8nSJSjbdRImyAetXHmZMQSS+VzIN3iKdBW3ep+
r0jVlacv/XAkV/P+n9w34Oh6JB9ENFGWyD6pKp4Oo1RhJV3GTNGsNL3c087wuoWzsFQBowrbCRnx
dwaMHEPOvsxvaRVLR2/IQlS4RfSBgQm/E1hB7dNwiyXttC7GNE3oQf3I/vo3jj5PMecfFOuF3cs/
WCcmIpOEuC7uCYWZtwCS9nG7N0Z/B+jgwJ7JsDWpgWpiLA1Gg/jKAXpA5YKA/V8syPcAV4fBW+jI
emVzUwVDDC+hk4Kc3YYPmYSv5HoLaVpdNrZWkDH50WiLA64tiqb3wRFvPv8IUKZgX5yt2JOlc7za
XWR0dSlthnzwOBL/0pQLGB0cw3/FlJwKNoHpcqn4w93aakzG5/tDy5Am9RO4cWuvQtL8Sm8jP9JW
ShuaEUjXEMneFHUvJicmVkE/o0rxLX2NBFPt8XhLCGZC5uVjLI17EzTSa3JdHr+rSGhxfKUsS3dY
MOxpuKHJihjtSz1ctSmgSWGyra0IEpg5fK2oN+ztP+12FYTjkhSJdZ0X/mMlww7QRvLtL6R9fRZG
Ae7Vox9Th/iv9nDqsO3+9yDijzyQ4RLZ5BDc+yL2UNVXNmR0zO5MlHFDUKh/ZkgkipjEhiqaf45G
7ZuVn0a1CYveXQyKuzOJ8chxx/VKL43gMtYZfsDrr4iUoltuvN9VMWZ4Ouj/G6hVpXFGKUYIHl2Z
0RhX4QgRWR0EfyzHjAPR5NnDsKPb4DMaEXNXO17N8NN5BWRE0NDrcxhTxQEFdsKeTEypER2UvCEK
v6LOnG6/6vMpNfQ/QoWdFLSb+zCnaBZvloPANhHTLGVGalnLuzmJAr4iZ4B3EZKyl9a6J0Zo2l5A
hAe/MoHLQze8LFUPcEzlcSuCCqesYOHssCft047iL6W3BkEsSv+aKeMb+DlJiMzcfcTeAR0AT61J
oHGbsY+HuidsuqruAR7FESkB2SN3RRq6F9B6EFZ1b8bGQNJNxsWHmHMJy7McOLPh4ghkL6M5xJIG
i2pkzV4ZcXKUvlhKwX/gpj16HfoMkAaJCP+o+hAluMTHYIHOL1bqInomAXuUahVIIUGlFdjXph1h
Mbq2lPss1f55IJPnWfP0litobRLAXIlNPDGJ4+23hHtELLifFJtcNkdJByFSuAWtCPawzzPZo30u
pP9hwBG2igAuIA89AA8uJzOUCSDt/2xS2XnP/vE7CfR2Jnwa96ANHrWA6z1KWjFMg7Eze5Sf/gSM
VAmmRV8bylAlXDsibTcy1XyfAVCDwb/SKi0GS9S/VKd8XjvIRBmOYv0WMmOsYJV8RjTNXv9HkWqb
aXQvS2rEmdcanvEks6o9G45yi0rBUGtuYJAaIcQAB9V4F1ys7mEyOXJQ7/OW8gXGPgguFEsKXqIW
SuajRkoPvVgVm2OiMh7UDVFEgbHWz5Tc4d6kvwpf3hAnnDgVj9jE/wDDB5Zy1c3qjhE35rEpJ2/k
CGxQmFxbrmErQ6+4PEi/NNXKdI0yX+2ycXsbbl0KovnywhRQ/3PkPxto4MRaaziVVSj7A4TA+xMJ
Lfj5R/Dzs6OgMd/1Za+pe7/yBy4YgScVDAtRee6y7tadkraJy8Qym3Svf8GhriSsalRkMyUyEf9t
PS4ITUeYetmiMfUjPFTAKtxd37FnyI8HYpQHVg65bz0saawKO4JLolPTFm0SrVUQGKEZj0ulAV/V
Z2fbvayDYKHLHsp25cish58QE5LiLkdeCY6KLevXcw7WKSJzBlCG5fXCOmzWEi/RpSSzyQI1vcJL
ujhPU/SScOPXCczJGhFUdgU83jTsGFR3vv33+mP6TmOk78LNe9g0shwFfS0HsmkUDdPba0ERpD/b
7+0pm4rg2AfIHVKMmzcZoFLhjgdLzue18Hp4xcJc8E4SRQyuskWydAfKpINjOlM5n/29Jtqx2PEO
dyeorNK+DhAMsYiHvBhLolZRsIpmVN/u8mZN/945wWsxEnxKCGTB/OdwToAvUnYzc51pfa1P4CDu
dfc9tYq22u3O96KWfL23I/oi07oqKv9P3dwwCW6mj1QQCx4pIO70cvz2pX5KhlihUkJRbdGciJ90
d5q3fC9+VSu5mfbGjeas0OD0tjGI4YAZq+BX16Og09eVpm9UhC3GSwW5CyflQdflMSPj+jmbF0cS
bIsmGAEGpL63xjIEZPaFH1MYQ0bOIHAeckmKisQrVbSHssyyRrtlQf2AcuL8sM2UgG85Mz+v7eB+
TKKRzJOWcJypY0N/6PbbeDz+tyCHVNIVjYezYiAFqTlSLmMnb/WsqB3SpoxXkDD2lQApJ1xYoiTy
OpcEe1h3I/oZzL9OpajUTQ38Io50U0vCR67ZRXs1YgSYe0bOD5Sj7H4R2/5i/A0LuIX78unNBUnR
vq3EN25z1e3IY185iyYUHZMETeTf5HapVp+8k5vo8EAVapkcPG86EYTIji0PGoHI94imi2uthNbj
FIIHkQW2buTuB9dftCpRHhjHHVORm2gjgrYM7drwYah2ebg69L16wzZmeWj2ZYxSQbSD5QOkMPxR
eGmQ9oKQ4iYHRwMJruOJDMbbUy3MYBOKrByc0Nj0f89cjktlY/SSCPek9gnlk81ZoM1hxi8ytoqa
DjxMOL4vEWjeEdovAiKQnXl6d+oMsLLqLilIpOw9Zcy1HLmUNN1A1OCfClbMbxHqJPkD1LjOUNsv
obTeJrnVur9HVVes3+RgemkkBxaRUNKbwgdbpV94MIkD0DgVpzz97baAU41Insnr1L5kf9BgOM3M
j21F2ehnyTpdqB9O7DMykVVfbmJsX2VOXkzYOSBI+7HqJx6kLPLdM1xh5qJFsvowy41srDliiVVt
PCE4LDpCmlpk7kaGi30+BGyV1fiehiCd3xMjgX30lTGwRUyh8bsDY6bekUJPlQ2eDjqjtV/PO+oI
YCtzFZI6Okh8oLsllbO5oWlf0WFK5yXTQNCB2V+2JP1+soHK0EunDLUAcU3usNxOlGlCwc50ze1l
tAnFecOP7zwdWNnmyPAR0sztq58PMbGD9AHZV1bicqQqFlcq/+NZLCzedcDamA+wQcD0LxpmFU/W
lhUpNABZ7yZMd/WD7hbxsRjTMOxOtb24E+3/mqrzkZ21pBCO7gyd4WN+qeim+etdTg+3qtFpFdoC
A+aM13grXsgpe13T9MBSXzYXGZnJ9p9D/hkoaDXRgyn4YrKCqK1Fwb2NXJMBOzae/bXthLDKRICM
q8rJj/EDDsTmkAKmwOTVENrFO+7rITTyy/DrJrJ5j1C0Vj8deCQOwOjzUpSP8Qh+Nlp8eUP8XJMI
8DibgNvwIi5jJxwWr06thJD6uvkj1iMsAjNAvvuJVl69ZhUEKkbEEIzzEvCW8T9RpOFVgbdBCYsX
zcq15QFiEDc5c2xbsXDsyII4E+vGlj2M07Dt96TUZTl1Rt3L8ANiRPjuIVQuvaAtI8t0L84NpA2s
0KLgx9vUer40wfP3jrJl2HB21OI4WfhpdcW75xX7stqhsVPtEPg9l6RjvaYdj4MqQz75zTsgFGGj
3pRImojRebNT1w3OTwF52rahxK1Gsd2KdMyrQ5QEoqNpRXa6Ox6XWAdfHuW3mYZ7A04VD7Nv1gP0
xVB/LqFd3VUXWXg+wigcjg0rIOk+Z0jlIhNO2fEIcQgK0AyWiGluXYqIZoS2FcJ5R1BRg9+lg3BP
/2ar2yOLpG/BKORl3FouzjQiBBcbl1IznOisktvEYRCS39nfQXHfSkPd/t84Ll1WCaRR/whbv/JQ
CJzqymserK4CcIwJq9aAeDTSxh3iClXRbZir6geqfOgnMXtpzf1A+UuB1ue4nNa0qoOujUBjL1N2
ODztyRK7UNe8sUnquYMCljw33uDxrZBpJ8Bbo4UAiDrtfNG68iatDs/YG59AOTLHV+exq7zg153e
ISqXwYx4MHnfodVcI+EhyyGl2UUuCg9prYNRCVXMdvqj/HbxW6CUsD0CD7TWZIrwJs7NZJeGqIzW
5Ft+vpRXBa8RMZg+t0vVzs1pYyoGsXNluBNnagUVa14uGrzmh93qszshnHcALNBK0lhB5IlVfXyK
4jdYH7JDP1ewZXGaIWxIwa6TaeEsGHouyfSJsLQkIqcmYYiDhVcPnBvXa05VhpEwRSJPMB7+1Ae5
m32KG949HvIj8mMbchQHRdk58EqPkuZzfPyzlcdsybT/OGzCHdaD1Fxy3cCmQe5Qs32o/Q1QBhTN
yIjGxm4k5tg1YVqw/E+hnDSYq3yHvFLzHwfYNejpD246cbZn+UPn7N6lQ9h6Eh8tvnmYlbnKI3uz
TH47zVTwJxZSXkq9lyxpn0NFbJBZOm8I/I3w+fuXpzv9wyHWkKqNSWXrvjzK70PfSbkO2Pi4w6ay
N536KeKXRMFULh2cllW1Re+nzRB9oDaCvYutsYsA3orzx0EMvsLT7MfmRYQkg6ynyOQgHMBknjYK
IAjKAeCONQhXoF6v8DeNg8pbHHYqnxlpx9nSBTK3hrnok392lCnsDYEkPwZOhLv5FX3baaa1P+e7
DfDBbyZJgkcZd7cvH+4Jz74v74yooHuAOr4UJIkSdNEQBjIj6mCewIDGeDUjogm4i3jwHYoCSKCV
55Ypp6UPfrVWvG4BLO6ZTu6OVdCI/+CGxtiedjmnaRVa8+4veNihzQLHvYg6H8koZDaM2u9Fw1GI
O+fl+it2nEQsIPcpcRw1XmC8grazL3dMhmS3UriLNdmO6hiBl3dOjVcE/JNd2sCb004hM/oMPxgE
PN1a893z1+ZYzYWvvTXmQOpBeLNB2gTgeVY/e4j52eD5P6l1sBUCpduE//nFeG5fHSlLaZDaCxDs
CpIuoBXmz1cdrXJcX4wsCxAvUglB/tVo6KE+vKW5/aaD7Gm40NYF4sxTAm5A+JOP2d4bGWFY/vD+
ZzZWXMxucEHOEdIICJjxsKr7LSulF3VhbRmLC5S83O1vFXVr0sqJPImbJ7I6nrW99Pn478yjl55N
VzmEieFDDs46fDtL7L8usMgqz/W5jV6mjw9rB1UN07fWSwSlJaAm0wAhObL9nAP22ovdS5f5d8Va
neyMA9acg9rlI9H7b0zzRHQxqPAANmD/6H18Z9XQuJoBtSD73W6yF5604sWyQ7r6EEppZVFRFbte
OI35sIsWP3HKT0vICiAMKa2UhdFdLbjUYO0waLZUC46hJ32JEr4oKUL2FJJ3XCVKApDz/5b/C7Ve
x1tPfaY3tRNyYkkLfp64M//Tl/wviipotEispTunxQbnCAvA8OB/wtk6qQMXpKC041GzTq6y26Uh
bD1mCQ/1noUTBfETabMeZTAYUfch9vzG29X54hhFjDC5idBVG5cS85GojAIBMLgpG0EjbskSwGkw
aWpHPJPIlYT8zqRDNJbDY2qVUFfBJR9JDJxFtoz7gsdF9EVRncYJK71u9NRtiGMMu/MtfgCCviuW
/tWNHmR9oFXgAJVrMAlI566M1szDXu0+O7cjuRF46hhxg37aqK0MCwAZee2opzwsHzC4QhUiJ86Y
WQ5C79Eov0ILsb6s1ABdHKcFoBa9zB9xCUw7RSj9oKcTo05W9Q9xJgemWpL+8nerDlx8hnkKo536
bS3MElppPqS0AuFvzDiq6F4GswTdf/ppXU150qHxSchzron7eHe9q1XHxjX+xHqBhBg59hKpjCqm
GwAw+Au13GiO98gar2QBAPGJ94D3yvmN5LR8SqX1XmjQHAvLqBYaLnZZOwzxJTPnB7r4lqz5HqNg
j8zCgpJQWkJorwhMVx6XEWMphVIqwsVU3vf9XBnfpHR8G7NyGhBXkbSJbxG1ZlVm0YbajacsgeWF
NqyO7lauajhGWskt5BRGeSdqOrsLfRualQt4/UgmZq8pGbSgyS2Y6ZHbU9/DWsUJHD8Mvh9M6UOT
2q+i6km3sswp3VIvDMcvkEY+iq0sPOvjGiCfSaTbUTIBBA9Jl6UvH/Gz8iLUkiTkYqloEH6NiOqZ
hry6vWcy4U7N6TLbRwJnMr0Ke5q115p7N73WI/L6s/Jj5HXSPYeXuFn6Cu8Ob2APRFV6Ifq5pTzn
3Ca99kIL5yuS8IOVB2/hJVx6GOoDWBN85h6Yt1/39uV7lXgDZ3cNpg1Qx/30suDPyMoG6ZOzwKRJ
GKdd5ktEkWrGFmTrsKfXdiV9J+IUdVU+8NqcBcPDp5N8aC2Ui6Hq+6MEYuyJjZK3lCOHew4qFkM1
MMZa3hN+Uha3oOLzHiSGkcIYDCPukLO3lJcC7FQlP545fE3ojXJZOGV3wGaLnRUXlyZ33pW6NmIC
IZ99vDKOAV92ry3pLRJk+qhsFI/cyr1AKeFi+o1PGEr/SVxrz2b2IbCNubT08wBXGwpVuXpwNbHD
JnrA6xTCz/OVocbfUoMyQteJObr4r+ven02gtDepSQKLRjZLRdAuVfrjB8Gc32/1M144+D+jwPRp
+7w7HcXLamXpPXPs2K//JNWEwuKhk1EJhJMi3sbe6RaDme2VQ4vJSsVL+gzlOKkE8I+4jKaEt2XE
f8VjYaCC1jCvNKB2dnMTVuvBo9VH9clfLPPWmBVR56BXXYIMJSSnsRC0eNeBHIU9H8SS9EchjNRN
snov4DtnZG9PHVLXaKDuWF8La/jJDD31u/8jIWCmtpQS6Z0toxIRQCYmDEX+mPs5JsmXrxGRVge8
ektH6EMNQUT/x45UkoXj5+CuSK3Eku8Y5aRNccwhO4dukytep60aH46Syokq6WV5DxaQUWIhpUhA
BBBN86D80QgXOYoqNDOHRgIcOYuJ0R9SUbTLZmDqpSB60+RuMq/oKEITAIcH3HNbW4dn+h5xbsTM
cLeMR7vDKkXL5I3XXFkHklIDHonetrXl9m0OrS8up1xPQtw6VwZB06WdlMoByFOLJoC3Y0lEsPUT
XyVCo6IUA/va9eYff21q/2RvFuF7W1C/wroTg+ottYGFSk3lHDteQO4UYecaeqvAYA7Q7jQw40HA
agyQR75xkqJpJvxSmeLAC9K3DHe4i9jzm5jOP9drkT3ZMJZqAFDdRA+CuKOJAxb9KM1eUa8OOZZc
YF44qRB8VvBJr7D1PfGGYF6iqdrksKCZmPU1ymE+FPJcbT4Q/lCnu7aZD8QT7NYHWT2yIJjnR2Hc
LYfEBZROm4yG1NSxNHhZ4AU1LdtA6fALdwK+HA3JCWRk8EEX2Mx9E1JkW434gzYFStI7nUV7UPUS
C2emIIbOak9PrZaAp5cm9B1ORpjHj1iEpy9Zb3XmiEb8GpqDe8Z++UlW5tIFZyPthMX8J+SC3zPS
TOGAjd+WqPkqdgxm4Q1TwdafrHbfYBt+XtFWC7wFdZb9h1Qsff95QdyJn0Xc79+73S9YfYb3eC9r
G+cSH0zkqeUvN1sBLWVbsMl+OpTLVvVOJeBZyy3v4nSoagO3X1xGZV5NdPvFgY6eZmitIq+JuTSM
o6XsXRN5CTuCZ8p1dt4nXPSE5KNrjfYw76VDDkTSKiTSQmm5uraqxu8dt57ZbyXFxdS+omWoYk95
Hk91JAH6HyT8kC9/nahWXWp1ocvZ4BmplZxKDgbTs/kBaJkxoPZ3nfqcrTVUcwVNczBdvdsCPOGi
roN8klfQF2Nm4LnySfQ4eRPK4HoHJBCT235Nbp60Itk/PO5p1wPL+ht7aYYVgX1iUrgWdnfPxCp2
q5Rxt72+9SRK+wVyDAVL3WbrlhRWhvsj5+CwRyfh2LiNkXVUTn/+drCwLQD4mYdnaeyzzjGNiY4g
3MFrxqh/Xxlm4eM81mFd2a87QB7cQ+BGbiJPO8V10QiI2dby86EY7JNcBDHwfBENRx1dRocYgT4D
YSKLe1nGf1BVg5xOL8m4tAKKY+lvCeG2D7qYwvSrBT9sAwCSpazv2NJ1WIoRt+hvYsz6RkKUNQkw
+WD3oUvGGbrBHoJSMCY4kSzKD8M/L4KWVigksScv7HxS+bYbs7xKbhg1zEFDB7al+ZSz4XsdAtYu
hOjQEC3FUgzK/CQoz13OcASX85AQbgV07RL+6Jva2rOZ99ISOxJ/ieNIV+6NsgV61siYab4kLR9g
yTLCze94EsmKS/0hertZoCYdS2ysRYhBD5CJ9QT+qg9MEQmmf9nuBh/YiHcxZ1EZ5feHY8WC/kIi
HCru34o3LGokc0xkvxLq7MUT5eWZ0h0x+Vh+4KmW2NJ+UeYa6wqlhN+schWH8hXnd0rT0ThbdV0m
/FqF3jxRFW2m1HMPmwzaC55FB1ErwMTueBVHc5YyO6HbikDSUBWxme3ieh2wy6hBQ++JwdWq1tc8
/rQjoAUa41tYUkATEZzjUWXW8n0+2kbVwXdX2pHXrZSY8o3BjAVde9NIfEPEN3q9oUMRYPABGDBo
XAik2nhoNwFhkpdtBhE2UDW+6ijfVncFnYFMI20H+JhTfd1+hLZ7lh6EiMYTC0Vn/IpiJ4ATN7WH
d+6Ogl6j+0TaiydesMgsTB1pKIwG20rcOtRAaymts+eeMsa83MUdMVUBhqIb2QCA0xxxg930kexz
oEMn0z2ozYC+f1Sg3isk73CG+dcMGng9p8K8Z/OARZ66NJ8D1Vk4QN+ziPltNc8+qTq1j5Uq+vgw
vt+hqm1h1/JFFD3e4ubUINEJeoYRAt8benoAumenJi433e1Vc74oSAXhpAThvHlZ5ybaXdR05HI5
d7jI69imSP4o+gg+/wnuk7aax4CrWD3tWrU29vSgLUOiS9PxUvC6M3DQZHd/dKTuOzjjIeVFGNNl
+YBhWIILslNBQ0GZvSxT7c4UlqFIBILADCsFb9sLn7UewePcVt+9dne5QOMqNL0tqE+h0vymT1d3
cR85KgBqHOOWWtxtI1hK2ZIkoVHxKYyHJUVu1e9SsaF9x9bmx1xIsHCk/U/S3n84FXMAHKFDrxZa
SSFlvkoZSqwk8KGOtitkvRCmKlRm6ny1UhaQatq3zi31nvcqMg5j6i8fJKc8VEfjNhBLvGmpX0QI
lCE4erQbA7QTbdUfPY8DHIXtrVrutBn4OkZ3XjREiVN9YBYAOjsC+WdTkoMrz2ZlkV/ksr7aOfX6
IVYzLfPj/W9iznnqdEe5qp4sTAeTDkZLa8n+4yrlaWrYdoVeV5oepAlA34ycnORPpfQ3CviHeXVt
Gug6JFsA/28yMz6Tl31Ae11S8FPHlEAwzeKT+XHX1hg5smkZA+ORjbXSs263k0U52uLjmGDKiO00
0AvAH/UDL9Gpv+UTbgvm400wuwRZ6WAiQbVCvKmrNTLL5Jt+GFWpWa2d9zH1FFFxyRvfGhAMUcp5
L3mdZ6EtDntU1NUNrlBGhOLA/8FXS79z3i0V12a+nF1NzgZzWI371rzC+Y79911gq4O8PMRE/5hu
EmuASsyqzAuXbZkpw5KdGwr3lC9eMjP8zh9HKMMhD9wFIieogJm7yzUAIq3FvbYrIC1YbODnxZx5
O8+goqJh70ZZk4AxNf9hwqd71OPDDzWb0nkaSVrFQFA6QQ5bU9QTs5LXCvMREFYgZkww9so9bIsD
adKxj4PvkSSgb9gnckxEx9kuGVRJhTisuJauHQhW1Gyl8ifPspUKYjCdMWVoHGDbttIg5KKNaOuF
bI7MNa1wKB0uCO9sHZK9C7LbN3pA/NSWSeP0ESHgZNT52MFY2E81DMBkDyxm+DHiyJZjGTShAjL9
y1hjHLTrJQrRKMb8y+peCy0Zkt0KzBt9kTs822Zqtvo7roJFIzMdk18mHEuROCHe97ShElLI2aGT
5WxRk34Tg1uxATy8n5y+hBkpC5Ipcv1nmt2CLsnFAnJkNPB/kV1FxMEtHpPO6+Pe2fNMEuwUrJlE
TS1nse1SvmM9SZ8L8KR8pZtqtuKEjxR7vR+Do4bzfhQ8TkIWxGMOj9U+5+BEXBAmiW7lzSwKGN+P
LRmBn4OC/cxLPWAZAGUdbYDPOFMZiHqv/29E9FF5iTyLecaksaYsJXcPuKLHJbeliV6M3xwJyIHj
VUoFSiWy8xaZDuDsxZU5sL505eQ6RRkFGAyIAQSXZYuurUA5VYhfsB0llrqXATybh+3NCFg5OLOF
mt6y/yKut0DzW4nfl/2dHEqZQVc57T1EvEOF+ihuf74Oma9gmYYFl6GJo73zhzhNIdZ4V/n0xvlH
eW3cyqKQV4vzHTwuSPt4v5F20R27bIp80ffMFBZbo92kTlyiQUseK9B3Kq0WinuLZe05fQoa9rFb
RQR1x/r9QtaipOQ60JQ4DmRELHsUXmfnMde5LOaC0AdhTTq1EmMPfdDKRnJHFbtXeuAMLD3hFJKi
xkmVmcvY/NBpBRz9nZylC28KqGDFbywYXbd/Y7150kiDY2BNNYrOnQAacKlWP1jR+fNwJwGlGTdy
IFazettPI82aoXN5iu2SxuDdkzMYUnRUn1xQ+MrvP/75H8nOV8ixCH5myrjArGMQBX95psULESOB
8GtM083QnYJclI6QaMSNRQZZ4O1aJgtdLxul3zy8j6NtYHp92TvEWJfIU4Mxm1swacS+9/CrsehV
eWNMJkMne+gijMHWjKg5HaPpgt7R7JOVwAdd2NwwC4HOvjLb3bor6GfrHbpXpVwhtS7TOBAVhve7
8PZjUjPdOGKizKSKG9EdCXcDjJogxiXdthcPzlhhCbckjpZJyKSO7p/nmwd7r5SIMRQYjWOTeElq
EK6Uw1JmEYK/eZ54YRb70TYiDJosJuTwMizabM8wGMMqJJVDPri/kdYXZme8jyNgiwdDVbgObww5
7KImN30lPcsnfUil0kEdBsDVjSjIFzFHx3Skk4YekG0VxG7SRzEx08cZlOZI8bxLJndlRtwf207F
iw7XI7iyIiC8zV9cyl9KEei69gVt5YA7ZyO2cj6okcrkt7gBR32Q5XMEoF310rzsxbFGAK0sbGU9
m0C2boi3ztc2iUSDSP4YSyfpdYy90YEY05S/C1wpIyVKHJxzGsL0x5IpEr/q0MV2b2M608VUHLz8
j86WVAf4SH1w1fbdYMwq30QO3dP3nmf0B02atlc+ugIk5ozmqlLLtFZI1H5Y8yps/QUQ8uvyzAtU
Zfj9ifZ3W/QqdeLOyTgsSflG623O4/Sou78ppxyM/NmROBzDhodzK1SiSJRTATleOG1nbL34hZdy
rBds6HOFBQZDo+odDeL0CtXzrTu2SrRycFuWRNkkYuVKVUJITeRgU6FDI8l8teHTh6ryL5H4bGTp
mNIQX7i2+Fv8BHRIojCQk7RFwLeppN+kqyJ32ItlD+8KO8xIRdyjKOfvG1rnrbhAEanj63MWcv9+
njIfyCT4Y+swnBUMyahVT3nn8uhjJvvBwmR6sBOKN7cLS8wQCVZg0Ij31GK7hkjJNlrQQetbv4Ud
8rNYOmDxyDqRzzqFA5HShRINj1MsirGdo4QGTWklTcKMrAVPcmdv0W/J7FPu0+/IxeROQx+pzSj5
0lhkhE92nAhD4U1GjvgJLdi78XJE/wsGpbtpnwWlNiUiJ9pHEbvEYtKt0yFuV6kv8zTjpd/C2icR
rrZt9tGTLMnJgwhbK+Dtc9JAp7G6kGVhT+dOTEeUsXHMTB/ECsIq0btZBFdvtLT+P9ymskWiD6IR
4e7A6eFKs+iRLcuJKBpPCHTx49a5STTVmqhbq2d7tdX2XLsvlfUHTfoZq4osZzbWTjLjxeQ4wnEh
O1IY//6s6EMHkArBDljcl9yg0ZQsT51Dm0iewxjA9NUpdvI6xAVhw4syZS39qkbNbAePFt/pqRTL
6Lh+/BFyvVa6v26twZPoW5SnyFn7I39c8q/VQLFvp+48cP4o0Wy60j4voCK2qa22BiPHvNrltTEN
utPpqqSyK25JQvHGpQfM3cJdAPE7+0vj5rFw7uoX51vF4JbwA4Ae0dAgyjEa+mklsa9/YtnMCLED
FVVkE0Wi5ePVUIpx9fBlW3nUH/l5alXNTw1Je1gQlPk8fgik043bhak9lVA1IAfjADcUhY1MHFVX
09w3CCw4ZHJ1N5gNCZzwZ/5Y7j99iDejHby3y8zcbjI5Zi7LRBwExGuLMTPwNzpe1D3q4O0GzfJj
vFhTm5UHkUSjq0SOByxzbs8ruWhFPBTYGLydTX7v6NUedT++S4l3/Bz5Px008HvVnV0rWFhSax4B
QtAJ8KUn0vlml35WA6OfKajkm5wAUp3R6vWQtOa/ZEfFHIbotnZi33zLqiNDSvfnx/7EE20WZ0MU
yq98lFTnFcN5FniVDChjOgdR5LcXX9JYlNsOGsqmanu51rHFMpBREHmfWup8pWwWGqRTJm1xk3hz
sPgbuzxlhStKShGlndDrqiVcwQvk+N+7k23lt12aJPShIb94DQ/CRTvAzi23eIVbpKoBdANJS4Ux
7MtQcPEgGUJPfMumxpXiVcNc3ZbpTs5wc1H5yRJpImhwZoTCuQwzvEDQfhhkepmJKwHRn1ZefgGw
hH4g9CNifb6cTpYG1g9lVKYGn3iMQnKkzAk+y9cS1Fz2miFO0zKdaNc4qeZysPNmlnvJMFCLiYqn
jKoyUd2zT7fo6My85oDoVPVhCINAi83dknlkbAYFW4ZrjieaAWkXDNTYZTr/8khWQw0bSgp+Bxg0
TTLNxhhd2LIkwRItd5PoJwUj2UcjwzaeyLJyo6t28yniFacg7oe/Tz8idPGsRw5ZjlVr9Izt1ZQK
4/8I9DCWYgoqO2qdHUk4PWT3cuM8hFib1iSpzUcOQ4/Lt3tf8/aMVp9C5C8uebTx7xz+5qxYjEAe
amOzFbyhpA1Pf/YIh4sD8pVHan6kAVRI1YqssFJxOEvu8M/fPhHWGVrhSVrJDHnphRvFfdNLyFZ6
CQc+2NkcA8WA2wu+kH1eKAwj5lzo/N7MWu/vu6He1CfsXp4Rf3Uoi3jsiRhNaGCUflisCdoFn5he
vgs8IkaQd7/prkJsnZIiLABwL9IzfeW86Rzc3qvNcARNDgWVKgSusK59psI4FTfAlMZVDqrbYxvn
bl/9OPmRe7zKG93105DX5PA+XiO0k4OPoL6b1AYktxi9ogZR7rmAeArZsdviaxZjx1pkDsH/GWjW
8WdEop3OmlNWVT5tqrVT+FNswvLEYjgVDlNkhiKF3dmS6K3YJoz2h5bGpvBvUJCOuKYZg4IqJjYZ
T4NQW8cHf9sEOHxpexEt5jcHuAH8Od7Prxc4z2tfqtZcq0Qvh3GwC9dIi1TwNpwl2ggsopuFfZ5f
9DmldZpONZNWWyL0rT+0RvkAxvkR1/Xy6CXbDUTciEZEWV/Pj4Oay8Tky62gPj8eRAAjkc19tty/
6WTfmyAEB5aHqiz4333JYro+5cnuzKdOhexs1Wy4Wn14WSG71n6OFdNT+XT40vV9/GH7577zjaG8
YCrXoCTWGIHxmXrRRQqxkDN+fz5RpPO9k8v+uN2+LrwGW2qIqdpmjOKQdx7WyfSH76ps905ovtH7
pl3eUBOy7Qs6NoDm9BbnsVygMSFYfL2f6boVGoSM4qBA17sWyRn7ffgnpvfLRgY8KI2reniy8Gla
nZgxdf/gZf1uI+CAAYBqaAbMkGc9WGW4ceWMk7CtSpOyZLPr0EEkV3ytYaspZeieX63EQPudxDaW
mlfmY3ZTE+HG7nkRccFVpjq0UyHWzAHGuz0hgqPuiFyOSpWKNQIn5YRUP8JJTMTEsIvp4QgImJdj
viaVcX0fNyz+cJQP0+dp5gmYF5PIYa2db0sz8nxUYBqNROyH7WxqESdWmVAZpT7zqc9ZUNWgeKGF
p7ShX6Bn5oQHDYc+1c+NdPtNvkAzzfktP7kmmkDvMfcinmuUDk9y1/QJHXTDGx6W6UAHHQNWOYkr
s/HUowdEaLn4OdUYPAMAeQ0pCI3uymocVUkOltkFQJSMzLttUnmvSQTUA22ql2Fe51lcAjIXd0Yi
2groybAUfZO7L/zWFErwKwey6wUNAqQfd9AeYf+qc3w21LIQXzIb0c2akRI3Il41stON8fNBAKKf
x5Bxyg8rooalpS/HDOMayItC909y6Pwr06PnTe8SETZstGoH5jgH97PEObpCOh9H1JPH0aSeRIdm
EfmZL+WZZmsTnijYHlh6c1E1WejrUt0n4Lt92UTJp2JS0+KH4zGEPUmByWIc8mJURr68xIVI+Xh6
hVsN1byLAtEgacYMWGhwkx8JMhUnf5MdhUHaoZDAE8eswlOPGdBTCdqxJBSTb95zfrFqUygX2hKe
FJ3wdmK+rrR3T8RrEAoSV5Hs4HFtWPvxVKb236LTeGJIVUiRd3iedaHVl8cfWQsVG2DvkPMbyS/v
JpkRvlqGecqEj9kdJlTVkIiFu0PdtLwdoTBD8wXgrJYsldHc4w/yEXVfCvHUh/YEjpoAsaTnG1wS
/37z3mOX6uYrPUtBAkTDktW+1dmIRVKfuyM9L1n4e6JMgmcDZGEbaiV0lM1YzSM6eKCe9vaywZwZ
HSEPncMnf+aml0hviZuT12vXpYh1fT914xidZ+8ENyLMxtMB1g8BTK17Vr4DbsNAwVgInJ4kzaDC
TtGRdnERiCwyU+LH6Re2DllVWx/B0QX8/cV9IYihFO5PSfk005LycYNHfwt2vfQhUq4c55KmhmaZ
yPxdq0WqPe43eLl6HhrNASGn9u8gbCHUQW5E1tlEt0TM8O7YdY0+nm008lv3vwo3w/AKDCdXsV65
i/IXeVEsB8X/IQQwfGj+5enSpL7gOBDpd3s2MOOnETI+PS9wvYv6wyf6PbNniVUQCVrOIpD/Nun5
uck6j0msRYT6chhJ+JJzCng5OGVJXz+99Ne9irtsbyzoRYLJrxediiighGE7z/Sn1Ra2fpuq5qnk
8Oul+JKAr5HeZ12UgqQIF2FHw+j3QZy+3jHDUkM0Wj88Hg8S8D1+bNLycB7g/LuLPQnIwegi6mcB
1EdFwGCbG4MYUVFin2ucQV52r8S+gPi5cGJwOgkeqMcXQH3JwYiAfV5+0dxyUGUyot4uxiLHCx3y
8nrGtHkCmsZTK3OvbjutwNJX1RW1zxSZfCeCMYMcrCxHZWKREAlhJq1FP7vMj6UlZXP5ug+690wQ
/7uMn6M/+NfWA2zD+RyqdAw1RBctSiD2an0nKxj5yJeb90Qz2NFwGbv+wkTu6dDkYLX1tP++TCml
tYDgJilElE4GukTF0zweKM7iWv6CwREqI2m5kBk93PZ+UU/Y4KSOS34fx44utBnY2to70Y0CNoXQ
nQNoh7jH8FNlp3GyRp6LKrQp9zDptq1plOJXDpfpJCGWru1bL3J/eh9r3hbgjx/gxnIWMLByN/2d
yGI7n36x3hsSFjQqjtMhf/pAwN/0g1jG7Rctm00/Zq8ArzXj3wwdPAprZrnWwuCRKoELdn6uO0n4
XYqLSvjdgiVkrOZWKCZuZCiBm0XeTo4ni1HuQxLdcgHHzzLEmTgg7GwzXqQnjpC3lTsYITPwaEVd
0duRIRZ5VxCDNMN3Lr4UiyMTjoYDnvTphr0l0WiLlMBX40DEiv9nLr5xDJXn3BhELMVkhNQERj1N
NwfKegNNo7Yzt3BjrEhMhXTRFjrZTUwU10NXYoZ+L+c4faSZmydzoExXYIw8xqKCYSmoqepkDR0y
2G6xctgpDlXTn08cylqqNcOXEP57miZ3GofipjjyT7/lAtPH3IrhDhPcoFdE5G1WMRgV04mRzg2A
ZJIyDhG/tiGIPY1GxBzNB4KluOZXFcsOwNNnChDpmck6yNWDhqVID3eEjqhI0xLhQh7VqjkqGg01
2TXfDd364kTnCw+Rfr8h4OO0485ERPcs5oFTGAkqQMCt7iWlafcsCU+WUcAeM5uMuOGdsqstwXP1
WddztL8gYVx/kJMR+7svD4fCZulAfblNZ5H0qc72EVzyCFPysoq2zh7xsic3r2PMTED499YeShpy
YkfUybJBYyF0R2wpiy6D3kNVeo3+DpZIzHIqg1EmLU0elRVFtr3L0eVbEFUczqBlqUsXqtWRNqMG
eCIGwudo0coJ/MNxo5xKD3/OXbi++Y0oMtJ2TWZg0DvSgHfsDCioXu+hurbgzflxEAK9w/F3+RfN
+ytvmGIff6hMyDPRqRs/Sdhwe+4s8YYqzw6W475XM83dq2ZvEgo9xerQ+NIlYo/ES/VtHEdqnVv8
EGM1wXdSb816shRV7ECN7MmCGS84WaSS7r8jtmqUrGgVRdMmekeLaqWRD1UeRfYMySabPYwFUhJF
aI+z5hMrjCkp2PgWBXwLZdwWNSmpl0ewCy0ZGBNT1oNmxmY57E5KJub2J60EIFr2Qysr9PMdBgxb
8eedMguSryfXHLvtmi1VmI1a8h+V1zEyubm398jWEEZLcU9+Md1xgPGeRucPisn8Z2gH3GDHxd0b
SYR95Y/XgFkzmUNm/VxuBh43dkoSIUlRxulT6ptcukTbjoSlBRSH5qyQyI/8oTWX58SyfMTqgV2P
LlhUKEtKIt3CCMuasGXdQCJmMopVf7VhY+rwvFnm1bWWBOFTzsWpXFhjsZjOphyqDKcIk064TB8y
bxj3OJ33ZvfI9j6RDapeoQx5YOiiabsXaKrYllj20H5s436zJUaRNUDTPjPWZisVkO9FwWM67u7u
plCgQ2uy0bij724ZHc52ds02dnRUTC1lAoPKfFd6dxOuHKNYAXHK/khyacoDu1lHb8zLMBJayW6k
dbOMorM92NH0rKe+ndi/zSDPuxBYrTeEFJL3JB2BGMqN6lzFrpTubiYTfh9N+hUAUWp38DrLwuL8
2DjlrbysNbzEqznS7d1BCS9OUgVNI59AkYQGFusnHTsPeeJp0U0xbfzlK82/U/ZunZERC4ngXtWw
FXypRjsVb043A66rJ467t18FCXcBA+j7wKoXIqd4KEeSyt6JttvUkWu5zvvD50I2S+af59F4P7xk
rRhX8y7quKkgmcjHMrXN6BXVrXO1VYZ2X+8U/EmfC3UdhNN8nO6d30OT+ktIBGvCHgVuALaqsX6c
tCB0F6pvtM4AEOf4D05tLIk87ysLgJ8HP/4pawBfXKWi+goyjgRKMLLmtKz/O+e3lvg1wAXpllvL
WG+98PQ470r48enwr7p+bj5xOffa/u0fEmMvbIrGWo23NVf715sYYTGWCeXYPui7RWgdLEIx4dZI
DKZSJUfTn2vFO3tLmPgXYx4UvOjNvgePHMOMUaBxoff9t5RTCNIvvxonupuyA1mMRZYvQ1ZdW8jQ
+dH4/hzYce6m/7WQHkkHh2vf52Te4Tox4Hg2HvjgDicub33t3Dkkdq3HxSuOJX/cqpf/ABw5Xu1t
PneyxqEymVrIu469JWz2h62squUiWj0TL9CD/BChvxd0Nbk0XNr04e91qlKqCzLi0WHMx+L0EXrS
ysbG3MoOwhjHSl6NikkxSRPxlR6gaH+7CSHc+jiTxkXUsb/DLjjKtV5ZZQOQMFlaLz2tpgZFm+je
8238zMau/O7CTYa2VRVTUvunaU6i+nzsTFRShS2Vyh4l1+3kUQBtULuaWDd9nfRMBvPrONKJsB0y
N73VaRDFOpb1vMpTYBgM8LZJSlBLMoj+oopFNIomgS2weFAHqHwpFsVXRWq9M5VwI/bNwVc/EKDF
xm6zUx+y31U0EexIzOJ1tkhPxGpAmn2oDX/UVVI0MJ+FzBdEjc3cSl0r0Gkt+1ipHMWHmPT1vUZZ
BmBQi0lEHNEA6yAVM5QgVLkd1rAAbGGBhlCl5YsR8lpaAY+U4mFP2wzyjwm+yOP5IOmIQeTnYvE9
jnjoZSNCHLmM76LhApcvFCbZa80sErmoDQOQbXEcJmsaXT3ONZMsZnzC/bqG9YesHpBP9Qdpbs3P
3AjgSU0gPtg7y1+mG3bhtBmWEml3FNu7cGB1q6W8eK/Dhy++LMKY1dSCjVpPskTow+1GA08PmeF1
smeirhbo0uiGdRJOoCn97QF4KRn/y1VQoCk7cQeffyRGAhTlYEztqhAmftV6Y1pu7FTTr4VKZDZR
mbjc3hHWaeC3EzPX4xeINOVqQgGWoeX8PqnmO7Vk7/cfXBgkwpvpjptRY7rDZIvEuzbqjQgO42js
4MYa6z6S5aCDkK7xcCCWnv6nR+xFAkonMJdgyIWJfi2k5E4cOP5II+V15mgZgdxAqyNSDCxOY6ns
Y3jxzQ4R+TvOdLiNUJYahp1WU69Aaw23iZGPsoL0jrjoNfJdC3Z+iY7lYj2hAHBYeEESRPWDG02H
/F/vlXPvhkx/zNXSfjh7UE3X7QOLeAZWKwzsUQwqO4cQwAi9g50UTpB0z0Z2OStd7fRImOVVcCxx
uHq5nK/TqR2D2Ij+uKut2jmB03BvUgx7GlT8KNi90ziCbodMqWAn3jpfGfVjfmwmxdWJteasFJaI
mz0ss5XUa2CpP0uMBRL2LRj3Siv/kZoE6ugFicPb1hyVF8ggwvd8Dl0sFnk1LwtBaW3tL8mu7Dgb
AaBfpLqy0UVrbSq7+0Jh4rLoLE93BA7dYKxdbsCkz7ycKjs7Y7ytay36htkUYxvZd+/i4ASdM+vj
PY7Wceo1yX/iqOIaKpUsGrbUr+TRVbBqOnTrkkIjCmWd4Tlv/mOjbiBi6LK0suVDuygirdpVhf7F
IgSw6STpVDkrpyVkkw5AHYMWCj404QhJ0IqRMKP4vnUfziLLWLc3RW9ldwkY2gVuiaJl7oE1GSPf
EP2Kzow+KOjiGvg+d+YTNtonPOB74zkIZ5LwD1nG71wi4KoEvlw8TlRN79cq4Xf+wgmx7ZC4Xv0R
dZHd78MmDpgPG4SmzVgcm35jAHLiW5PIXm7B/lpSOvNLtSYlW2ZX955UulfIyq65hpxM54CXnPAi
3tE8wvc0r+RjHs6c2/aoNyVi9/zyK+lbtxMzcKyc7meyhLRhw1qgypgtfLEjVmbrgp3DOQBlh6ks
VAjCq54BV35iXbEuMcneMqdwB6JPc4krtzHgToP3LdIBJuHkhS27bPbFpAadR+bBpWsl2XiJuhpn
ivqcR9Skck5I2MEHTs4D03OcYBjCNFVHW44NSSL3AH0ZEvFcE18DGFOA+L3x5UA8+3hXB/poGkrG
jDqa43sCe+fkG0/n/O5kYCBn6nycfYOSntTyIX3gsgS225oZOXyUQO5TlzePb+Ps8+s9jtqYCJuE
fabaD6VPkxQLa+Ii9vWjJxgZj5Ad0XQn/xUkmLucF8wAw2FDInC8zsO4oyxWbcABlfEVSJRWmjuL
EGYeWn2BvEjKabJZYfkklmhVsDtIdx9BLXcKG6uZ/Y6g/H+ztNEU4Gnf6FqZfWI+evWbWEKl956f
5WLox2HJoJKdeF8DUxE3XF9TvZWipwrl0deOSEXMdPdG/4FHU579Oa+HWxmk2O4OOCZAgl6dwdUF
DmFX34gH0494+XpGH1s3WZ/XqNfKO+S81v38Nsrs0twf3vEsY9Q6eexjmuzm47gcp77+rxv+XCns
wdcVK2mHA+jdm8E+T3wQVqnjmABD2Di4A4UTIn3So7VZSH12HG6CRT8Bm5/DgbR8EUXRTwFw4Gge
i8a+2n2w3ha9ovysizlqZJIqTkOo4nlJo3RBwTBrRy1AbNZTlbeGpdeRZfZtzDDDpwKpx94kBae/
TMTaD7BYVU/CtR0LZaWAeEAK2a8cWinqv5fzDRLag2APn7FQu+JCdUTbTQ/Zc2u1s5HK+tlWteR3
aj1BhQ/HDQiTEKCoigC5T5LFxlsR+h6UJG7DujxTdI7FZwjdhYJbBY0cObz1zHkVhUFRbLE4vRnE
J65TZCumiIToi4xn5qF36Ms+t9SS142Q9oruK2npTCG5NmsteMGTtB4B96Yd6HhffYy1fr+H8d3u
+cXqL217R/TxRtFQbMkyY8Zmd6WX9SDOnzI67+U+/T6DmjF070SkxM+rpCa8K77c2RrKaJHbaQWv
CX3vD2fO+JdacPlX3G+gsU5Wlh4VCZv2xrRkS7VJAsshXw3LKAsqfk3teukqRJCjQrb44XVX1JPz
xz5jVtflMhAr9wzceGXSmmsOscB1E5GcMEsRu73GeIVknU41tRWIidTQHqzalbBA4i0Y897+GAaq
VfdigPOL/O2SeM4rYu9umLX+83mPTfdfHFpqc+lbDRkYiHSYfGS7bwsPRvagzWbjPCEPO+dyBO5E
fwXXF6sOz6tTrhU2rBi5tzYLgE07YSDRm0eqzs4lI5x+6dYuQFRF6uvGJ0zgg8gzPPJOpDtFbu5o
YOQfrE89K16yDa9nP+tRoRbz1cMKUE+fOnGMucY6EXVHbpDr1/ETABGzWSZfwcl+tEh8d9Wh8KEh
5WV7krhfpaKIfPa2LqMiwHrxKnGIQUjDjT2Hu33q2DibHB0/RTj1z4+hap/atylgJUBZoQ6JUY46
WzGpJQyxlvIsf5bb6eG8jbWq4WjlxctHkUyChEZdzTypyUFIxa55SAS2t/abCcPJ+yYr1qA3oJbN
/uhdAWNSnqVezZIZp/p5e3wCKjYPXEtn9vKhTRe9yzn5Ib4d9WA181AvcfmoDok5iqy0BLbkpJQp
D+X0LlvhR6xKgHYXtO2ZukphtoYdowaffOpMU/TcWdW0//7FZo9bzHrF9OZzZMjfivppChLS2jWa
B3uUBkNPlBSiehbN0eVaipBqq3oaIls7CmTZMkHcVwZWFTbNRmaQYu/E0B8eALpvpfNmYR6zP1vC
cP7+bWfnF8EFYyrJu+4DHUrHAOkRLyLkuJ2v3mC07krec4Cpx1pTyYMlrUHzNi13qGAkOjtyT2Md
4+tQkY+oo0zZxhZHEHBvsySbsxBedMv1UMEBYBPp2ymZ+wgO4AVXAS4mz1imqzADC9W1rQzQZlZu
kOSx55HAms3eUxAVTRwJux3TEkGNvJIfuZ/h21pjQ+KJVXZB1n4xwLu9NdxmPm6r0HWKexDn3Q3o
HqgXTskJrQHVfym0ABZpmS0Lk4vw8+2PU0Bq4hgFKn27F+IEl8nZ46cTZ9dza/J/gbMuViPfpqNT
YOSh6kkxWvzKLOV7cZhPWzrPGA0JOvn1Wd227aWvLO5Ces/e+cTPj3JhAToN8/IkWmHJ+B25FYZs
hysnfaBIVyV+TCW93iavr7+x8PttdGioh493x4jkpBtUCx6oF1b0/ILW7lfA5OMjz/JqE23n63wM
YFrUk13uQv/U5AHOqCswJ1Yic15x2GFGFaAMDZm4JOINUApbKIneHDjuLXQKWKtqAFfBj7pnZ0k8
upVJvpEwTLuAcVTSakZ7xfgNd1gY4na7EDaRKarIhuojVOdM9ZgAozU+SN+OxRE9NFBmSKYOPkK4
oev0jI1Pls00S1fc0xEmdEkyXTlvOZPYxok6otXBHfUtwN+UWfUqyhVBAR3hDIbB7F5P3+upUUz2
nwH+KOPyltglTuMGC8rPQ2KrNGNpe8Unx0sZ6QBNyDD4UMMKss6Qk6p0ktsNSfLJPX9WIUqhI9Z5
G48SBEG68Yd9v4hWRkhx1ve6qHVP/E7gQcI/CssZJU6W48xc0Zs6SKredAycgPzhzalSl/AhOs4F
sroQUCW7cMX7tmo0+Mn0NK48luFsTPkpa5Rx87zW4Z3lhEboaQ6uDlEeN4Zw7xPD1358n+teFYvn
KLW+CsffOtZIZQRY39zBlsnjIT+cX03E8n/2m7zHau/4rsRI+S0KPAiGR4nsdMX26uO+F94XUCxj
xeRomp/q7eHy8WLTCZgyzmJdM/iwouZb6S39jehAfuFXsVzz16qUy0df/aGiVqNkszmFcSTJ50Bx
K+ifdqcJo7Hm+cr3/jsjLa2lMkuObEdJqabdvs21/0EHsN2Bgbgc1jTpvfkSZGZKEq3DOoL9AFuC
AVZE9OEB7/3cCuUjqD+rGR+z2bAnv2IJNEuWxxwGmgWzU8mjUTiJpDIxkixMhZCEIsHCaoUivd20
jdOXiSXfa7bqciS6WBO2t+Xt38nH1h5NlTAJ6HblgKVVL6e7q5y7VSmgb/5yqtQFY5yJ/wyRvKK+
yXBb6voq6rngjtGSTtrnyNlGSDGkVgYUBnHMrP6sMTiimWs2Nf6KKCepuioEo47WbGqnj2dZsmGt
u3jNFkqHk3fF90EBs2fgf3qVlSB+l6l0f4Mf2u19Rc/ulilOxztxT1r2ugJ8I7l86NszFsK3jzi8
QZkHiuqE1nygwGifOkbe9lt3Uy7bUdKQq1FsmrWhzxpgU8XGD52vENT4vDqug4aajBOTzniq0ATS
VWLBIcSJjgXCto8n+xmLFt7cXWv1vzEST5MNZBXU9+AePdkGCd+qOL5/CmGzQxrgdjBrzCoJv4ev
TyGTpfk7kVU0NUNyQS7+vqCCdn/nBnSWjp2jwkSJU7brlnOjyaOeHo80cbro0B49vTDfLe09J2kK
EnOvoc5hJHzSklr+mgxQbsOD0FW9mW3Ueg4esKXwO8FHURtJwdrkZwmtq1PCjvI9swih8MgQQL99
ECs0Zc1NtJ/BEsiF5T7h7baz9YUwx90DJ3A5UzE4BvIaGgm+ZXoH7mQxblVhAFnfUV4eVUm/C4aA
u4Oov/Sl1l1G+teYv+AvcLSYH9J0q4UgF36FVG4MsocNp+0dWWjiZ9KdseewYIqlVtAzEzQjWRXe
zM7CmwEYmNguxJR3m6bZmUZwhG2/UDBEIcr6WKgJFSEQ6r90XllzOIbyKL44jcv8RWyMCaxUezXB
CuA4ijqk3IdQdOCmHvcFQDxV7Ht6c3x9dXOXHOxopH0pFQHvDTbRKVU+eRZG9BPph/5Z/Zq7mRjY
ynAk1qzx/B/SnqJtb5v7ORA+UDc5HAFKkg138FEXTsAoxds12sfxASdMVfT6EOnacipU/PKQRShx
gjk7UTbCBORn86yZLVxIC3vq8+/iVbJWWFH23K5e1ahvmP0ZxRSKcGPciv/cI17fBoTa66seDOAl
0iW2DqHJcbEI3J/yHqc8480Lh852GO1e7FFH1bJH+qScX4d100drAS2mYfSGG7rhiyH3jlZfCNj3
vDoErWYPlRzCTgWEMvLY4uoaIXuqxHFAFsdexx0XSXYrvNnrfx3A7wjRCMCgd9XDdy8WreftW6GR
6gCFwEsvcGxMdn1Hw8QnRYuGBV54W9Vi66vouqxPdxz4v13vRZsLRDTo9wV5xmo6iCWcWCAUUnik
Cii8wXC/QZ9JmwoVfqs+pfnADIFuYNzi/g03Qy5zK67LVm39JeLobQ9aiaNA4akC2xnVgzSgUfJV
0BsT3a/lG4Twga52Y1C00djJytsZlqgg8K1snac+BlTg/ml1l7neTUVgt63lcCZDD3w0QbqWEErq
SFSqU9vK7gbz1XPqsHMcYiNTSCDx8vrW0PKgB1kTuNFT8ljmLC9kdkqyO7eP54eNF4YtMJcJonH+
hTq/zpustx3f5FKCOGdAPWDjB0uRFj6Rcd/lVUWZXF6IHRLcdDJzGqY5mrc3SLWI3xfk+mK6eLYD
Qt+zWA74kuyxpeCbfIfALlTeF1XPwYulXnnJqDU+Ng4cw8nqHc/oWjQhABz+GxgwC84HoKiljleF
2JmUfLonsPRlnEfIZb1x6zigd1EjMjGkFPBjDETCzcKPb67TWOy4/1boGrefFX9TubKCNoEzWjtC
JD+ICyArxTv9Wlgbramjg5scXb61ZN6XF2t9nJv5U2RYnsPn3Eu7aiKM3q3xk7tFDqtlxT7HGGiu
p+uPHQKPHDSZQlCmW536oicMhcLvO/nvOVZH5hYHij+pXfoElGA726sRH4gX7cdcihwvTxWO+b5e
pP0BhQrs7x7ufRXC9NzhBsSRzvNBh/KmOSqotLY1bLKS/5khE3iiV9z7APA6QtwdJbzj2c0uB+HK
WmlUoQ9UeZJZlWBCTnZAKgKcHpvzWKD1rQw7pGMhvwi9KcTj1YplXFCh5YVUYFqxWVLd4enlB1mv
ZkAowLiVch1egb2Dk5q0LuZeesgEZ61qmurxi0DJ5Gnip1mjRBNp+qFO+hU8MpgQQh3wy357logQ
O4bZ79142vOaosRhRV3urhRMl8u/Kxc6n9Nf/NKf589uec04HO/YeqaaxrHi9NlTzhx0TER8ZTR0
EePXQdJoYlQZOd0AetDPHyXJ0Sgd8Z9qVbyQ3kdzhWsoaa2WoJoe521zepaZRD3MXt+fmV+Hsnn6
NRxPxGJPhZ0iy46krbyTfqJ3id4VctNhGEcIus0aPGDlwWWemGGlSLHa5YiicSWEn/SrfHxJQZNc
x1Qf4n/988XyGyHwSCMUQSF7jXt5/NyxOXUP2sSus896CFfT0gEciMDj2XdgQLpf53IO2fkPZLWv
ViuJ1+85Gh3308Y4ZrUzlu1NbaYsSF3geoc+wS7FXPguPsfR/btohk8rWWaUZD35wTYiDXNPAIYa
LGSIRP5boTe9Lgy+f25khPZvlh1asjAV0gxacsLd3Gk+FsJJOGTt9KPOqB8/oG0QRgL4QrNVvpE7
xq99MqEfq1ei/TiKndh6/5F2NkBOT3fNSx7JqT4N2aXmy2nN8qj+xXYcBtsqFeYs1Oa/5fchFf4d
wZvb5x2jFKn6CwaLtthsOPsSr7fDnyhazvwq30LT5XigmJGLtgKny8oejeVSVulO48bQUlPynIaf
yJfFvZZgVpTsqtc7SEIzudFaaQKD7aFe2xzEBw40gZb13RS0Fg8S1sEzh8QKbhJYJGPMFa3r1amh
cGvzS/gr/Xz8RVOhiIMZ1BRD/e2ONE4KHV27rSfxxXg9o+n1RpAViL/AsXVFQzDJX5oaZTAAGfjS
Hv2CGXE2++4PyfhN/KX5Pbj47kwc00DwIeTIRuhG7K5pRnwkptii2WywCHwstSqqm9iYVJYCqi9v
3ajuA5eKKz7HUE8nZEAxqtQ8CuWmmaLVHUVVgRR5e5v0q6GFfWho0f2Kq3NnH9GBZgqBo5UQGXcq
9KNkuJoWUb/V4oxr9U9XQMFm4v+5U9TqepxU6yKYfC+bnNKsMpAYi13dNuv2CSdGW3yjrENsPvJG
kP49GALiM/aOw38Qz0116JUP8WGenpIyax6gIZS8QwAu4LbpJ/yJCT6Q/swhAy3FgegV6qsok0gX
LWak5VouG/G47bDMYCEgllfU2o6hHW2rgHPcUR0Kcscl74tPJEA5nb++bgZln4aXpNXZjpOcmkvt
Okhez3OgUXK+pY4/1Lwz0PVDGQuguCc+rjG13/Nz7/YleXmrUnoCW4HmLWsoLgOjAUXoEjxsQw9B
RgrzSTjdyEI7ng4c2PbCw6BwrDrr9QVtZ+zDG2Qbe0zsVEUiCbFXm2+NIenIR9puzYZvwC4zv/2I
najb2xzYl/mRZy7+Fm4BIx23pkUEeoyvuhxVMnknwOBCOFwOie1lgCx7ownz02bGcuEaS5QCvad+
5Z5bozSACMfZRXWbHNVPC8/QbUt1Eb7X0qOFNG2rzVMCs8emN+8dTykTtF5Eae+W/maKsDS7bpwd
I82bN77aPVqL9wQqFS0ySOACOpq4FQEaGUXGJy1jVlqdANZxTWRFtX2XqKOCFqJofCZCd9o7DIkT
PMnkRYREl0PehEfh2/XoMd9DO0M62gusqzbHS0hX7hGJ7pDO0HJYFPvPWOUHD1jOuPnZs4dJHml9
2X+dAzSXbwYSw0ds/wSUBCkb5Vlt1+tadQPEgm0QirUNhMplLdsgv9Vp1k704cWlwOxxOfXiRSO5
sXVQpZMq77n/64RdWIwZ+NaETOGhFlKT0B3f+1/tziYwy57jDJwFvczk06LSsv1VJwCWei7V/dNs
C9uPw9eI7biBxDDw9uHtpcRjj5oguDzcqAZ2HNQPU/SPOWQPW6NmQMDatJeqtLY+ShMt2IO52pSz
hw5xg+DR3PX9VUysJOieRZkpZllPWn6JyZR6q54TDybknfsMFmZ93pVme7X48eBNrH86bzOhsGyO
YQTghBV2z42gjA6G662ir8t3LhGmVqJ4wmyQcur78ZOj4RjgVY+I2MQ3+r8zzjRd2K2hXY0fu8CI
KLB4KQckczwbeNq4tgWqvGldZR71mXoooHrjOscXeDQvSV014hC/evd8Rp9j8KXHBk7CNBHKqy1o
oWOaJKFSWnvnEdDQ6BsEy1Q9jnKLDQdY3SqXRaaWqkb3I3h8MDEV6/I5xzbJpKl+t4BDPD0VYcZe
GErUGKCa1tCJUwTGgAWqjtlRDxKAFdZ6ngOd0S+csOTK5PCT4Tt337eV6lUGP0R88CcTl+urZWxB
TvEo8WZbrxuB4dko3PtCD1abo2aUR61+z+zV3TF+8HOSFwM3fYALxAzYxqKsY1ecI3aUqCtozoHL
PdgC5oQiR5yb+Tk8egJu3ffg0MTuMAeo5U6I2loNa8Htmzhd1VUyegx2HHN0phJnvBKievBotysr
e3Dr9xQq5owjnfuqL8BMPGLNBfgHuO6t6xzocFCeCsTgQTrJj2WKA3dWeAR+4WVsD+4l2LK72+/R
sFXK2Lnzk/kUCVnyVDStaWzjA2dgUF6OQWQSgUhSUoUsKptQKS0VENEZkTbJ/0l//vqHyY6wOHgI
5o1Pwz+pn3FH3AwpLZA6J72G1ohK7Y/XPNddSagM/aw56bNnqqZTq+SQlt0phNuaO0Jhw/CkPKdO
T+XtomDxLTc7w0BNEe5CsvQZCq0jurB/Oppp3z96hioox5YeZm5kV7951a2wcV12hzj0OcQlE/gk
GFAi5P8tmocBby8jKAOHNepBhZ0oPMC+HpUDzFxW666MX0bGA31BMRrfrLUsmsblp+9V8L8QAJZS
DoB6Ys/IDZ/YO22KWWHL+3ToenT4Ju3zvwTGF6JNbSnWdgngm7srYnqH8Ft8NjbwSxZb8hdx5zxY
DnCzieK79vmxvpjP+zqypilKwGDrj1R5b44TXnBbgzIBEIKtrkjYe+jrWre/rbDP8EYLmKhwAhen
KFKlM06+orsXW+/bfNB54rOTkI76vycDvktR6bnJQ9PDHyXO8RXlXnD0Q9IWRn5XOdPY5Cjjk+gP
2tr+UZITlktWn92DZKRm+ZGE2aEGQQzZkB3HapNVI0H9FpZuvz1h78j09nnYxKqswLVoPpMUDu3/
iMcEvdkcq723FbDQBeI7SbxdUWxreUpoMpOs1u3CZpX8Ky7Jm8rYalXdK+JnMLPMAiIJKu4lKLA9
2m4vSlJWZ/+FFtTewf3+oHo2t3e+PgjqJDMrmd9pCY2b68qVf3WiXENSVYD97PYsXAoB53320lUE
f86Gj+DGrl1wd8ljGuSWHSoB4PgI0MMWoLpA85RcKHS6HZM127baUTQqc8FakKl5mnP/3e8TzWq3
TSmPdnk/1ecYSFoESgWAvYTcMwLNiPgo1PLLZtSYHvLXz3YoIR+mdKbaBobt1x0tG9gYkzdT7fZ/
TY908dOtU1q/lyfzuBfNsxZ9BiOsC6PJRqxUQMZhjtRB9F6GsHuz2otVC9K/eCKnFI8xR2Q7zwh0
Sm6W/WoRYHCdYgEZlFME8WtL3VZ7oaO0LzMPIJB2AtHTVvOiCVmkHSpbbAxl5gjbg+Zyzrhb3fYz
UtzcHuBMkIT6al4VlVt8+h5t0v/JOjM8rd4Wr4ObCZPsM/C42Q3lTu01Br7F9MxgOsjF3pL0vKt8
2pyG0unVjbGnPwItZbKIByW1/0KZVUEGbuN1AU843eBW1dKbauYAst/EoU7uZGIx4HfWjoEPTend
E74srT9DbQjmHBVRhXwl2csjUBunUfUHWZCD4/19L6eKmms3ZXCAaVW0j50PI3+aJ2ghfOlakQj4
yQV8xe3KPzGqkZr8vjJO4mlxSU0a/7T2zIFHO+YK0YIbEAD3kaR2qM6XzURxiVwFaQz1ZH2Wem6d
Tbqy8sN76qAYpheS/oigqjxD9xMEOHvWqreN5btPLnwqZ4wOiB40uu0GL6PPflWhoYfEcOK0Y4Sq
REjGXxqD4NdhagqqUyadpHZqAnGhRQ4kHlROYZ9Q+97M6nI9RTSiZjU78PDp8/gWxe2dBMyO0pp3
8dqhtCTEsCJEIVNXtLQ4dgTMXbSz0fTaytNqLInqJyJP6lJLk4xTCTNcj21/z4OG2F+IB8Y3tpU7
0oYvK74Mxe2kpDKWU0+yyc4dxWQwxILmTcy5SROMWUJEYhPxdK7e6baxa0HIz2LoIjWoYUFV8b4Y
vl5Ejgpu/V8qpCSuZM7l78bcjqTJmC17dPTBZfddaKE01MciZxMdu6x4edyz+1p5h8ejb6prkOP5
pN+5zffmo3ET42dEhLVnZbcTGKWatkVOgr774pfEaLx4TRrOJNX5SFZNT1mAUFmDEkq+9idls4EO
DAyK3sI+HPYaujyTRh8xehITI6gGXkRL+JG/npfY7qG9/qJgYjKaayciGz7kZQY776AqxkG6989m
iz9v77JGDR2j1A+/2Jrwz0ySXPvr0Bg6tqADi/x6rsXgV9G2jk+TW58uJdjB+3s+x/3fAKrt1gl6
F24emVEQyjY4oslP7VZFZpqF1+rnugGB+FnFqZCq69iDLElsAEdcgJ1X5a0OjuaPPA/zJk5Cwc+4
m1NQwJxf+8SFYPK1vfup+c+anyTMX1sK1XX2E8Vit/qz84T7HUpfPwSyCL3jwPnrgxt4w+ye6a0y
huUzxVKoVk75er6tI+kDSBvDkC2qJYvP9vVvtgh7cUjWx4ov1Zy8XyRQqKcdt4kCsvD0wrFy8ojx
pfX9vMtOcZFwc8K17Rh3em4Q4PaIL4az7U2grCbvECA9k0MoEcl6QsaZeyLivu1mAMvqG8S2xTry
uUpaKgB+fmw1MzDs9AP33wT9KUfZ/Ql0XE8oqqgTymXbcgdcKuAflBn1Zsbj3yBp+wUQ4w3zAr/C
jPkdmQLBU+ImhIkNhnEdnJKpJlG04eg+jgDPNYvtgfcsBb4mJwLN2w9fHuQiAu/YfFV3iZ4kY7MD
Kk41EDMPKS1zbgId9873AQ4jyTUEjDovOkIhcwf/tXKboWgnVPsQ3lwXmUIiyV882DA99f5heWXj
qqYKMMZMNkqnBxoiuVKX4SEL7SjzyfErLntgwCIUsIRVqOTZa/Aq7CNN1IY+035m2Ig2oEiIzY/M
CAER+TPmtRxr4zszZvCfaeH/WKXjKoqrrdIceVv22hK8C2UG7Q/D/1RvUnpmxm9mLFUiY6a9us4l
kbQe0POZif4yRdEeGXR2UzIE2CDj3x3HNHfvV6I8/oacbnpPwfUMUB6x96IRAs5pckj/1NDdyGDC
OsgSuMNJnJ0LAit10wsQ8YlFm+dczbtLbdBptY1LzZBDofgYu7T60WHyCe47r0bhbdgWZXdInIHn
xALtSIZsVfemS60p4j6kmtLsdUzqyntdCwfS1P6RaqEQR0+0Ag+vRFb/fC2gVtwdgvnbHNF0Fili
qTMoU8quAcY5cB9i/zbT2Ag128I9ieivBuhVMoVyTqviJH8FjO1rTp31uhREeCYHFtorLyH04UYW
1bhWLrKyTtlB1hrFszVTUqEIBvCxGk1M7EwlEYLRJyzR5BsWqxK5Fu2WQiJDFiGfteT1vdYFcU6C
55OGhDtLRSlwmQ4lLTYrBA3pK1mQb8zY1r0k2hBAA/pCqaYmVHu+7Kc0b7liM+5GLoR2i+7Cw1/k
O/yXHTkcyYyd6ZK2OwLV6XhbEHFUwxcaK4Q9rartT9NuudENBiqgOt9UmEFEZ4KEc+xH8jL5eTK3
wS0g9C/V2aKufqu2DEyCToUvYHNVmJGTisa+CwWoKiA9kSMdACDOpG6H2wl7KIkvx+MZj5hYkD+D
vmLNRr/NZZr2WvufDEIW1ZQYv04w+6tNPVBNXZxV8bjKZvHfKBdKRlLDTGc3aqksgBYneuD1W1tk
Lp3aUSkJgQMzsl8KC5bTS0YIMW15/djeyo/0n/48YqfRljP19wTQswB9EiaugJ2nJacub1+azB69
q4Qguc8REhUS3PaeIjInuauWz95nydAz5DqXWxatd7LkcCoStQ1qywuwKmfXPxWjfSFPqEU0l/wa
UJ9jbNvqzJNhpyGVZT9oHObO3/QVwtwuDJFfap02pszUy0kqe4sELQS3WiK9mT9ZALG2FUIkuplx
aumwibaadNt9IaKNRYQ1DmZ7H+iUKstXPnHcoPbm1P/+BZ8JljTZw1Qyc1//8wpusZ0SOYVIt5Jp
TjjrHn12KP5p1dtoJd4oDgCPwtCEkO7p4jWcbtZhmwOv3EQP47DCzzBies1btTkF3AvWMXcbTwxK
9enrik+o5dGk/bLWtxtFKFHh9vG4jZ0bHhz3ZnsWaFARHEmvfGA5G0+3OWuqu6RRpKvmSKcXjglj
ycJCgQ3BhUupHL70H97/kcWAoBnHgKncjGMO/gn8v+V58VFwiz5zOIZkoMj4FV2jAg9HMtYK+uoB
GW5kFdMv9ww2tpHKHT/MrjEs/pU++wjWJ1uj8pRHyGl4wTJgXdJ4rrM8iAY4AblAWcv6t7kDt8h2
Wrfq9PWXAdlcSeYXKfEggJATbGHCtpHb6/60I7sykmuXcHePrkhryrLaexYwN4EwEB8t2GMcYJ4d
/ry7gvFIJd7BrQ7OQNnZoWr0uXZgLaJY+u+aP53FCFycJE7vvxX4c6Z7/joPSpwDs2xhdX9kUGdU
ffk7clfKOHGU45AqIfSeF+Zutyzx7bK0MxSSBMPPS10PYVUJRPDyo50kPvtJc7LofkXxNcHwn8aC
rjnI1lHJ8Rod1QmLQ1xdzOinGufAfrViPrakRmW+Ibd2uPfnAQKPvv6TZHEblm+fZif6ZYrwtqVc
A5z/rMraL/o37koyL68SNnizbcLwe0uU6tIw2cAZSsCIFaRQhXgcS7KFT8scpBL2iX1Pu+D0ltc1
HchgBDg/BlcYnf+ID7CAdG4HfQJf/hzksf8qRP6ljvB6jWHrpqkYsFmHT1BiMYy0PuJSxQ/RHQSQ
gJQ5Ugorzsxf5YT1TgaIj0DeBqIXkxv0E+p1UWLQzjp5h9pcfK3IsBvvlkPHZ7ennrz+U/J733AP
xLhhMnrUBPZV0hMhUU0hbhFLGM5bGX3ZQqASUl8m7U0a7RIYnUtZUoNFDsxEybUuA6zGQd92mzNv
xb/v3Vyf5qlJrdHU2tb6CgbrudqpUFjfMI72O3MGimO7q03thv0dfbnqavWE6QeQvRezcrnAncm3
fS2nnx0uMbC3p2XL35o83EPfuYH7c9BBI5T+DvO/9xlXrM9jDZinFIx7hs2/cO66k6Yy7C0yF48u
WPVJXPf/5eohTc6G8/u9ECye/oXJl635RVi9jySO0cD/NPRA1uDH0rzeMHgPVR/fbr+TzWrxCIej
3ZyUsrBl4lE6r9I+BOPGXb+NFotEg1QO3oxHC0JoVrvjdGdzy0N7/tfRDpxHpzRjJR4PnNfbRhge
coBCF9psjIDQWfJefUfCPsfJkjlruFjl0J7nNyKMyj06uB2T7u/PZBJjHgVtsVz4LSz7Ru3RU4ej
UsFxHiymcW3/46m9pJTqETRba/ZR6iXg15iqcIW1mTPkxoHU0zRp6gsuZo81JJcVjOs+DQPQv3fr
tUfJ2nokd4ATWC3EFbNi5Dt5R7MEv6seeCrjmObfjUq5Ur7nr7viv4ve3gM/MftsFvHp19r5kG7z
Ud8udO7R1GKrFZ6sixAM4zqw4jtw2XVddYjM9QornLavLe0FpAxFt+qhJi2CG5OJbr9I2tOvO2KK
+OrY1TPRHmuRcXkhAQ5NXV618e34l7nLrgZ7UvVP64pepTjbebZbng/MV9OSoOqz0P620dV9Lgky
vTddF6E4vgBMtNNF5zcz601WfnzpEGB/2bHDudZ9u0RZCJh1F4cYNQkB2fE+95iu9EJ6Dpb/6fWy
hOT8SVe3QU4wCdoN0N05ZIsqCL5Cz7qV11Y0bbR3Wx7je8UkKTQsBGkpcQmOf5wrt4Z/wterVjSP
Dtnzo85+B1wy/rll9z1jAID5VwywgHUfYnFhxeCKVC3JIOBT0b3yDvR3Ekcvg1Iijl6I2AncN+VZ
yLoJlZBC0hYr2JiwVJvBAOW2CmSYH6Put/ndQygKTcmhpegXYp8QppHpRclODSyI+WGxzzi9opDs
5lxc3vo53KshMUSb6fdZvlaKK7KEF/fhtZF0Zm7avHvI68N+vGgpWP0dLmoFRdX+UMfUQnHKaJyz
IP5Px5+bnPVpSg2Exm1UIy+9IJ8TmI1IRC4cDemxS/wvGQUW4ExeSLZ+p7NOwRReCVwN+pPw+P46
VyssPXTGz+aesYT7SI/1WysAjAfJq6BIpwIWBDf52g+1vFoPAKrsMu2CYHitkMoc+9sE0jOsIDLx
zkz+0zMHMkalyJLX8N7IG1fZVJTqFv4yEO14nG6yCznvBEtJEhnsk/2vJOvIoqRUWwh2jzZxg254
bhRNrgzo17Yrxl1yn6iW1LJBSGH2ya/rHon+X/pAwyCTrlb4BP3swGSpJI7MaJgJolOQUJW9ApnD
tJ0KfDCTxns1qXiTi7nP1irVTrzAKrK0dhSZvKE/kJcCvmHEu2a35cDDNqjkeEJz5yQCeE9+GAHr
jEjLmhTRmKE2uZk8rc4vkbFsRqgPb14ZjM5na0kEOQPTD5s/lg+UeJgXhKoo8oTxZ7krdo204YtM
9XH65d11xoLOSCrW048nUFPjrkLVz5sZDlQUKXcN36tDfaEv7Sffith0APBSdQCVw1ytIe46Dluw
b6a3GPwVFMFfPfkjRT6GdQsnzUSMTyD9sYFYm8z8lzdjordUnTv+zUFqclHTsr+2WmrKNPrzrsAw
a6xXaXq5wf3YZxGAtsa08epksSZr6mpV4B6eRZlD+VQWu/xPwVPYfyjJht5ur2D3wDvmjyko1+tn
lzWmF3TLJceJ6TgobU1TaZg4tJ0YCPE0D4iuxcmT5d/VXGetdbtkz3dd10xEIJtE3/E3IkQ0wve6
cHPpIOvJFnxrm/x+hn8YbjInTS9UavgIohEf6bKOVPmUYzQrNUssgZloxN6KzHAIAukukaf+ijvE
EssJy8OlfBx1nn/P0wM4pyNuNFpS6FAdNlelk2OzwsqNxa2D/3MUqaxQDrCG9NwP9G4YnFwFDH8r
DH6TW/RPWQxd5ez+8ehWsp+gV97WCHpTxwhDOl7VBRgNfJ1oDwMKfTvD5R0fmCBuKwga0AtRidHX
DstqPRb5vt1i+fUHaKIgs05aQ9UHUG/LYaeNvn1hSA9Dbo5c+cP84lf2rpR0WXLbWiBZg9Dobvzf
S/12/OqAsF3DZRBb5PfLj3amMkKbNS99jPr0sglQFLx5KJglrGNIUx5rMdFy7fwTN6AFuZo/uwJq
goHTsIZSZ/EmcCcjtUdT+WnJgebymrR6JLGLkeEYSLuFVryMJvGC2ZR7aA93KkoI1pWC4bF+84HM
vSsQqz4uw768jb428gHrR+Hy8KFvWCH2MjSLhcf8ZA2lo+yNKUsy1Bow4ojPdgR1tZN4V/9e3TmU
fT2Lo9BR9Tv90gIEnGQBd5199GUyr2ksZALr/s4uHTtSbPBYHFdUv12iaouM/fYy6Isk7i/GyTic
l4dMDaQOx61uBv0FURF6ciulOWH56MJjXZO/2HDcRY4/wIulNjlFOpVybj/mzhheSaPTqC02j8Lo
ujAJJo3l0uxfd0lkoRTvjRs1lCSvSsGNl4eklhAAhScTpDjZRIykcC7FA4gF5ulo17nSs8tBaI5v
hOf7gaeQAi+RhwaklBqQxmQtrg3ccn0ycIRtuhiObaEpBLTX/PuDPu5RaO/Dqvign0TJdDx66SOv
DGfLYks/RNiQoDL8kETPQOUjWxvXguwiDDAu3qMnxJe9P90+E5FaYIbWq/JJZJJK0mRjQG0KffMj
k346gEpOfMOCvt2Y9ytwb5zdWMiO0aR2obzWZyPV6r+Gws1cNSPSuerNjO1AoB8oPYyukvuS0dXr
C9ifoYKc6QQ8AKzrzFhT1S7sLu08EN+wsH6Ie5ibDefMWkB0d6lGsa882G1e59BYPUOvlIUmxaGw
8BSQJoK9zUtsvpwZrt3WcpfBup2lItx648gQUnqB3nG/Biny20GIIYiThPo1BTmR4QKQGSh4/Vsf
VMxppKagaJRIScLTmOdZChJ8AiFsgBCfSdYQaSIGMMvpK8k1TNX1S3B/k/w4oS24iXais//96TnQ
XoJy2AKdikzUtDiN9i6Bmg7xPkv2ei4VaE7PKB+ft/VNewv1f7k5y5Tahb3nsz+QAxhNAM2six0q
0y/L8XO770+ebG51oizQIdCv8bb3is3jl9dZmI07ZDNPXSKF3URhVBVUR06UXXi7x1YdzRe/+ZGw
Tr7+rr4B3IpQsZhUWXbQlrynF7mSSD3K0cCpSmHK3kmeYPmHGf8Blmqw1/ELwftb3vanUMu8PVga
jbeErCMmnTyE29gzyrbp+d+fC6FhnxUV66zGdUyFZZOdEM7GIxjasu2ZuVy28dAj5GXRN2lvqaRn
eKA0FQIjQ2X7i8abrOGxWa1dhUdJQNcU4lagzlse1vyqf6YMhicX5W6yGkYH9uld2wF+bjjvbHTa
9DVroUkW7Y986PqdSYQmMLzx44E963OBKsY2h5f6v9j0sNLrHGE0BEmXdyzzKoqP88Y/pDv0gdMO
BOxpeSbuOBqyMrxKZ+inczLPpj+bmbH3EEKeXfKatqDxIc0Tk2lAW6Xn77m0k6ZnX3tb3kR1ayR4
kYk6YVfXHlHDVbgaqEmgne9/Be569pR+aVUkc9RgbUbXHvvDfG46U9BPXFwhf0c/lsKrmiww+dG4
cRGVpjIZ2RZnhB91/9hH2FJMl6Ig0hJaqaPquOnlfkxHU/ZcQEvejR4KZHQWMWFBg0RK74BBN21E
Yv3brcdXqn1rsV5NNfK+I0BA7gC5W4KUIbYUDADkF93g2mPbYPAQBRrrkB4RnOMhhl7VPLohIoI/
hiEedrwhnQm2E7NhyeycKaF5CzQkQ/s47VuVSfSUYKvxLxpmZ5PpNxpDd542sttymi+TBQx0DvHG
ybl7O7QDNA5r5AFplRLCFP6juVTY6R7x86s+xAImVyZylbHFHAQAfM6qNw6mRbBAelv2+avydAIN
+oYxGRcBNDWt+1jgsdSar4eXt8+yu+hdyYtv0NUF6lEQIbAeXOvDq/vJu/lzwZkR21vtMHY8xfyf
ZuMBmMGsZae9dupsgNA2C+vLWS/1EqAQsY87sBCZqMFI+omHsllA37i/xlcAsxuciVsfYMVzK5g+
+csZDytVu92m7qaIyls120mDkgABlC5ntiTPMDjLqKW/ZAkYbrlY13ZV7BF7jwW/BfezU5Zxjyz5
dqizu11bUa3dtOef10LHf7aTfv5f5cLArzgkj9zOwVXFduzDihFtBRHwLillij5PfXF6ZUbe++eZ
soHUTuImLopjkeYZxuwCPtOimjrGUw/mMdWIWb0Vo0RQASTcDQwKfH3S9Azo6sdr9NahJO/Rt0TX
wlsY0XPQ/L7S9e18DB5l3WUdBZFN4LlkeEYD+yhYMHSdwRk35VBeifPne7JI6mgbIn/vUPyMQt3L
KTVXpF/8/0b5Te9dZVg4Yfk9+3VaO6+IuAoHUdz9jh5+guUsFPWv3BiisghG8C8a0yhvFsN6JLna
Tws3Ss4YhvTUsp5OEjFv5ivbClo6iWiE7id15ec/frX1q3c+7dGHQ2xjI7l0C3b6Z4e8AAAFp4Do
0SLPzFZw+m+EbJjwpfTI0GHx76/Ls3qhgyqbiRr7Tu6tn1+CRR8g5qnvDWVXJN0jhm99i8pRWmnP
h1zlR8X+gEsrK2FnntvKmM6UQXqR9o1UgCiDjxvwf4eJOBaRqyyTwOHsCq5GZuWd5hQbKT7me7GZ
h2HKjp4zg7aYVp9wHLnNM+r5hBBp3oGGPVGhqc5Elco3XQgC2YNw9avB6wkTxoDQUkDqrpDQ9YxL
dUPNruEO4pldxFORycv/8EcmMYBjf8pLojVyxwMkpDOcRsKTQH2+uVeNtiFzIkZl2C3uwhQEffjY
zUhKp397RI0eEEpdKdneCI9uSFtDwhSGBwN7xRd9GQKUzUvetU7UfD18A+nQ1jAGqLOBOLChBId3
PcUwQgDeC5feTzad38iqLQD1Kfzxf1a7uJXvXf84YyAE910UpnOA1bL4oZD+x3Y6zM3eYGTxkxET
mTwgwuGr95cfrcyqI/r6Vh6wFO3jm+pth3pMWOnoe7J4b0Kmcgu6exKJOr8pkuQhAoE1iCXeIts+
SJ3Rz6nNmWSl6pBrh+5S22duqpyKnkOkZo3EGyVLCpb8LlUyVPkw7T674gVs8F0UkQEgApLrggIF
ABwUjGJl7Kc81TpskkWAk4BHCJxDer2DpUY99TlLClWV5p7HpLJuuEjt6WZ/dZUxM7lTp7D4P+m1
ZflTt5iiiA81D3S65hlHj3NSOwK9Tjg7Yyg2UNQEzalMCWYLAgtAVpzAClUi4mHEkpxAgLK/y1FJ
FyRZlmM3imT5p20cT5YPlL7B6od2nAlLKcoZ5V/HfnIzfj8NeVqyhONVfrRV3v6RbTlhWcqQSjaQ
YnLy+n1BT02mTDaD588+Fx2Ijc3Bdxu1V2MjfazSDoshhfav3Cn6GmiI91nzcKMQf+dSo5gqK82K
sOJyKdJInXx+ZavntaQ5edCOpo+lh8tCmW0WlGHHAbddYCknOJ9g2LsBfE9/Ur5marGxQx6FjVfB
zIhVMYYwbkt2Mq+3N9JeEYSUuxRCgGpncuS4pp2svrdEWtpjjh/qeg8ns/03gZN9zHt4dI86sLCE
Rv9AhrlY2b839u/5VEbvD2fMG1QZcCSEyxhV+oFu2jB6no/MasOClrO2e+/Pd4eDwhAFm3kVB3Js
qMuMRe36KZmUCnxws0JnhnDqGFrYTAUbiyPIkyBc6V/K/v3lqRg0QYRfkSJf5BXCAqqneuz5xqp+
qoes0zdNZw3AQBf5MSWtrIwpmAgGEtI98p1E3hbulUeoZFe2XLsaGLMbZWJN2eNzFyJHpO9pb2fX
CdH3qybe4DVTDIzcT5PxKnrxiFODWbDJoEv+fnQv/a4f5BYQkMuwlBYqBwBhic97/iBEA8uybhJn
0H4VZ7iyLCEnBhwuDNZdE5V+gC0j/E7GOZSFwNT7cb12oeRSVJblm/kqA5168z6N/tuD/6am6Ecw
aooLgc+DyyO73mJJ9ZCj0sJ5ArnQQ1QdQbMqzoJFubHKMH5qk+Z/QeQFWjmHqfMEeECMWrxVUqih
P44jOMqptXTTAOA/3Lj1K6urt1g555bsMUbnDd/7RsJ6MhZmF57/lrjFuXUchAwHySKwAA9L7dvt
HOYX7oNGiwn8GCNASdV6J3yQD056+fxT5NbDfKdoDgiS1X8WbMXdZamM4FLYhE1DbaB6hBJYcv8m
rlB0sEZYGg3DuNxuqVz+gR2pn1tDHPris1XUVUjksGjzCOJpncu0Ooup6AZXopeV21xX2nIt4Zp9
V6XYnYZEvHgtYLvToMdgg32w1oSl08vV6wtpOEqYzySDdy8zLycQfPlJKNn06/feaWT8bmiYsV5B
grvDJu13kX3HxAKO0k4JJIWBWgDzGv4RUyOkbCBm0oeNkobT0HCe9ICQtdjKdALLeaQsEkImypYA
mQiyHz88gZRGrJTO01YUOuxY+/T234oQcQRJ1pano340NurZ7xNoVzZv+RgpvAj5f8qNG6D0hrWS
hl1m3zizyu00zvgnZuiE3PLNQVgm1rz9EbfU4+5CXi1ug/RQJH7hIap1jl3CXAoRQs6teMrCv/rU
yXOS9Ul/5k1fSiEluum9Ye7GwZQ2R/RjuZtNuqfRceywvp7b2sPtY1QmgvAQsqU5vDahgoEaGSkr
qtOTtR7G/CMfwanlOhNJ/4gz/+5Ta0DdpwaQzNZxV/GssaAfDrv2+bYiyi2vQZ8L6foXWEYhq1Ov
U9cMzxvPNEHHR/TzxwU9lUJUWrlegjU1Zb4hT3VYnUi3f05MBxaVow4tGKY81r+M8Au1SmEPmnl/
a1T1mBMKbAUPFNTLEmFsMoQP55abOPI4vr5DCKoHM35k8JKYYzgHf418wsInha12illl5THYDxbL
iufnOrEe70YP9dOXvvVh0i5W0UTunifpQ1y6x7QBoIju0y47H3nNwDEmrUiUR4pit2V47qR5t1zg
0Z+pubRy85E+pQQfYtd/UPeWLsvXQiNdBdb2sFQLpO6VFGn/ETu8yOo9S7bCJ7f8DX2/pl70WMgf
r3RkBzwmMeczKUZsOLzVOdPtKWKBA5fzM0ldoy7JgPInCUcPSh8ICr8xoLVyi+ahwfmD4EYf3o5G
T+ETO5oyqyKOiSTynL3i4TMiJc9KRMFKibnxrMLtLmQAY9buRKDgMB2cROhwbyhfSdeGyj6xmijS
0sePH2PpMM2qUSAkJBcDrVqgUQCNi1WOb/zSiiYzpM21MObKondAeV6/J4iVrE4/KZkhJaeO0UsI
CiSzqphScKKm0VKIJg78KAkidxvjMwDdwU6sXrhcrzyvXMn6pot/fLiP7TFE4emfSBIrJrk5CN0p
5jq79KxoERJssELobLTUF21kM8mYqfNpdBxpPHCozb49pnnq5Yw7o+7e6KuUKmxeFQDB/mwbe7ZE
57WuPB8ZRBz3iEbF+7hl2Pon8fGcZJpifLlg6HlCG4MUI8lCGzPg9LUH75NpVmMlGg+obKuzffGa
x71ux743MoFmw2WhoGrXURfnUkeDhQPlqjQCwr18lbfR6K3H3wocF7JWlNhkZPlj5/AZvu4r5jsk
kMSEeGKj6yY+YZ/Czf+OsUM7QbLbBuUdu9Bj8GFG+uXPkI5ukKNl45oaiGL2synZhoiSxG2/K/q3
nPA5wdsEJ8Q46I4XL5jAXltG/VcquimGt8xLI0v9Tw2KwfVQnr3H/lZ07LKQqzinZrLYO2gLyC2w
gYWSSzRo50O23Fo8zluJuA97T6ier7PWJOCZR02ZtUlVy8LqFMrqdwv8eBVqiWQ7KiDGnU/vi9PB
bJlzakLEpG2dYNhqlk7eHnaDHjQ7zXENoYwFcYExjfMgVmEWLRawWTdFpCKJY9RtGSiM0C1mnJBJ
v4tdeMXgKW5ETwyVNy12REACoW2PxzwIUfsw9J+GHUaYFi9ENC6glQ9wK2UNQQxyD00anyNSeKdA
6e2WzKiO45zBvT7YHcvdAdCAeqyzVvKrhznkgjBrBvW0ygqGXM1EQ2H8CJnVnV5hpw7n5Ma64QBH
gc6DGxq5dfNYLDeIC7sKRLDxp7an3i19iuekgWvwLsUcFYTD9VOFRhS+uX1vAJPhOstbU3fVPkv6
DSygsQ3qysE1OyXTa0QQtq3VYGYudErLvd38dV6NdYCt4lTYT11d6o2riucjOurqLgCJN3CHqx9z
qbkOEnneuR5VkOp5dfQyHvvTMc8kKCy4tiVsx/6ZnKCZC/aR3S/RNMODofrbt2s0fEri1Az8apKz
FZ9jYpB0mkwn6wNWtvNdW6x+O/AX1qjvXxg1KZvFpoZZZdcgJr9qht2sAn1W8VbfgBdAkq6y3M4n
GMro57lfRgB05dYULC8TEqyELT6gO/O+GHHpxsIYY6hb2jb15MDK0Qdc3vij6M+cjqD2B7igaQji
5P9y4T1zZSqAHw7dIeMiKaheBuxDO+YsrRD/GwCpvu+Cn8AEmJUcTegBUv5fAV7ABlkBRgKvyhX2
Ie7oVFaak1Nnazbth7Qv9X5aFe6IIwqCE90PlSw2QnhAN8U+6WfuWe8emcyFoUj9o8VbOwc/oIjS
rFjAsGR4eZx2R5a1kWZlSemf1CSYoL/j7XqILrho6FA6IVStyHSve9xIyWKa+S4Z10rxldLbjG7w
2zaZQVyfljG/azedM4g0w5Qfd0ylha5QmrloI1TA0TP4PK5NlrMsJ8+bjYs8Osi24F5LyjwttyG4
HLXWSE9U1rktZbKRtcsFH/NPuOoLL+n1DK0nNM5gIL2z9WE9ZAg/QxHWFdIoLXBIPZRCrOtvieFV
MpdlQ8abmfm7W3858hgQboMva+6kwvuw2Kvx0LIl2LT/yavJaiSgryEZ3c3V36ngwW83F3vihp/c
Bf3FBl7xYEqHV9Kfrxad5WUPobVeQ+EnfS6CgHJqH6Bir3outJlewgJaG8Z2OZcjyqMBNvbdRRgA
gl6mvC79He2dbWcOAHRcLEJdJkd2PEow6bWOKEAYd3xc9SWR8EyTBe0cFpVDmDJm5gX10i+Kn2K+
r0Y2l3JT28Y/iqZlppdszr4QpaheaXPFqBbTwyu4m4vpCYFVS36uHGPdkEkEUJ/IA4rETfwIF6Gf
N77cyt3jOIbgi2aYImBNWB3ADkG8acTfaabuGXcBhxKZQR6SV8Czkn8r6b/QWnIm0kxljs8uhegg
keODBfdMm6fqTiSKFXIw9Ir2uOEWYlerdbSuChqikttnXGLoQwOxTzYeK6duZvP2qDfHK7H5nw7T
ryEU4DVYHGNAR4Ss9wKM9S/e2Bd1E1cbrw+9UtvVs6EQwASJvvAU4DQHa70EtIHHOjJDGX561hIj
61AqUrhL/SjO2tUPTNkbYUYbjEDA+dPmf10w1KRh1cEncErPEtSWkgdM1e/BaKyrcX4Rf6tcm5T7
ZH3xjt3LhKBCFZAvwA1IEI3c3QW5W3GYMBeNTvS5KcQfp+wzKBQPV8j9chJtJPEHo/RpPhEXpoj6
5B5Z3nzxNyf+yXHTZTvs6Fg1wFWHmw57jrHreJ90QJrq0tLuTljjUJcpYl+GK0HApl8GnEQAy79e
tMZuvzQop/rIb2ELfUEvivsz1mRRV9J75IlB3yOciWWzT1pEIdVizJahawJ4C0j8CuW43lSyyBIp
k8cEVUt7NuyjQ7vZq4F0+ff+wMCcYctWzSc98kAvLMLR3kvpvDL5oiP5JPWqomniBqGKCqbvQFXO
vEWi+u/DqwRcN8ykmKEnk9cwUgORxGm2b4H0djHyl4WBL4RP5sQSAnlLEu2IKXzrQWB2to+ateZx
gfjI3kdzN/5dbcqQ39TFvvWnUN1eVKxpJJzEJhPFkflJifS9qc5ghdlOL5CsPPTIm3ZjdFu8STyt
zKaNJiX6xpX+b/3+AmnZlhuxr4cWx7t6q80NcMVyZrpGJlImfkc3n5csoBG3h7qkquVpewyYSBS0
UUgX9rjOag96d2TukGFxkqdZdYfSniztJFkFhEe4DQ1q290atdIcGhf4i/JG/NY1qQbZ2B2dxzlh
0VvKjifcWYEDvimG94CwE1C5WiFhXh6BcODP4Zhi/avb2jjJAvwanP1VrH4IZ/wkR7OW98Q78JJx
gftXBu1Sa1QuUecqQPZK+dIPUhiD1H5xFEh5y72IvWBf1FD96Atm5OKMuoXpo5dgRlwgpalrywBI
xiN+HS5XAAciTPeK6bJ9nDxaKsX4N6RbEQ4DOiWS4ayWdNpgVO41RApnURfHXmo3mDwxPfg9rP8t
uEeHXVGEgWLqAMfzGbfJe12IAVTEhgnMUhNUIl5WO+g+FvEsVE4In8N5X236YngTgHAbqnrdPxW5
TmejTJz8TJ11DdYT8QLU6nhNn130W8oE/3KySzxT7qS/XdFtTM0DdjlmyjC1hYStXocMpSMzb+a9
JO1azKezlJVo5wRz/VYD0wHCKqVdBc06eGSfN1unAYLjTBodPd2wwyamU9HAQRTKRX/S34MlfUax
+QQfNARvKe4ByvWsiqUD7h/bTEd3vF0i3ifeQJKe5GJgHBC9vShgej8wI1r0xt+YUa5aAW9ZaMS0
LSA4BM1DF4VS443xplyMGDvjvndx5ySQZVZQ7bmhK11SAdOvQbMnedQTKnd8lVgo8L3XiOA5NrkJ
wxYKQcJd4GTrOh6BDqpqo0Try6na1DyH1dPrlcmjoINeAt5NwdxBy9S51cCiLyOa5cSkzQ4RSY7R
TSB4TNrdHZJqnS40Fvr/TP7Qv32/P7xw8tygZgJJJT1V04aTqIxMGHW/rCzF7jtcGUERBf+v58di
vxQNZLTB5aelljjJSkzgWD9bR3aY7c0VONvZztvEF2SANnS8ImrlpIiERtA0TngUvvGhGQhugq6w
KhssarjTVg2cDWX9JAfRdeBo0dCTTXQsEVbpar+ejJgehgESuTkcqbA3OQsO4EDQIOk/MEmlf4Tq
TPTpUbdgsyclPHuAmRPMU1WbJ5gKVqb8o3r1TQp5dXBrOB87Zp7/SWuEgM0eu1bIHUEdNN5HSSf1
6TXbFCTE8zIN2O2olodKiL5f6pdYMMoH3H3DVP7++5Lff7uG1M7+WMQovsMRxXNPpEdB9BCJ3Qqk
TdlBX8cAIsxFgJb24IiGJMCO8iuq9vmH6rpt+PSpBbywgxJQ8nD9I3kqkkcSKrdDn3VhvJu8KcXx
h/19kwFAxZTIvHyTz8ObVGGa/TSwryLjVo8sLwX0oBX1LiVhY+Y6PDLbMrclLxQ5ZVX9kDvY2tnY
+l0IMfrRSZcpbmpycy0F6LgVxU1D3Io/sKYxel85dEa3dEdV8fsiDrPejdOgy+cd7PtRnYcXLgvG
b5Z2xFzYRRX3sZy1WTL6M2T7gEMDndOdj5gpUkUfIGIVDkZA1XHasfi2tN4gaicSGUHu1CzVLeWR
fUxkIL/AycLzm5A9kLd8KRVz+802YfTlOynxh4tG3SWdiyrvOS/SHy3MzvU7WKvvHoFMsqm9XFjF
yNwVWo5A/5+68nGuCCJgXDdFZiii2b/XLxvUX/QQTbX4o44XyjZjLco9R/HRoCAxAROeWUNlgWSa
gPCbKvQPwrKKSiMJEeiKKqbXzJaitqOY5kd1PwBdboLe8gOFSO/KMdJlcaVFZUIDtA8WgCluPH6B
etarm9YWXVUzWUm46+iHh1nkhNO1kdV9AgWvAMYnnk4DyG4tyG/Z8MFHCeGLNkpO3LV4MnaKVK4e
kQbR+gcLiYbyaAvY5Uku6n5ueJ/zRNU2WRZlkqQIAjws8rS6eMhbCkpDniBPApmdhOkVYxo+Zvyo
hFtjBvoLIukufYFD17eNkJAanM4RqbSCaa9oJ3TOUvBJ5WuXDEdiB28LEYLZlWifVkqlQrv4kKNT
jOKnuMoztNCKUD54g1u2zK4aQAbAYgWmPypY50v+aKyrb23mAXc4TPzVhByYu9D6jjHy4Wu1veV/
uEfWouO807VYAyTQdY8TDopRzvUZnPKmOJvIWmd4v3PfJH2MvektSCoJ2I6Y146qOEviohSxi9JM
hYsKvLRu/y48tmNUfjkiSIKakgPTVZMoNeTU0iKV03MA+3fCY8uQTGQybgr1QXqhTY8ULRJMfST7
a1wnTiVOYRk5I2Qu3JhpgpLvrbIu1MfwXg2uSnSUr58AaT8LEGQYfkH7JqgQuaNgPiR4v5AIQkR1
Vm00+oixbtBNBX7ijqVatTtPpJRkViyss/kUGDEuovMG8YMK5XBzHHpv5dOyBfttyP17apN3TKO4
n/3PrikI6fc+NJrLx5PGD5NzxfmeEPolayKI9nGmNvAblgixbqX/x8VGzg++fdc4+O8wSPXm6Ymg
z33e8JDO8E4Dp3oXT8Pr1DXr4TPiQeaJ3xkNiPUH7vShUyv2lCnF8F7Nybyd/Kd7UacTVTc0YgHo
ja9zaUz57chijpRqeDge88frnaIb1wdDyOiYpIYpe02LcD4dpkQNHDBWj9ZaD9DNl5HWOKdXsOsK
0J4mrnGpra7XmI+AEoQ1h2QcVWCtx02zJPBthlTi1HmQCU+okenvnJwbVgufKl+kmceHFR9xxS6v
J+GusGXXX6ysmlWULL7XvTTnYvQOqqo1WqDb6eMEbAX9HiWQkGCs9bKCD+K7ayPrsBKAMIngb+hC
RTyafqAKGMzcDsTKK2Y/3YJrQK95SAODKt3GMMuI+Urm1AJemzL3bogysAuod3GpskDr2PVFJZvX
djY+QrwD12uZqcPRfoK7q80c1v5GFYgqu676ZOXOoS3U1GftJVc49aoVvrIg9CJRYbvm1mUYeAED
LlffUqI9aHxUDxJ1b9QsALQVUsTlmQuIkBQMlx4p7pNoHsoxp6y2gg+1v19T6shCSW64s2UQudxz
0nL0UnQ1U5Eg8+RFvE7qBxBa0BTv8hcNaXyEUYpzbfUle0ek/hNfU9YKInNBuWumLzgAQtLnJIqj
lzR1TIim7MkR3R9WpZLfiNX7ygw92qQzWbKVKMX3rbHvYR5O5a1oGO+Iv98v4sagM0VDcAcViAw8
BxG7oXUsKo9xgRspLQejh2oq2SG+9wHGU3sMyXJ9cLtMQ2vXXC4adJbaR9bDd8qdMNuNkae8+JW1
4BnX1bDky7IhvX2AbS94A/fqPA+8XGaxUVE1TGZFcTW5mDVC/3AMKQRFyY+SoK5pFoI34GTJ/4aT
EqYKpBjFMvfpeHmlDE+liPdYSZ0Q7tPSaPS0LN+GqYWsLYQ5DyWTl6enTl72D71JmXSkPhKiZNDV
OYp7sEj3sxyV7o7KcT3hSFEL8k5xxfDkEu0KWV8Fflx8Ogvw4/iET3vXuY2kRH4ekcbuLZaIqHcw
oho5jwrkGMoJ4zj682YvQ8dgTqRmqr6AT/fVQZvjDFMdsmY25YII74jgHpxE0L83O80J02nCEx66
t7LlXngmatxMP/byHACYB7MzeFgxmqbpnerkUPWdA9moC7NCWo5D/V9Mi5zXrEnnYVC1hkHyvn1f
ChuGqbVu1Ji8u3zxLhqgTf2B53YOE4MFj3vzrrm8yuswmY7qI9kfu+Xb8H437rOZ4sIdhfrfQeFi
5EVXw/kMciK/74oLTGm++Xrga33zMPCXtA84G37mC983VUSFugs8Dunlue+lQpF5mPICTuSoSxYi
PxFzj0O3p1HGQZFBBGBhkRSbwvIy0DXTIfUDmJuNqeoAksr/dM2bwtZURWpA3ggb+OiWduNSr0k+
qOtbxSwQ734Dg/n3krkD/CD3Z4mPXJN3QIxp3xg7iCqEVTj+Adzlw9Lj7nb0b6IxV+O4U6BksRzD
+FkSrY5Kb7Byz9itV9ah1lGvY7ltz7/qd3L41pxPXRUJIARd9cG/IGBemP0Q63KqtwzJvbp+RrG4
LbgSCd0mlZ79M1zRpHJ85rENT/XKNgXd9yyAXGWsAoGpBnaxS77wxN1v7cBRLXiOl315qLy2JzPc
KhAk0HThEVdNGXXX3eEbfr7fkw4MtaaXs8faAN6xdQcc6FJX76Kp9RvbUrUIylP36FeEQu6qGwd6
y/5echF70txMwQLCd1A4FR46QYo/c8g/oOAxS1aTSuEpQs1EbBTlWld64SKd5L2z3UE8jKsLry6P
NL+1H9x27/Tm2IZjIHf8RveuAdxaVLWfvzRndfmE06p9HTC4U9gdJELc3IUnHfG3isIJogkxTB76
bz09CC0Ss76dMjb0fclr60gvGCLmHf4BrrlAtf9oIOssV/0qAglbfnZWleDv1GDYgAEV4nsQdeze
g+4cjHLONZcKdSwqDlfLu31dMIMNt12PlK654t3d3OO8y2HgMbWdGxdANcSCDcp/6xRniZwToDDu
/nT0a6s8bcr/o/cDGMkoua4MmFSGgk3HRdWABc3p2V14a7XBlHqwOn42DKJ+1ZiUwePIWULzt6j3
APYBhkv0WGBXc0e9acAqSHlK67i+S/p2WuOFmATZBB8wIJy06aFKIHr5kLO1ZLY3ADVWM7ng3foq
uHwUFjA/rZGhiswA6HhYP3o/+XwuGI/DgJaXvxYnnXJMWEdPvR71f+bU2CjeZ1EldNY0ayIu5gOR
IIwHSfvhs5BNOybkSkIu/O3RSVPNbWipitl7OmeWEz+liQkBLcRtVK6xJtfLTzmFVlMSIJPLCG0t
VSUitq0NeXeqlbejVEam8OuquFNThpxO6gUrF3lpJV2xc+rndX1s4TKjKXVqQHjMCoU9YsYmHIE8
q9/UfzMH2mbvjn9k2aj24tus6WNtbJtqeQQ0v4eH5Pcet8WOW5lZo/87LQCeucxp4rwHrZUGJeWu
PdxZ/VT45Fa/vDe0L3YZWlIDGpT0OASxmhZ+m35b5DwfP2170XdSlyn5gEl0w18h4QDx/qOluoY8
6o1JXl+8pMGOdpTxnetZcmUtq4BvzoaCS5ivaGrSRGCHWF1KfZWTFJa068V+kkEcN/MlWUm4qdhc
FhuxuSM+HYigiu/QEJTCc0znyWVpXSg1JeW3JmyMFTnT+uYRXOxw5d/9glkYNpaLK+fWfmYejYN6
obaK/X23j3oyU12Wzzn1eAmXJ4isYSBXk2cW/urscPv7YzwTijMqA+k5VDV0RpGlrbOPRk96H5vV
RrxrPP3aPAqKgLYYOe26ZQao/oQ26PxXx9sMrQpCiXtExjGPBlhjDAMS1SbUSNzTtTrXc5B4VKuA
KYFWMcgc04s+7b4+y2EYCgxcABRRRUJjhfZEfZnDtFUfDSayOZ6IT4JXlvYaPrwSGwSUTYivNVL8
e2jRoC2rk3ZJ6xd6NVPuAEVN7qBqmY7cSj036mRD8CWf1Ei68XFTpmL82wHUaG5Gn/aqGhIinIh+
kGCnBi6YK890/tkKsZuqp7mGEAZrD0H9CDkmfxDOnLa4KfzA5H3BEZS9du64RdWujx4dfFmYAyCq
mDt2sUKIQZJJkeD+YKbYJaU2qkVRs+6ts0CXpj8Lywf82aONSn/MVK6Llnnqa1NkDkyGga+b/k8R
VBh+K5DCBbOCyTD0t9r97EjAE7iL++rXpJNwi3nX8UWELwNyE8n09dG0l6LPus/xKjUz7DtJ+zQE
H6U/rEhf+npgjILCuE4yI+imHQfI312eMeUB40DEy+uNOZztGQ61cixcVdSQDRmdXv0ta9dY31nw
P+ay4/JWBiKN9Txb4YDpOeqzHvEyA9czKzzcICVumYu23S34c1PAikMBmuNtso34drr5/vVZJCXG
hPy7A/TS0fVqiwN23sNSh7P7pJhMKTFrmkLMUItZGu6FaZWDtFXvz7D+utnKc1OawlAI5Q/26//9
5HidIDoohbLK4h5O01a0bL9b0VZS+OKwkKhW95MBFcqSFdgffT34PsOk0kq3XnRC8hNP27XjBzIM
1WbsHooDFAYb1+HAtTEQSs3jMPlplN0urewHDNsFrHtP9wLTacYS3MylzBJRNcDg4mlMJ6ntkrel
77sl28qYpFHGawLvHEBzmhJnxdKIAmDlkgxO7b/OcYekW1ZheempnTVtwBuLDm1b2zycJw9Rw/5+
hOdUcwFKnYjlJwUdq6xBWwO2zLrWjavc5usR13udclUXWxTpM+XDymVLNt3eylnhNAo4vHFLUL81
erxodVF+DxSRvJd5vCGVNynlQNBS0z6UBf+5z6ypYDO15xEQ9Tfcrhi2XDVx1EhC/Px2gaB8szKl
4InYWqI/SkS84u7KHHzzQ9dZaRRGMSgEA7aU8dNmzfL4P+nPDzcMD+u8dcQZMHoLBHl0l4cuwv8a
vXSiWi5LRcMlVUqJtib4iD/ZKKHpvJO+IUxWaat7O1c4wHMvQZSqYYTEG11IutXRyHWTlb283A/2
d57/eq3p900xP3S0yHoll4Qaz/tWtK5A2/XcFbhfwBTOTvxeI5kU2Tgi9TpPXhRm6lt1O+MOQfR6
Ac3IRw8fwi47NuadtmnwA9g9J9RDKmiTNuH47jCuQDWjhvTeGVxFWjRJBD6Zoi64aBUEuEjXVu7x
8wFwOvCDl2haI2JpdjL0fW7GRNiNWkgStaf1rIhSoWL9Ioa1THLPPX8bHqm3NCevE3Hm/i69Xy8F
pEijF1k+wJz0Xy2bfveQ7fdFh6dTgeTcR9907HPUJAnH1rOWGalEyfOrNZFGtDnEr46vcDLJLFV2
QHyMi3mzuPCmrRL76/Z2LyyfyC+6qX+auWhi0sP04tysZzdI/oaMy+6YMe2iWPaaOqRz06waG7rP
zjZJQKdtNeDcIcuVkcMJv9goNcpNbImrGE0M1DZ8TEYMWsL9549d2g80FLOFDGYAvBKpAFEam4ei
zbs1n8BgeLHF05/9kBh7yREiS8S2U6mM4yDCq9FGwERnJC5C+IDs7Yj+qltWE5ZN/livT7ahx08f
GVDC7zMuBgC52wz7pnyYEM3X6hwoh9tJOwNJ+gb5rlIKbh9qXTDxhFG/5r9f88cijkxFr1XMpCLA
oOr/Raxy5DWg2wTD/pdowtE5aNexniBZTImtJI3T5M1h3tAoyZv2TyE9QLMEoQ1y2EiRAZNbcyi9
EHr1IWeua/ukm/c7jiIczjPo1Wt4RmhpVejUzG1X9GtLbSrIrCgk49y8u9qOP8dzdxUUcNN7GNoN
D9SaVVDRViIZLn+8o0s6Dn8QqBRWIwMvrg9TrjUnHYMCDSq14irYThGvt06+bjKcsd/7/ymQvvPn
YXd0V11URTKHNM2fiGmk8g3JlW2PQM7MA4YdQmkXFxaR+IGjI7VwZ3AHhcoNgKa8BNoqB7Hco+CY
EBYe86+HQOfUd7PO9/9Ve1S+1RH3uu8YPwtapRuhT6S3iXRlzDfr2k6ycO/20vaOOkRwhRJel10b
v/HsDqadxwVC2I85lLcTeYZPXkRGkHUUC+D21/1coQDwONvYVi3bHCx8cGrqfCizoFH1+oxiV1MJ
uoWDalD5PCosmtza90CJYDlMWRzEyINGkWilzVk/Eg2QxDD3s88RM+KoCw4+JNFsdxu0RBAu67aP
GL45N/B9qvm/lBC4K/JdzveginnNyu73aMAb64JSB3lwGzGyOUjTc381Lpa8Hil/MbDbzeX/iysh
XHq0THX4qvtLZUoS0fCXF8/Y+3KuJFX7hZu510+2598twPRxz7I4aLoLVfGRGy4LVefrZe5vZ9YJ
6t7mTaaatQjBsMDfu5KamcA4vYNRlgNAyZ8ldW6F9BUl4sN+q9k0460mNYcQGcYxrBmkVLO+A9ez
GaCoMLeYn1iisLD6w9FA1O2ZVsaSGdIqWtYOpgIUdRi7pZ0R5qb6/kaHgiIGEfPw1FoGuIOS502J
UYGMJdUkrdmPnzReT2OmcnQbCJPRyOeZj6MUuROa3QAZKQegaGq/znXwAhbQmtnPU35OsMQtx01m
SUANf+763XoucxFnnm38EkV2KOUcRNipvP8cE+QMDC9bjzaQLdtOwI4/SqVaWt0V2a72MSwws7k9
Bd4A4ZVgVvhwDAJrFsHBtF5SHnwevUE99uHbS0ZAYV32K09wmFeVsi7OFcE61vEfY7D1vK7gH7N+
yYFYWm4+svpbHC8KHcjqqZtVBUKrcHhWiSFv1byi8btKlxDZ7YRloypUss+3JQ4IJl1DU0JViIH6
8kWCTGHChWgi6joT4vq/OTI+C3kAL85MCUGw6tQoGjMgkDFpmL0JSxVIqJ8FGiOMTMTJFMDM/H7s
/xhMaav/s8IqhU5dwBDZHEFuuffbimHC9xFZTYCpOgTrBpicvpe6/+1OmlWK/lbmz6L/7aKo+yZ9
6qyUcZNGrEpkIESa02NCTihm7dzHhrWS+xQnBPejf64Uag2p6gCMbhVWcy7c759oOkjgMp4iGxHQ
mJK/IhTZxfRvKQJCa3uel44ANIE1yCLyoqefWBvBRsA/W3z2/7LtCPW8vQw3T8vq87yBEFstGE2t
mCZcvWITJF5X71NLZqanEh9awAZHwSZbWatrLwVWv0zYoPlFV9JLRfrLJ385FgFM+Up+MsBHFhIx
n2SaKfAgWtelajHhGghyCCZEUwejqMivOKQR0fInVC26QFjD0YbAzxZja9WvX1M/yiVtQVa5BCG5
cEeTKYN0ja06OP7Mgo+49aP7Euyr5juLoEWSwlyumYRRyLTbvneRlb8erjR1t2YVGtQNc8SGVabG
iD7XvLVJ6MLxQR6qYNEPBx75GuEVqU/ugi+eHWiDZBedXAR5FdRrQWxvNp7npJjRauS1QuLydBLy
5u3PeRR2MS0ZEpPnDwbryjYhihZGfiyrB43WyXi+OwCYstxWOhpWEYGxQFIAblokngccgXI7m8gX
KlHhlbGSi/8EEr8T7JneVa3mT7Wam5Q8cWK3d9x1jKO6BA4cv3md9uo6+qZE0lxGJ0NPBDcfoB2r
Iz6XpFi6/3X12ayvpQA+iEb/t9vrZAxFMN8wWun6ivsVLCtbI1eqQJ7Xt/nzy6QACgcrOZQqUj59
UgfwMva1lcpM3bsT5sB1RH3qi/K05931rkbjpgjJ46h0kA4LIQfH8C61pFnNkrwqpf4JVjdDHQ+a
o40sNDtizI3y7yMFxhsRRLzx9j3J2RT1zTkSAxGaSBSHOkXgxZgYk7xL8jqGUtbtwvFWY7evYRte
aLr88Dqt56G4euX/nGlIv/UESVzk9nPLj8TYMVDzrmw8Y1zzjflzGdoWUXFTJVBxPo/Erco0QIgs
qKMYu9V3dxkP/4ypPlQdyxt1hDC/trNWySheELkRg8AKtIIZ6LyIkMmzbQvyFiGnV4v6OZ4qnGiE
CC+DtlhlQTGh5eZT3b7D7sKBD5DlYks/nv9A67gul4hLvYJkx7x4qudY1I8rlSZkLPo+ssRpA81n
iFQBYCgw6nyhlZo4LQCpXLKHlOVU1ANN5bLBotdbHAj30lbsJJb9mFZ/ihZHpTjc3qgNQgN8XbfB
0sKg1Merd+kfiXyJl2Ew8kJNcl3mcXmI72YtXW81RFIaZej28YW2NKayNji1Apks08VNIylts+v4
9n5GbyI/DCjYA9QCsjbFTQj/+mGFmuOiFkSWU4dsiX0oy5rxbnFpDI05MZb/4hRjfDIDOV/qYeJt
A/VCxQ0E72ExuqxFmqxtHrNYtRQjdf7sigBdmgAWx5CohZ0CMG9ncQalyUNsdV1IhjE7/fjrL9sD
FMkzA0JspSGQA27cekbB4MLgPO3lesg+kv8AgnnvPfMThPHaiXfSw1uo2F4fZy2y1lPYPvxEuA0b
JJtmeCLCIE+VcFGEfOENDhtL/vJMyCKbhRoH08XtdfwvaL9jrB+3XYmAk5YL8RmY6Ujg1drbX67O
ZLdYihdAT7QPY1KuYeKjOQi5RFAPJDeGExeUC4uP9C/kLhYCe7Az71V7ALacHd4FidJ6QpcTvpNy
/cz3GY75HI2CrgLpw+9KCtMG53ZaFl0kp09A8UGaz/ArWjtuF2D4puEzloG6H6/2Mj4cJ2q+O8+c
w9Pdo6iCPQfxYZez5FPpFpUi4z4zRH/jHHLagtIpz9BJ3qLuTsAz8i/2VceBFqGV0iSJHlCztjsJ
IBL8ZZHraSgndjQ+eB4Qtp4vRPU8SoyrOYif2Qz9RkrVG/SdTtedvZIqfJmZmTKhNs5DGvLt3JSW
9ybUPzLtQhiApwBklIAIx7Jb+kqlBTMwiJ/vYbvrGg28zGLHL1hGHNAKkIwinluzNgtf5AV/OeCy
XKpTcaaPP0EShTQ1PVx1bfCskTwOhhDZT8kd4sq29V8nHY/1URnuPiS4l/y+cjZKAcWokOc9OaNz
UdfBr8ji36/wPumdem4e6dn/uCxNjcP3vsEPZe9cmz4RGa5ek6yHaJaMn1I8BGT90aVe1PqmS1k9
DRh/6SUysGm8TduTbyFtjyFLNcpjLYG9CEjUoidK9y9Z13Mick4IYIstu0FHFMA8VgvnYyXmpHMX
coXr/5uvslHOUfEWkupF6wnC+MXmQsqtqk8Rf3KIpAXDEMlwPepsehYKHQ124sxR1vDSxUvnnHNS
lFli2igpLLp6Eelpeea9cA3rWhoZePi35VOrhPBqjZfxbfKEPYt2toZt+zRnVhkjjXIKcahDmXwu
n8ZvifH6VOZM1J1ozRs+MGPhsPWtzPZzetr0FKH14NcHSQNqZGdPvTMXgqO4JCLnvqYmazjXdIy2
TswaPBHKiM8EsUOra1KeXNbzkhMvxmKeH/0qB0fyKR6FWss2W4fsXZ7zRLudpFmXvZQXMjue93pK
DCvv2w9MuGTk7kjMBA/IhCXq+SWG7Lx/p1iSY/oLdP34Z7I/q46KCWweJEwSFtl5WteVTNfDLGa6
4i3j9dXlhmC+4lmv6wbqB+FxOLo7ODXd1FMDzQoHb5JiM9kx+zhFO1QtVVfMBbiUHtO3H2z44wT5
fqNAeV7XOHYwyv2u4A0a6lqZ+Q1+hTjTh95Vd7QHuoNqwMoCscZqfv2hWXbycpybIHbPcxAu8Fld
c09crA93ce9oSYVTCTjmek/21umog7b8jb79ffQSBunkkfPr5+3JzpMDPkb3XVb5SLvNlMLyU2bH
1pnujAJoi2w854v2JzZ4OlzcebFzOFBk2x0j04PZ2FH4I94xD/K3fGMcdqeIMDUZVxXkj7atBnl6
XPKpDlMiLUvXepYCH6sUDohZAAWxBkMXsC+ZlliLlQ6C1m7oO4U87Tw8tCJ73tIw4/eltDatXHqh
o/aLuT5hpQKDi22QtABKx5Ak6KsRoO6ZVobQB1rvJ7tMWdW96octYsgMS2R68w6cqhLjfcb3jY5A
CxS9MqtaaMyLctTe1j6SBNbVv+ZMfZVTDwzd0r6VnoNHdOGOEzfSubNtdmJD04dBC0OkQAfkRuAz
AOGxaTa/kEIK+fwdqiWeP2VUncdNlzcmZ6Gr27FPcZo9bD9ibpHO1tbj9oP9hI/7z8rNJC/u/hS1
TZD222P4BgL0WdjgQC2pZZ0vhVroBda8OQ8KrTzyi+7M4EXNnbdEhgKtprCRM/X1CCZNmGq4/E0U
OxI5vSfnKPLmtJBTeyEmZtZRFC/fC5LZQK3fiZ0FLyp84O7yllvx7Yd3PzUy97KBLGDgp8tooTap
bHI6edfnm9lKFeZatig4po4A4NiAl8/qoYXnJbIpOzgW5YFn5NAj+sEBDFlzMoknRyQLzU8QK/jK
u2sI2ygl+PcREjXa5dp+42PxY0ctmXQiQyLKvk6Vk4roAV89m78aQW1drTcs9HBndYsCy5fewd6/
9v9DXQNSToZG7OFNY6c7+RT2oQ0Xfy9wZiXePe/YctbZiaOFacPdm6uGeAMdpFbrU8E8xAXpYPGy
Jtau2k9xdvZTAFDB3ujT+QH3Pal3U9cc7HdajOVrF4MKN3RcZMDrwdnqn8pCwtA9A3XyapqwF9dZ
U0bA4SV+WVTFw452JLaSEKBlkAONWmNR315FFN9z1B4jhBhPK6xodukZqSN3eDLHqm+UkVtONBtf
QW1yzHhQSTT5cutlUsxrWgqMuu4bKZtn9529UkSo2JczoJsbxDlZahHHFdgslbzzXTMlqelWEGxE
HNV/Dv/TzWzIheieOrwtpsyQ3tJbDiwoYKhGwOYvboUtRFrKO3ilIbd2OoZNTX2+yF9yZ38FONx7
zeMfG/pM0k7OdmkJbHNax98xmVVDzRClUJcIpqj2LBErCpFloKxp8gcEpHoJwWlZJ7QTfNsW/vmc
o+IHh7O7h4apeooaBNvyzl98arOZoCLO5cAGkc1KJjsntcnat5ea8P1GvjXuRBSC8jVG14bZ5YgR
iOSb+eU2xgTlWHQ4dF1ui8vmfN6VCe5Xvy7aziZUZ6iWKtmLwVuQrXRlkoVfXmK0o+8yWxiyN95I
TnJ4kF3nTvZ0u5pflidr+57MOo7lqCgkzNOj7YS65saI6yAtIzAmj+KnRkgpShZWXDGZpFMcre0z
yLGeuq7C4t5KReeKXeODhY1iY2hDpJYj75Ic5aNFtqGwhCi67olxDkBjCVAJmFRRUUliGoi2UWAn
axdY5EPm0lOhYNqLyUKGYTmhd9TKxfKq2OOKoZDvFF8NlB7eOhL5+Ef/hCwLU8IdAuOIDXNNWHX4
kf7zGAEVzUH0aECcE7kW3pZanaggRXPZ9q3ogPQX7LRLF9d8pR93KrqE48Q21cF2Yd+agMmJNpyA
1+E2rFCDelxhNQjsJbIcQHGEoGco3hHLu2gJYFPYlh8Qk5rSCqYl2bpYY1v9x9R5yXF5ccBjsYL1
AdKyzclkKTLcaIqQ9rhFR5bB0qQgFIzitwGQ0qWJCxUiHaBLdsjl+pq51ZeQTJZt0J+vu9TPTF9N
EKIxUEIdhKJ84Sk79p8y3kgoI3eZi8JWIITR2g8pmG3ckb1BHivmncP/CEvIvHHlz24llG4laPCP
ON/FSzECjezPF8TW6s6rkWEtPeEsgbp3bZOuXq5aC9XJ1Of5i1hXHF/12LgYlYRc7QWL9ELz7naS
5wPexf39hF0qAE8bMt6cvsZnmppEf8/ZYDHNtWJdGYNNgiIDghe4mRd+BEex4i2l68Q3X/XMhzt3
p4DM6a65oh81w64cRIOeJ+cv87ebt3w5kkNQdp+he/I5OLl4k5qcU0uJNTDmoMrynxge8GMPN5h3
UI/pj650xV4rkflND9D4fFhjdp5EUWt4s5IiblVWhPp+CSEi33L3E4BElA+kV9ozPEwvq/gHcNFF
vnfgcqeMos639Dxgo10pmbXjBMW/df6hx/NsdlQRyA4SOwMpHUGYQxbp5pMCHPHI8GHW203L2WHG
W2KlWld2TQ3+5I4vrp7juZ7pxtdPlxEroORptlAIDe06g8QQ/PazSyXGApbUVfMWQCJkkzKGizmw
OiherD/BGEdn0OmYmwcDz76XqO6B7kFgjhl9NgtPiLzwsEnYKKlU4pF/gO4sSSvUrb20ZvKgc8SP
lwd1TIz7+owjqqARY/p10mZiRsVqwvE9I4dc3BJlnftnev6n4LM2RmNvAai7vRuJQTBzx6pNF80+
vpilf8N3ecigSj3gBvNwP3OpqTLCN063XNAUG6eW0Yp7DKfqoIC+tmS6xO2nTlf5WoDvwgze1nyV
eEHkHj1G5YhGrFuSveUhmPoY6z3pGu5gDupDDfko4oxitLsSbbqFbGH2RkVj6MW9oBmiFAjLcb+F
ac5dIzuW3Pci4gqiPckLtsphtfdl7N2rGAlESZgc3auu8qleXyjnFgdrQTp9WoLewb/6fFO1XK8x
UWt9STWRK0Y0HtmaJmv4//Jh/NTZog7WA3/zBIp3D87QauVV+H0gZyz+bowRG2t+URKrVUNlA2CG
66D7Ks0poEmCDznZhw6NMcJCvtlnmfcoXhtIj6X+lh5+p3UxVza+P1DVKi5oJEJUE+aSPkKeNMN4
DGVhxr1hGkHMfnBEwteMxHyhbtGtbm+DfZU+Vg6UFglr40i0W6EgXkREvoS9GsfyUe/YoBzD7DBl
P59BOL8RJ2c3xIz6gVPlW/JVNDyxg2SdlMqA+rCaBJtsD/ruUaiSdwnPvw6+YK6wmG7H06dRahIe
LlY82aPJgGae6jPOfmF5LkPZsI2iqvkLiNw9pbSG9QibJkainCb9jAQqPcCW07kjpeN9AMD8gvdL
5qUdl3YMiKuYmfome4VfHP4oNd91Z26e8w4Vj1v2ekl8R8ejbj6ICPHysMmnvFx28DFa86yGTIMk
4ei8GgwuPrKWRE7o83BEHZtDU14pu/w+0j5UKUpBbht7e2AwCq+SHPg4lKitUz3Bvy95B+Tzs0PS
cX0n4oc4ZN+OsnsnZBs9put13nEuKGLgjFNsLzRBB0YjglZ/FJihDlhtlOL8tr+0PAlE6b9RPoz1
YXDcf7R5epzupl22GaQeLo7bBVdEWH8jniTLc3pnn74WXIHkL9XttTBVWTlU6RMV06yeQMtyg2+o
baLmvmpzRfQGJEgmONkfmCew2HMm/aKEG23uxT5tnQ0/8MGRULCUAuZA9WELzW8pWhqdfs8VR5Tf
kmAqtZeCNFK3t75tAda4e6/R1jeMJ0q73jIfGaKbDAG/1EMQeSQ6wvldMpu3vYO94IrWjJirb2bh
k2qsAyeG5eeKOhtdZ25FbkPQw9HeMDxiGO1t8ZR34r4NIgfP0JedxUX4F9WuI3UfG9a62VXsNtsv
LvblKv5SRdQ57gOgdsMKTtZI0Z8x/gzhK6kEfJmGTatsNdWFCkiwsTOkcSh+z/XO8VmSZLxs4c/t
FxFL1qz+5dbWKpALIwN5p7LiYHyPw8xddepf1qw50Uj8CQNziLkGyL79oKo17JVx2eiSscQ+q341
eZf6Qflu7L4Kn873jSatZm9aO2SFRUb6mHKGF+FlOeeDlRIpyTQz/bcS3pQWQGDY4GeilvlKQZbC
uK3DUk0mgbBrmDKCufF7liGOssBf167g1ptopwpQ6scmmqJFRxspdrcqNj64o2rN61S7JT0t++XW
WtiFNYAuE6QdW1Op7Zuu9PCDwyO/+BC0gd3E10NRYv7xeAq6Yk+YvfRfEJAa5+P5aFSBiePcpxIH
2TmrRA9D61vKk4/giNcKUaZPLbuhXWcMRO8Y6pLQqLNrvARXOO0U2FYYYGkUqD9I7wbVM4OydbHW
fNdrLeh3pVLAVlCmksGS+8WB9lpb6W9pCd355W5nJIg4YBWZKsCXMUPUGcbB5Z92zNWqKPq0z9Ha
r4jIuDZlS6xKAt4JSvlloAJScO42HvH39D6wZCQrPnYlbPcW6TCwSLtXE/KRrmlp71hbL1e3ECzd
178j2NqsMDLO6nJjMGbjdJUbMMq4GPeIojcjiPUoqS4RyN3LGi9nrFqrS7KvRFpkTcxoUL726Z4I
FmQou4AkxQyTVQbShcwD8gRdIBTbtbP/q3WotCK4dj9GhieqcKrr1txPGYYAPpHFXquNIv8Y4ceu
6iIpOUyS6bJZzNKQjW/OWxSBCa7aEC2IA3Ze99S5y2X/lZiJSU1+524foT3cw4Wer3XEMqs7HofP
rk//XWKqZQE6AyyrFihrsqgvN76pN7UAM41ImM5w4TdLdtJ9ag0hDjCh7IPYMrdaBWOSwP00vbpN
A223iOSa0jWSQZh6OXDqOiE9ukY4acj8D5VJvJTooyrlLuuEhp/R2ezU4+05LjzcbuiKhUcVuN/d
kNJQYxuNpo22UHnNhg3TDAA3N4mbpsE0/KGhFleCOizvmd/ZLjqy7NuejAJYV29yGlpqiSPknXvn
8fDOkSNU03OewtcPdvYReMI3v9jla9iRSw6E5l2kxI8HcbZ0xAY3YtFpd58vSFC7pbDmjaGSxIdf
aaSU3qJFrpTKTy3gjLiULrr6aD1AqpxhontygC62c26nFIc8PsO2c5FkxPB6QNWvsSzTze4rQBoo
CF3K17P7QlPoUEtaa4QTVlmYputOwvDd/ftUygP+QBNaFF3uJt/6OJ0KsLfbq9ZBCc6DGuSQ4AMc
wlfb6cj4IpGKQAqVEY+NOXOAF1kVCZueGRHIL8TkmHOa8IwEJEMnO5mRCXpYY6kRHZvwEye6k7Y4
Hyao0oBIk7tmfjj+4vUB2ebDRRG9HcZY4ARzHxiA1WfhU5D+xLonlQCH5dvDTS+XVxI2TQPcav3N
jWK/4rw14D9GbZ5+f8Ij1u2/VzG+EqdHlOeMaeU6FU9/jjef8AyBmfQgqHYn3/yaqXOuR5yPEAHx
iwkQSKcXeeQMN021qjrBGBo1lpBzVQH1B6AZ5UNiHBRDuwrG+IMaDTz8Zyed4mNAyU/UWOA6nYVk
opzFjf1KHCX5wJOiOEEMg0tdLhVcMMxaBLwSGA5jg4DrlZSONLuRx5Mfu6zW5pGdHmDwy7fypjm/
+wWxHFtoQrojgI/pw2tbrscwSj1qqKwDaeLQPlmdQbgVllYSqnguWm05MgH2TwkNDKa+mWj5gUGy
8k+Gid+ZA1kCRprSp6x85HDlf/AqWwssc8G5ICWW3jdVHQ5XqACpj6+JBv+knBOqLYiqWkL0CdxH
rz4J7do2f3qkroqI9GY268c55kiSXEdVuR+06tkrm/lR8Crl5Ync6QUI2W0AWkwav9V8Va3NY7Xb
S6HTdyACfrw2rhy4FtDyIMWJnypEH22ZnERkmOtvzDxvHfeeeXdGvDDydTGfr3WwdGPD8iVQzTRU
TfSJ66qmezk9d6A2fnVQ5jSR9mMUh2bqHb/facZFgRNf5JSWM6SWIv3UyOew8mvW4Jb7PZ2uv+zQ
iDsifolYWo8VAkKsdJqr53N1jTVh4Kqdg/tZTsOoO0ZqDi578s2vN/c8UOs9zfrsqHfzil98S++Y
Pmkp5GdsT7LzArV6T8c08XlwFl2dKtHqSfXWfkJ4dQkjqhI99my/Zb6NMB9ZmI7PlfFaTpY6TiM7
fro6Dus++bs5jZHbNqKLEeitMENeFY6UOQrE5aqRZWSIYT5J6ObiVqiSN4iBfY6gRjpVkvDYD+SS
VGRVixir98FT8iZt5/e3iF3hmWHBZw0es5KH5AVB9PJrodb/AUifqs5KObtGFD8PwVat/rJKS3ms
AVa84F9iFaWtwFwEDY/u1SGMWt87ysSe2CB0QWNGYjadOs37rNNobtcWtuki4Th9yfOaqJljUFY3
X0vZOGaxQUhfTPyGHO/fMBnCzCZ7CUjaZB6H5fzr0jBwsvWtbnUgO2keAN7zTgsDZqpnnzWCtLIT
5nwbfVhE4HjZmFltN8AxmQCBGyr3vQGATndn6Lc3qAw6gDODyVWZuZG4jjQ6LQTpXcJ1cmqscg7/
i+2tnymzyMjaeNE+mvf5xmVTos+jBYEUSxw1SCCTGrKtPrkdDeA+tk1A7GUFGVyRgpqBTSjBQJjI
JwRVCMtttaN887tZ5YslGO0bIr+GMUjD5zV1q/7GyC0IVH+JTSe7PFNR8/87mXZVgGOiy+KBs+O8
T1LYYKolqOyHb19eaiI5AZHW7jN1YYIJ+m7G1tJGpizQYVOczEGarFfmriOGXJ30KCfinGiLSqA5
TZrTphhfCQqaQ/TsVq8GdyvP+pZUD1O5o60+a8fHA6kX//n2bMYwl60Fbki5ja3ZznFA5rzpgHwH
v0jhnbuW0Z9vucR0SCD+CpRr9KP2YMchcXlGjhGSGd6dgXuIHf2+0Gz/1/AQYeNZBubZIkBpvUDy
GGyl/O67kRB6JE1XMVwZuyBqJXI3spKPbpB1YJkZcI3MQ4p7E/p4tgtccL4jRLPAGj8fY+4lyIsm
a8hfBua0l2ToUyGGsAAEy5tAx/Xb9lql+dZygqaijEvTF8J+leAlfgBBBrIhcncPGnituvlPoZzJ
3xGrj9nLnxYnjajUp7TyW3h/hI5dyDlu9QwzG+xkfFxvFsBQRTwttbzfb9sFzDZ9w7JMV5sBJ6s3
k9zHpGWUn95iZL3LHZAdVL3mT1wL5ruLSVHiAyWMJjiqhjNIST+R3oYX1t1i+cE7Z8+J62sAj+Oa
HGXRdouFMa/4pjYOVPlv92dOfjKx8QfKVtyuVbHPABCLXbzqTIWs2MgZ2uF8UYBUUDe+HC7zmkEK
vHquqape/KicpfGPumO/ppcyMjbpDUHKIaPD5UIslbLrrDw/pxKGOlh1gzVpXy8tw72vtks986yD
qkLKI9W1pDAzHcA3mXtoLOnBdSL7OQ1RfzhtJrIWXfVJjSeormLGpu+9KUcMJkbaQgfZ2SDazABr
MX018AKaN7SrnncafjtW/YtviuSkR5cPzAPLoWMlIG+Nrh1Yl/r+jeX2fpvbF1EO0dMPo5PUtnQ/
WcAm2uLTnB3tB8znGC/35W5yPpG5GaWhh/XAimxI12Co4AY9LK2tRMoIbsVS7jIOzHbsRUNADHla
Z6HnTvsPUrCp3Stzb9he/YGmype29VjDewHa0XA0xgxYlX6bqMh1hDU3iuA8DTZr9TwxWn78s6ad
WLwBd/GG3RNJKkdlgCJcEdmKlFUmLzKLR8hNmt/AhjqEOPBnBe6tGM2tYKn+WowbmyjQasIBU7dS
qIF03nPzX3hSgny7y1zDBSP9GR+M2oaUm2Rx1soSvyQyhRQIe9WkMUZihWpLXqa3XtkNYrABr7aO
lv7tbmqWbgukhzlOqwnYWUXAkgdGiOf2bBIn4Gh5401rcgH4I7z/hQk9tlijHPrr9EY7dCZHlHxH
JZWQLsMc3c1sHLnRZCiTPY4EsrH2UXNbavov4hNpSOfP5UGWZJqnsJqmr7a09VPraCPB4U4OD190
RVWLBi7BsHqaDchscRAim1mLX06s+xVfeTXTJvSOkbdN7YGSpNDc1sOILFay159CT43VFBrbOkCV
z/Dw+66DdY6KA2RocJ3N/qOCZOFCmT/aqUTPOpzeYFMYOSbPzxFs84VvE10/JIX8qkg67/PfG8nA
z9VpLNLaKe673excxdTS+YFOo7hZSgQI7fdd7lYm2UOpQ6rWwy2GPldjNRSuCZd58aG0r4VSlNrH
WLzWRSCjNiMLyLQNt7QCXO/EUF66MN1+8/P06u8t525GaQUDORFvQ8eI3u4VlmVWTydbkFPj0dsc
37zMOzGV8EVtjoZNEYUpLYGaPglgh7W11dpNf4sqXsloljpdVVSa24p637Q/LyG31fq4WaUVl9ES
rsi7TmKsWxxX7OSDb3qb78dNUb7RC7wPRhlziEnlVBvjI6PNI0amPCyYNA9caRWF+64/GQ2dIJhu
P7Zue8Am0UebH+VtnBCKYkF+l/94LUmwXY+jvKarX3urQm6uzLlOmkZiTQquMni4QAH+oItzatWt
NJHv7LEVuwP2JtY45/EYZNR8uvVcS3ZSGl4oC3EEVa0LX/VqLrHqLam8eH12lVog9o8qVduyyZST
3ED4Y55FQ8MEGSwtwFR5OZSoVDcnBvw6qoNB/A337HJ21yUPluIlYJn6zqMgIMxPQjQru2mTOy1N
gK+6berfcKwRveBaRCvKPZyN9PODvOw5hHR8f9KlmWHD5/83vlq+C7dBPXRJ3igYtkNsW2z2wkyh
gICnZ8APJesqZQeFtlFll1M4QH6RSI3Td6Oy6+9rZCDP24dzHbKrHo78jdFnY+X/kkoezjS1TQYi
EaSs9V/lITkk/eDW7o1FMEO8sEXIN+W8pwf2ntwQnDwcddfHavaxdLRA0nBJ/rFufWnkcTpmpNXU
/i3hhDfqtl2jLcwZY7uDlocEweWq6hFyumIKA3rujJW0gTVdnME/ntKj792tPZwOCTHkB5npR+Nd
MaWvS45RmEtQU4Qjd5BzFLVHXgv0VYuQe+//NmWdN7mlU3Bcmh6x8Z3KbY4+9oTpFduHidYXJuXG
iK3qp5N2YhpFiAEx4iBuuMPrSIT3c5NNMUiHBYg9DlxCRux6sWiPX+lLKHn/4W9GtLSM8EZaRBNc
8J2vySJSrbXy/tHZXeHPBmmlIFErj9nrHl6SmNPARVH/+Sb56XYH/wiiZ+yXhPHt0hjsb35HWeKg
S0/BcJCFcwZtruxqzn+wZ+sE4GHasZEjklp6DfISvKUC4NUYD56KZ8MEpM0BxCLiWcJbwJUu+pmN
ru4f/Oo0WyKr/9y+OzIUEucb8T2h1Vkmrm+bSqdMx07Orle3lkqpS7WOCbmqiAvApq0mC2ZVW4Cj
FkD6xe760ennMXpjyZYvsyC6eGsKxHxIv+r7C5Ojto65mhZel6nYeomJmuklOWjMLW+VfTOwpmI1
qDNky/r1foU8MKQ5pMShPc+/tD/dYExsBRQ5cKA4mNVxSh2L+2iGUUFQ1gfQRAF9P0vDfZACXYo/
OlZPTXW4xwbnv5zTQLki95SMsPRayoawc5Yr8mAkN68ZwQWCAaIcpzAzT3UBu0+f8d61lfRVb8yJ
XmcHpnAH/d9Uobvpo4JkK35zRM72EY6L1g/w8Vvp92iqqOvfKj9UtCgPM+1fzEtVS4oxBlX0HMcI
b2N6ZsVODHCH1NLdd1iEpLMoY91e5Ybg4jc/exZdgniDjnL99+s14byICfNzZ0l+UASKiSN3WPis
J8HVWjs1mdLNAQgT63guBR0DOIGzFBRHfPQdyE8ZbTk88og95wKqBWeicebMnHktMy8Ic3vmfo2B
p43hOyBG0E5aMZlWB7E9M5SyWrRc0sq20BQ9PPb76Xa+D1PSl1Yg+7QORlp/tsvWrcfjdzkcrSGR
T9OfuRx5VO7WmMyepzWOwbEK1bvwRd9OhZwr8FmHGHbQuSM7X7hrp43SEs/laXa5ENFHbvQjW7iu
HTCCrYnt9C9Z3Me0qF4I09mSF8j7ciqEyTpSoGbMFgNzCC63f7IPT7b7gDMB5vRzHW2+3222K49U
hQNpVU2ZVroGQmK3UTfMSlPDKaJ5Otl3svDu1yCaGG3BIChWlSahanI2fmQj2Uhy1LBUx0eaIcHi
a3fKp7hsupuG9DXR1cxnbO8UMCxM/RRsizCKZQ75B3kXGR4TBLFZIwvG2LnYWHyslgHJRteepgcW
TlaggA5GDFSotK/ncwbLT6+wYKRpvR6APRjVcb9Mx7ksU38bI4qX+to9pm8Fs99gJEqanF4tguyJ
ycWdFHFM+V9A0F2Mt9Q7tXofGcDm9t0Xir9SqADS1IcjUgryanXIJjx5JXjjGT/wBKWI/n5dz9o0
B4CxK+8QQ4T7K6gixditbdfwlTyJw4is4UdVGDju40ZGjZHsGD2cUWDmKhTshwoS220caSk1fzIj
rFkIg3mSik5daMF7eILwKHLVpFZp0XgaX4ct2KzQEAA2HLMIUNFiYKaN57pkSVISa5Oqj8AIln07
3cnk0lGdjfz/eKel7RLyUAi/5X0YqqHS9TtgkQwdmY+hw0QdVMpVWmQJJhvz/m0XG9nRsTa3Q20R
prEq0nogvHodKNHsuXMSgMdOWyIScIqFZDK+WPYtpKl+bPBuIifEA7pkqH7jUCeKdREQLog7sjUE
yPZUm9sWBQBa6NNtdImIyZEG8uL/GAF3FfNL5G4Jy3dHQbBLuXO7k88mBUTQNcAwg3zx/szeVDyc
oVGYnIiXeuxdesvivcvaC6gVh3hKxULCeRh3Yj+H5czZZwsZFFXewLLbv+FrMPYHILpzSmW5oLJJ
mGBy9PgD+r+e98Mjaj3JSbIwPhJd7MEOT0HOXS99b3JjB2CD5TQhpnDo1uJx/sIYMJOxCI4lNt1N
yWy96kRO3/3QM0PabEwCeNkn/uB9I4f8PHijcQ3K0TD+2shHkqUDwXYCNYFYMjy6aYDMj8QTg6X0
popf2+6Hxnn8HJOnsyvSS4MJUgxUiIsa3CTd2TbJ/Enk3hkdzC2J1HjfkBuxfnYull/JIXawo95i
sWHUzCNlpFQpfWkbkr/E3waqvZ94rpFt7DYlZfxg5aLUFI1hkR3/w/pzmaGMwwToPAbbjyo90b6V
+6zslngu5RZWm121rOuMXiFrEUAsVcmDYYu4H+VVhO1J/HFTY3pdFSz5J44EoQRDssEsTxcYYGgg
FgfbrWPD6n0JaXEWuIUlzP3nWtb1HkefbESdzq4ivakXE/+TSrQhZzT8V2YdhUMZgbKE2qXABwZf
iIzNeKKU117iSSSnLjyKSq5NIXtHkkxtfU3JjtHcWKeNryQ3dQgi0/DJIktI3RvjMAoePYw0uKgX
w6PeVRxLRRTttGRsFDpzZsOwEnQ5Oy0xAqH8uXuQgT7itLdh80fs+DL3u16qUFs8qmxZVHRM4XaK
89uo9xtsunI8IrsAMWa6BCL4yIXF0HsFRmTtCWAkQd0PlVB5Ruzob0jscE94Hw6TnkrI1zi96IvR
szAPMDYf2pnhweVzBQE8RIibJoh2JP8MG/gHX3n07SPJJrexywUT7z9eDZZmX+McXhF46v1+m4qW
TKC/3PAFBG2xfVfwG4gXfY2BqqSw6/8k8JSEFsAC0aI5Bt32NqextTXdWhfSRLC6KPriUiPZj8IC
iQWykuEPyeUsphSXPy17jzf3omRddXzz7s/P/BAgfbgNkYNNCwDwFS4fKh8SKubXraYQ13IxjmR8
DnjqatMZcJEXxTFeH/idCYXRgLLxmVoZAAtiXCTuetjLCYR9y7f0pwq5evBLDHNITKhWBD8ziXPF
u6fDtkdkwQW+arnZSlUytPrFpjKkyVgVE6xnAdL7YUJVZGgg9sFvuuXM1+F8J09+7MxESSNpjvFC
u/+xFd9/03/8CdcrJwbUiz8PysMqMlkyQQz9uGj6qItYGQETnlO4vM/D4V5daS2EUppABpV9ZIJ2
O0cufzVimbgaruSswnItU1l7VIsXlWzvJ80VCyZ6PUGg6hcC838hsQ7wNKyXSCYVHleVruzHGoIm
X6T0oplyhJ0RLBbad10u5FgMsEqs5S8RIKnf1BUafl55ywSmPiHyazqInIu9kGjVPz0GOr9bpn5Q
SS/1wQGCxcYfJhZQcdZKWAOkt+BhulJVbkBzSv7QFiLpaJ3RhgkBXqDWMWtUeOqjq6PAKmhEgVJx
4SM4svonUrzjuRJV4AUWW9Q9A59HskLHfNUPGjXdKCDpEuhtPJwPs+fxYSmwDLeU+vdSv081ONpC
A9EkpmkH9O7Aktn3WVXCQFKOwnozwiS55KepQteo6S6YhgliRQAkmIDVwJvfO+3a4MOmrg2vKk0I
IzLIwffmDXtzEVvocxDanbLN6W6gn3Qz8On1Y4DWOOlrzvdsSk9tQ1F08hgXGE4PppSNDDk4m0Hp
Ya2xOYymMILt/3TUjbt2/fOVUNxXVyw1L7HV/dzj7RhP3EteOjN7FYxNzrisvPL42LloaxTFh3qE
hzIMObOCMwvrD/PQ7wZOgHhC7giLkYc58fv4UxBFCOTjH/3/6qU6Dagfas0w8XvQRj4cihoPEX4O
9ZVnwB9Kla10xCB7mT20Igt/WQwKzAP1HBhsNC6XBy565h8xuNNSwAyWNrCg5FZqb2Uzl6MOF6X3
JrUKsYVM6H83pN5+1RHIHJFRZ3ppo+MKmIMzbxPpIDKByCyQga2dmE5YES3eX2kpi5mmW/KNvNUn
h0HESfZqTOAT4+gYAzH81GM/ayOn4NyahjcvRtatlniYTZAr3UFeAMxQkOsgVlVfSYO6YAxfXCvA
WM+IMdVEBDLLr64zt0kd532xK7LK0CeN2asVxiwpP/QziYmnYaAEDDMg9RHXCAB0xjaxJh6kWpu6
Cgj50m0+EDdVEQsqh992Z/DHyHdujjlC/oyJU2CdKcF/64d2DzJzRq8ez0GU59iDuyhgXU7MmBsy
pqw06OiqTv4rxwdCarmgfTNn7XPeNprQq3zOCuK5d9Q/IZkLAnBGUEpnBaVCpX+/5wXPYA4CodiA
RZWu7Lfnl6WFh6iLn1shY6nWplKa/vZRQ3H3oclWaxgElczVeWNotixD1o0jy7fvoXZk63PzrjCv
rAdgR9ZHBErKaDmR6UQ/6VcVitAsV9IVJEr4+CsJ68ZGN7pmLRULdts+9/ReE/7ux07FPaHHWAIL
jpyXWhxfT1LkbOOm1j8U+glt0Ja2Q+WPPS74Vto5wgHfMTCe/fKygM2nt5LbV86DsqXNjD8X7X1K
rdIHbe9x4+mAugMtLyGAaVq5GBYxZXzatqvMFBen4cYYgfTUq4i1O6++8vTWfMRYBD7xyBm3iB3U
Aval0l1XWG+6t1Ve7EEf7wFPIoseG2vsD54+9wmF0qpWZsCIYDemOqlthJbSgjC+CXpZRA5OrF1J
QhBRCOz8mLYqmvTpX15wXZNnDSsoNYpBVxpF+FMPECdNLUwxQgO2NQZRwgnRHNlhSHrGVKOsF5cp
poDP0kwnos5fF0Mrc2nAWKXZ+dw0uex9FC+yQ5wNKuYqm+y1+MYrjiTyWaa7NSuLZK8R2QfNsNlA
95aupfQ5kU1/wDEJCBWwylzXPdrveciiDVOQ5iWNJKQOoC7+ElvHvquiBRm7h6LOMKiCSTlNiffp
3Hw/r2w2FjDfRpnm73MEkgkMEJKx+FG48E+qvf6feuKLpoHv+kIqJfztocuIO32d1H4Zcc5bkW0h
V5eGyySNyClMhpAXRKtwFIHNqumCOluSnOYEdQEt70nv/dJziR1EpIhfbHVuUFjorislWc7b2MJn
nNumXg4bP9PiIYRZHbWuTHA0k2ryTfgL3T6hbe9vrYu+H0hnr6GmL0YfMzTB2LaYDZFhArqIMNpr
MaViEZtZSorNQe4bFtZ/7eknzvMO+TeQtbPaWJo2tmMdd54+OFgcb6RgCSEH9KBClO1Rhq9MSwm4
EV3Iv7gDzRw/NUKhaXgYE2AzhevvGO7bQRceF1p6Ay56B5aG8GNnWPSYgpouuf2+tR3IxzyI7IVK
NeuDB6cBynsH4QKEkd9TnDOdKVur5XVNw6o8bQGF9+2KqZHWioQOcn5AmJwwyjN/t1hhZwZYtArG
0gKudM/jj0ie6UUeo8dsJIdzQxdy/JWHdLDSPpaVPKWVStCZkb1xsoJ+z0snMhr61XZBmD2uKMhR
jpmRrxs2Djpd2+9tplLfrg7GIr8e473DiT0FyN7HxTL6cWS6TIIS79sGuSGa6pNkXHDcbQp2LVKh
NnVigYahQS2WB8jkazd0WxXee8tgEyemj5iDaEqTBvqmlSc+MJyMSsOk3JteKU59ihzI3cPxUtYJ
1RK1xpUpA1Gcl1qm4/7zLRF2EcvrvDzUncCNXtnW2KTmNucQJIcW3wNWGdoG0RTUkpZZBmRSIpd4
s7zp3vu38p456/4NojQvUVhWYYwZF0qlD1u9Y5I79fjlAgZGMCByS+34TK5sU1VGrh1EkIlABW4E
3U4pLiMuhDQMavpu6lCHqt5GhTw25wTCZ/Yo0jSOdRoxbLxhsyO06nB3d6q7K5KLA8bTu/pXWJGZ
YfR+HTD+6Hla4k0Nz8MZAPsHr4lGU5dBqbZd4l5m/SnADv2zScovlEDBcQAOxH0uBTtYe+g/kTaT
F636ho6s+ydD1GgEnKKOfkUBcUCBztWIAvjZ5+OfwDnFp/4HRkKEdLBbODl7484a3NS9+BzOMG1E
3hPEf4BE1MCESDctKhjLBdWpE55sjDd+x0T7aRnaoQqhgdbNekMweEIhJEYCQm0Wg2xeOfz/7WuE
BD8kg0+n28I7vz3NbzwCGJEObw/zoP52hlcg42Ec51ioAcqT491pAEGDDDbwr1AjhBscThZ3kOvO
VvrRKockzj/ZV9XmJ7gJcuyh8kGC7eN+h275W4LqYMLLnb9Hc8Pm3yJsyF8IhXVQW6M+grRk0tyv
YsNjkyY41t/IA1LbtH80e/f6PkOLf/j1IuuZHrrzHPZSwqJ/Ms4RCo0ZETXusCbK6QaMUywPb6Gb
hvNbX5gQtKEjG90WIJKfYF4xilF/n3eGVRKwrQ/RWXUWKUx+OYuJQ91blHb65J0rqw0+IbQQXARe
3yGGsyXTMoXMcLC3ThtRbCpwelSn5eXRPuPG2CiBsTJwSbTUGbdFHDxjyMSAdBmq97ReLzVEdFh4
BTqzyKJnOJGvWe68pp+BcOJlM8zVsIXse9vPdoyN3qABRuKdcBvun/9AQj2EjiedECkMzn1Ultj5
eTFDJy42M8Dbvnc/sSQySqRen0HKXsi+1axofjzn6wUkh/DcQIzYc1Mb9CnzFITDVPPGaIlTLPNi
h2MyO2XNCaRbXXYlPEL1v2MyAqR62FVQJmweMx8N4gxB39oT+f5gITz9MANQAeAVWTQgSnpuahTw
Q7qeRi6QdfMeFNB2iPg7OH7fvpqDohgLSTAuI9K3Ij0ZPrDTvgpqFwv0XNJ1ZybU6OsExwgot9JI
9JW8RuMBNDNEbveO+IDDoZZ8o7NgLSnctLHcXnHakR7AT1aKsA5nlMi8vvof9HR+ndNTYCcKY1Ta
ZyBaYUcXlewscUSycOkzBtEL/89yUeZQPkwQUnGaqk/DkCdTcmd238xuSUTV3Zk2Lf8zuUlSlHNr
t7BiTKTpgc+P/2FfB1490L038YRz9WhC/kAdCm03QSdPXbwvO93rKMlT85VCjhVeQXo+gvlQX3jI
NXZHfKLaN5ZQjn7rjHpR+yGi1IqY99Jww+9aUE5EROx8rW+ov3uKJy8xM4t1r9QKx5m+ALAef+Oe
Aznx/Y1B7PZ4YkGXJvU+ZC2raoEEJ4wMUA6S+I1lfKsfi+7tPje11ZeE9Zi1eb61fPoHhN5GM0GO
s0cm45LjozqdGy7K/IeUFDGVN7VV5KimepmQjR45S09+mrL/9bU78ePZ2Edrd91jJQoN6WEYKyow
0t/L6Y42IhVEeOIux5BJzyUX7NHVs4EzWp57HscKz6Xhj//ePd5hxaR7OQj7GfMbS534ldrMcu6e
LyLAbYcDyUILjhcS2JiSVbqNdJNjGNeMZWWrVpa5kY21f+xuQlsAgnabaaHl3+IpAEdXZQlJgQ2m
Wje1AtYkhuNNRnCS97Rg+jLfKukbb56VG4dRcC1HmJDSgnkAM3XI3KytdM5fO8+BPnw7uWM2pBTg
p/mYk9rhTwXv+5UyX4UkH0BlZhL5cbO/8fx0lkN/IJVMyhirSbbQvpJdbIqQPNO7BCd2OAIfeYxP
7omPPOKmP/fAH0GxEjfCW7mBQcn6lUyVOpF8N2Ktbm+pYiRFFWuv69CdAin8yO6IhqcOQ+0cc7OI
76sj+2xCPu4b8OWQQBNmiPsmIpdpqk7B08hn+HIPM9lrWjr6ndE067Q/DEQPLUO6A/VX+x8FVRSF
YTR8/rQy9+GqOlkUTcXJkMyOlrwDjCt+g+Wqow+rgcX/PL7z6ya49pDbamyrJAATAEnt7xvn83/G
VyMg8ALh6sT8YoL1lhwqmDnxt+dSXyv2Yb12j4iHZKPSoThkBlDHwbOLpTensVWh1k8C9qrcE0bq
zbEEdVeMdexXR/CAshpqLVHaDqbnCvZPQC+kYm4KQ+HNRlntoXw3k3APirdIHk/lm3Kz9O4avhny
QdRL20sl6gjfntyO98MGT40v0/nivKSw1UFXgKzi/ti0UIbDTzHmCZ5KppqH7jGDZQLHNamWIXUY
MO2JDqAxIcNWsW8pIkw3UTR+qGKL1gtz1093yir1lAp6OM6eOgBy5QhsDDwPI+tOfENdYyEH3iq0
Ur3dUL1VQ3A22nAChCPBq4vPxIBjI9aw013Uc+pO2ZbnMV4kiRefo13nMprBsU/CucSgOWLa9E8I
EjMXNhTQVRTM4Qg+KY7hNl5/Cvh2fjV0dS+URTV2wGjIwzliiKoaSvsoPVynbQQIMUkwfldOZxdI
o9KY5eCAyQ1pZsiYRC81F7MCChARi5fBGNdELpTQ3yrmwHBsKjBNrfRa0ByKDvcKLpAL7oC+g5Eg
ulgHXKD2Nqvd0Q0y1dFvkSWzDdC2VLq+luYSwcbL9rT1zoDaIA3mb9s7Yz8vc8YdQq5E4znHjPrg
NY9MJmNd7TxwpiEDB8Eyt3L2FdhjVngFPHwdX0rDrgWGujXutEKNf9bkL1mNNNElizAb1Z0uvPbL
ta//AdwozCd6rJQH0gOFiXTmGDwB0GPO3XyrFYGKObPe8vJMTKQUZyGDbaKm1ihF1oq5sUf2N/Ji
cWVUmuhjg8BEdO5d5cU0Frs5y16+m+M0eYLNRAHaMwMnlr9Tu93ZUqME9pQg+n4HO/DXkMlPS3Sy
U50SrsNt4obU4qAkGZAD67l83XwbqVnZASuF/k/aj5Qlegv8wVr8hHBKJ9JpDSUu56bFx3VA50eq
N0+ClxWiUNidOKMihSHIpWMc3MBiDROjW82bdT9NR3DROtWSvgC0DoER7j7zSIn3gj/oDvSSO0V2
l4vUoQQve/oSDTFgWNMgEc3tfSBUA4EpxgFhjh9zl3r9hH9s79++henkmpIwCcXZYPG7VZVOjgyh
ibfzARVvcVCkzV5ceMy/Hn65muIRknK4xIw27CoqxdZlFrI+G8zjjR6VEwLtLnNebtvrn0OTErn3
7xNQFMXiP5NZZmxBYTzWHkQKolI/TZ2KQLVTGEMYUn+tm83kRM8/UA/LvOtg8/uk6PtOzOkY+/qK
BkYeIaLoS3cC1MHLo+52zH5cuB0rakw3MCXR8E1hjuRVsNh07l0o+NiEBLPSzBzCN190U/8dudAJ
i81CmAUvCbDBuLZmOBAFYLnSxQQDxlWBV8z3AsrCAVuTsrkrOJDcxpImfMokVPShNerXAgAlIvAR
ec69uHX4Xfo4wUAVuD0RJoeP5+t5PUIPDyGVggTkijoRMFBP2G1D/7y9O+llGDqUHJKKeRdJF47w
uCKV9KL6eOLxTsz80p5VBi8Ije+a3JPzKUtVCCfv1uXGxQf1kAdmOZ8PGR8adQXLowbcN7JBQ49d
4BKlVsGT/xgIQ8qIo+a5hGAiN3y8dXpSgUCTxKq9hwJdeSi/I6LAAZMXUwjP1u1FSaag9Thwv7K3
Cx+vXvJXqiMEp1zQx4vVW2pJcLSqKOc2gNIO2CFmtCchNba9IGCNX5HpuLqR0CquZrnjRNCxRwax
LNfOrkFQytzerpeutdUfu8oWRJPpRY/+niCkqQjXpq9tFEz77LRUT8tydMf4WsdHZ6q/KwNAWyvR
F79UF8y8B7UlFUd6aYZsUTqMXwpYTY/zHO/LGO/Xs/OIIrt7GiHUlWfha+uCO8dTilyv1QAwQWeb
+6hBIBhXihaTujCVT24md+w5sIFpiI5l90dusIAKorY3SlzXpkkMbWCRk/E6S7twhdYO9difdZxH
ow73jzw0DF+caYNHS+MzkQe5J5cQGSQV7/NtYbHg4Fl8fXdxoZbms0akbkX+qP2+W02EwHlKmISc
CU7ywTF6CtQvkA/iv6loylvS9RaCVpxfeaQXmanPelEthkXYdjIdL42HFL9yimYRxplwG587EXq6
KJ38wNiPFXkThhWj6BqFJ2FpfAUTfs926vQmO0cHgoNx2eHnm+fAwzN5kBetWcmdGCngJQ6CxSuc
3N/IJqRwEiUPUQttEEAM0gjy/4FWv5YqzNvVMHzwAytg94r6wgHjQ+GQVuxC4uHYfh2iaLpTY9Gr
Ft022NaRg+PL9GcRDJ567KKk9f9qs1FHXGUS/0rMB0fE9OUu4TOsLU3c1Zk4UoSQwhdM9OLDwp46
fyG30JQZI73loMbe3uVs0jd66IrX0qk1jX6VKQMSAtufT5iWV2PzwOsUgnXvVOCmijsl6kZLBF4o
JL7U42C+mU/pwPJT4qcSkt+LcJB5HqXTdQn9M1EYCi4vDlF8ulD5ITa/z5+b1+kFyHNuWP+hpmcP
bMjejDExYtQL10N2M868WqvSKx8p6BrbKGR7AodKzup6VwS70aAshNugdjmYzw1rXRUoCZ9jxeqJ
swkjshubeRqaQI7s8w8Mmccz6BbaE6ppkHxpEnAZpYHRsqw9UrJKGaiMeNFc9L1Ll5RH4dT5qYX0
WQRboHTppzlWcOfTRPI6R5hPTCv+NMrvtwAxGojqBhGiHz/j1gs7tab6wUyASfLQFzwjvTJBDKi/
lsodTFXu+a8315o2d7t5coVqDpQkuCSbfhecT5rusFZPYDl3lz5nxschquVNlh5mxr4djqY25fLY
MDvzlkAQmA2nrSc6kiPqkMEjnvsqZYDt/YPLHmfo1LCI6KRAP5ohFzWKXvnlsSnbaVrFsgJ8GOlY
6TinxOfOO62Ao579+Ib2nWvFAI59lsxSFruln2uWtGskhgShWlN89d1wtTVlf1UnbldsOeWqo5Aa
2uE/Cyh7AfoY09kYgY+mV0I7wQY0uRU95IHq2Vcn2yHXo+j/0EtfZK426+1sGG/B9Y1UG8+g/vbM
ETQqn/QPgJ/rqMtkoGgPqbxdKkiEcNkPWz2G7TqpvaFEuGF/ZnSCqQEO7fRnWKEp3YUBKw/TLpDL
Ep70dBka4rlLQmEFYJPEMKd9J9XlwOkUpnqMpCLCLqtdlfdW1BKuqpDq8AF0dZeOPg0FMAwW/mpk
j6zsfWa1Lrwn+DTRh4wFMdw4GiEXoEWxy2NhvrMebdowmZWFlphqnbOIi/QeLmL74kbkTkoKu2f1
keCzbNaYuG00zrOLxqm9kT6hnKfkcw1Q9Bb8STS7+adp7/K+mLmJpqGOfJ+4XxtmrQ25vHtmr6l+
8Ih6tB6YlxQVf3E8kud7E3okTd9fQwf/4M2B9VRf3o4vsehx+/DpTxXUzMO/wSN+4WtfRyYwYIgV
t3B5tyi+V5tjOKmN2SRZ1pwG9uImzGITn9Ra3t4Ts7xhbpdZees7daMLCOykTHARAEEqQT89kCog
FfjvbqYS0RxTdhFlxFYR/KU4DyFy3SiA5+ctgcLlO0GQzHNHFz9k90i1ZucQo97r4GwsmcFzbhok
PICOezGtJMUWzh8vkoJoNZvuIN066A2V2VNyf54vQxQdPqSbgFCfQMmMbCaJaqkE4EdxSJtQF+y3
PaosJbtkSwfH03v0UOvjrNlzoFDdD361iDllWs2jor8mbhT9H3ZrCaxqqsk67OrNhcHq+CfVwP4l
FByYX8p2rws+djWwSmNfRuD3c2udz428oKODi8bSodk7oXv1N13eLdHPBRDqeDJYfn/ymmm1N9uU
cHFwcvS5fYftYM5C4v5YYty3lphgBIGOdK0zec5NfLWr/XUdG3/AaTePkT1s6povlc2ZyEt0WLdF
PHyr1cxByfuzsiOZsQHNFVVqKwC2M05LWR+QBiYL43r67tO0hZvwEfAUMImloO7Fgu0Itpxy4sSW
3hUH4uOWHUEJAYscJas8AY4rdW3yyCaGh7ZhxZe3vXypSOUK4aKKGEF5D/+sEeyGLjXYA1Cpoz9i
ISLtCD8to0DCdoPfIbMH5qWerXVEGKRF7mkK8zgalqFZB5/B11dyde4Y62K4IwZ5PunKY3wZlQ6i
aOgkFdKFEjWNPD2kebAXwuCzslGHvfo/AcDSCGezjjO0GJi/SmBe5rZ2J6mSz8kbdiJkKrp3nIWq
tlni40GzRDRhYQImiBheobgJpSLWoWWhBsSufZ3DjCO85o7hnnlzaYmEIppz8agaMxwEVcaAhguW
E2SG9p+rOZSCdjzPWGtZrbejLz81NCYnlgXUO+riptjZBzg4Mg1ZT5XAxxoYzoeVQBp1e8kj5rqu
cxJho44UqGsLSze/dj1b5C2icYI0gQGpIUW3fTGuHuRcA93rrlB2PbuQ5VCe61chdY4syU1fBiG/
yhYX0JJ4zEYeiDtpJx5D0dVu6DrU1z8x+Qfw5N82oQPmHZhWgYFslo6gDbN2GNE02d+79o9dDi78
mRoJaW4YXZn8UWMb/FeK7U4OB5npHUHiFrwIQ3b0Y34O/XVIK7l4yGoCbFudqOPvqsEbhUviw8Rc
L//I/WVr5ljEfZM8oHW2gXPVJqeDROEbWMYjvrAL/SpJVi6S62Hv5SBoiONqbshr7AJcLp2uxhmS
fT0NtChwQC6UbtTZ2KJ4WsetkNhSg6F0mS30Lia6lFTkhcX0m9v3DsMa4qYKycfcU4iElsam89LZ
rfCLu7zkrR1KLicP9p09aliM3OFgmvKgyH+4JwrGdbVlY+oQBG6o3z1vy3Sdttw9kNb3LE5bNI71
dC753TJDLfdU1ka9hsLAUcpULIRNBJhkGFCSleLM4ZbzGK5yPnr9jONViMEQRXyKrdbiSrKq9xgd
E9DpBE/EIvXrzVkV+cdpZUDqsuspZxEli8z47+yVyt7xNSSw17jZ0O9tS9HCzljFsQJWDMdl2R5n
55f7bUkr++UrgOUGuiFTs8ZHHrIEkzHmJZyp3ejzBSpKTfg4E/DzdGc+h588U4bSXEBP3+dPEPSt
x37hC1TH5WAmWSp89qT0gJk7kEG/COAJGdc6xBLjHzwf6YI6tC3SNShNyvYELatcU4C6NtcbVMLR
afdT41TOtR1tqV0DGZs38Br48JrbqwcRKMcNiTPH0Y47iby+UgbXLk9lBP1VxrsfUrRNyD7zfVgC
Z1a5T/72rtxAIp6WUcCXNf86FmR5okY4Z4xA+/gOTKYR7EqbziNJ6jQDFWfNppQ4N92NcDXLwfKB
pOATu/taOGpbONph4QAj7LIKvMWl+A3ATqjpbn9c3CoLY6Wd82eOw1iLhqJ3T+TPeH+iEr3PWwzg
U6oINJViAdre3EoOrlQBYntaVK80ld1KtVHGFZJ6P5JulmVIsi/o6fpBEzFF7rxBFwGvwhMQ3l5J
lITL/QD9eQVKbZ4BC269LhKCzbCl4f8bojmfwfzaVgJ+h5+EL3BV9rtEK0r15Kdphn3Rfh0u8LHr
CNo7LmnVgivAruGa6hb41xR2Wqm3zuOelOZI/S765dU2wRtal84gVugkfAqBx4gts2HuP7GadaUh
tMfEyq0zYPiWPK+xyI66o27OBUDCYz2U4uJk7FFKvpSLOXuBGyLTX0MHxIJ4F41GcQME9fvxC0/5
aeVtENGRhGDDNNh6cohsKAcEiwiz3d32gaGy3gJgtirOgeOCKJzAPOcaEvf2UM5tuT2+iPfAJOig
A5q4LPA2sfJEEWYpRgrHsMznm1kZXSAQ2GpAaGrujKcEcuItvnZMogwbUwrHJWzFgB9XTiAPTb2o
ZNGc0j9K2p1UnbEEt1uprg4IPfSkaN4V/JYGGAFgbIxU7v1w0O4iszIlTMgDctpIEIWNkMWaeEJx
8pVBeSqd06hYSKIkoBEe4lu+1QGoMNSbEObbreUzdJEgXjtTUclqu1J6DIgbqzW3OhTFrq+/c3fu
uWr/IkWyJu5qc/B++rAA/Rszrkd7TSxjxiAKcLSByjFsiaPGZl4VR0hRkNmPdH3bYcHcMzswIA0Q
Uk8OT4Qh0wCGm6BbxNO/JZer0LhyjL4xn5d9HjXroVFOvVqos+/Lo3p0SqqYJknAj595/YH3IudV
H3o9ro40MeVACYK0cUbXmH0pFMj8uHieIJaH/gOVrmycKhXUsywtV4PZ0i/320jxiYtmPnSqb3Pc
VDgRfAVgDTdmD7DQ+TK8juxbaYch4COXFebjAFrEktA2QUEmVRGRaIJqbKpbAEz7gz5NlVRLq2E9
M7CUrYJFQ2jtRgxOtdKTPW8/UYkpjuATE1mJn8RCa3l6eMiSfY6mW7R0rSSDsyqPDeZAjft7fha/
cVu7ULWHVOJrp6z9O60cxSybnaa1KmVvakHc0CMnKaavEs/095vMxQ/yOJdCEkgodanaO3kAta0Q
6kvP7soDG+8aKd3szLhpxKQkHA54OEjuZHQaKpePd+QHttEcnEBoP4A0lZ5wVRgbLOCCfKiQRuR4
mG/Gld82Utq1fN4fRGf2kEqrpQyM2VsvH2KW3r6yFCDKn+B5tgdUs7kTT7Z+Tx8GhHhoCtRNXUAY
6vu8qTDvP5AM42nJqI6i632Kcanf1Z70bhe++oZNLKpMcijOgZfIW5pXO4YePJRxUs8X7eV2afH/
FDGJyKXmrtkUUGqNyHaxUOuPSGRZeqDx4OI3JNKR7ySGM2ZaiEm79/NFfR9pzTCwEpIpQt7nNxCB
4bxA9tN1K/mdzIjp/SHJ+zHrJyMWsZjdCNHPRQW21TR/D2XKDLR2bfw5aX7aeBH7iLc1oWgooUXi
3w43ATCNlX5Bfc5obuw5pxy7FUa+isO7tPkeOqzO1CbawmLE68h6YFMTQlA4/FAk5mMQKVjbsBUH
mX1r7CwXnVA5W6Z046KBSLdsSTDJos/RcwNA1+mD6SQJT0Le8WsG0H0LhAR9OXXYGlnxlyJXFX5D
qUdfp0eOnJ75zkNrT01EuTvD+ZicU1Tbx5u6T6Xq6Y/HLfjPDhPWDJfBzEzDyC08MmovCvwyyyNg
B9/nUfekShIMdrLdog5sTzhR582IdUu6Y2Bx/c3rbRcR62k16C5u8rb8jQ5fm5LvX6a7QpSdaRHQ
+F/KD5tCaM/hx0jD6iati7cEQDNFzTLLzHEK0DzLplPOmdz0Ixzaz2rUDSYGTnr0kI+kWoCCxGa1
l9apfZudiYZw2mCPOKiR275El4FSwFdCAvk5iMRR6gG7LpJDvbgpDWE6OaCD5jfTSqnLBFm7bPsT
DNL46h4SB42xiRr5uAcoUbFB2h7W4JFH3bQ7u9djJ5aQkjgc5uR55QHeGPg5n509TPYrUycJ1FM7
vG9xH7eNL/jdAXT8UHX7L5cDYEiVF9FzMEbpT7QJWwDJ1k3z5TuD6vvi9iJB5JOws32MxBJ3BcGo
sP7P+9OHDDFCz16oZK8nvPb6T890FQm2mjZp9NcAYzJASFAPL55b284yOyjy0qGpQ9uSPGUcCcCk
TiQkFRK4Idy9CVX1qE6fRdLdb2253S6+dTEW/kNFEttelldBZgo5fKvCKiCYD6OU0JOVYmgWp5cR
xnTNDXcEvCPIbADVAFCuueKP/UVsdPT2kX/TeAmB+75nmRRA8FYYf3SQqB90JHzeUZzlw+Bi697Z
wPv7xcaHzjlMnCSnE9uUlskfc4+vzF/I9eZkmA/8U9EKKL5tUpTxQnLRRLvSjNlIHRwKTYjwjSU5
NiFdn9F189r22N4wOXM39IMfyFS8ysvBuCZRyUxPITJMYyMfH8Pa1fmuqE10gG3h7ILZRzQJlqXg
ABmYT28pKeaFYmiH4hEAhVqKcW4uOiLJmjqvpSEMZrxqr+gd4aiy9kDtYNuuKacZ0CQPT8IY/Dk6
V+ZfovyoXvNQ0I9AHA2UD8TSnuazTY/To7pbAPzZ3UDLM2ah4dRwsIFxM68GfNGbNW5sJAnLPlR6
R+Ooes/WVF8p9RROH31uoTlh/4nh2qtVPNcilFj/A/YTtUvxSwPvoqIctffgCIcGLYMYE/0wb0gU
OBd3aEzg6DI4AWRHAvEVE3MqWr5Ci0gtgxmTKCoD+xWUISdnI+1qwW6JDYWH0ArFK2omD6igbazD
JSE+swyALwVR4clLrKYVsNQhKpAdwp+U0f/WJV9suFAEsDceG+pclCvahGQyZJi2enZiikU2hEZ9
AUDUv2N9FG3KKT02bShsflQXkJtIXqTHZqiWpqAK56VEkWqVwP7lWtgMWFqnfgaA4L+y3pOP5UWz
vy9QsAcDISFD/X707caUP7nfCBpO2lKQ3nevSu5zPuyOAOP2195oQeihaZnFiiV6Eu9MDrSzsY6z
XBJ1H9CF70Dt5V74TNwq9hTuWsPWtogZKPdvnWaraC6FPFWModMsvlJ7iebAHHtBBm/5Ovkp9qa4
/fUfCwghxACcovoF2LTZtObDfTdsTKBr9BlYqiZv/A9yzfV88dCWjC7At554qbP1/SQrL+WfHUsl
v7wd5dBq5LKIHsK2EK+1YFPWJ/aIrc5U9+AgfM8HcMF7BnOQXIpYjehiFiux3oFoUIY94BWMRDcA
OFXZcrpS5cRg92gNj4QVhnhTiLSKU+vCHJyClmdJeC5M26C4ziMJHFmx3tOx1K8XAVpfEbmpoC95
P+SuqUJlKTWbI4tVEP0pEbUj7XNY766R++y4sPeO6KbtI7v1uUInrnLyjeUrm45N0vwlpjOCsuHh
P6D+O3L1L1r9ViHCydw4fezRO/c6N001d2WcCd3HSUv3wgCVP8UCSg4Ka6zRhDo7uX4W9Kx3ARsF
TMS1GG9Y2mMFnh9zA2YPOJS+JJkCQKonYdfROj+zYX8QSBM2YfzU5CgL90gJadTX59l2Ss7a++fa
IKQKsvl1E5wITEHfWFV6ghXjzS8XAlMUX9u5jRDE1ez/5sSHnSwb12v56kr1w1fXaZcFFRZiS82J
pIbhSHvq7CsXeliH4XMX+y3vCzxl3I8BjqMEgG7qSJiYMb8hy4Bh0nd3SPJGda4swZ+yDGwSkBsO
8DcEX9VtCRlfFGbe3B/UHJdB5pm+o6B+Nne4ArAwEO8ChmE962eBrqu9WGmvaqiGshaqcywdP1H5
/9vRk2FzObrh1xF8A5Kv07kJiBGnsj9+LZy5uSRaUVDScSE2Zuv4kyqfOD9IxxfzDpM3/d6rpKQJ
BTIa9oFBjSyjYrcKhbgGQGJOhzN0UP5TKPGo2FIqjCK8Gdg5YrcRmCwNcr1iS1z5X1TyRPDedpPZ
9LO45l1DhIwQszbsQcuYMeokRirCPooW7DcNCdaPOQ2LYkULmaBNvBx/lMBDJXqkpp/WULccf5qZ
3xBRgIGMagj7z/Y2CLOXhpvx9hbh1xEi/CkfAiEjBEPY8uQ7CZSP/XWLFT4ZYoGGt9xo3g7xnP2G
p5f50hAd3lG4JoQhzUA0lY56MtWBxQUECHMialNkHsSDjKqsrFXT30feznjijO41gZsvQe2bEHit
4Bw6HAugoMNEPXcRDGFG2hyykpEK1cUjVFvVe3UUKZUBT7tM8VkHJY91Do4MJMS5F+oFuUtlf5z9
YSF+JfJjZ/d4o409V33A/y1w4W+zv7Z1qxviAKPMY/0xj3wTfBhBYTeHViw2VFvk63ZGLdjjucxI
qM5+2Po+2Ff3qEy0KgdP/GjiHlAEflGKnb85k8frDThKUolYYoEaOX2UBZfvfcoZXN6B2V0YQTwm
wdTm5DUQjh6D7p81bBIx3WhVKGb8m3Vpd5HzXrHnMYlthheOGsph1WoFFSdmtVXAADNGvUzydalA
NpEUzzIhthVji4YJujKPC2CXi8Zk5HrWoARgeJXgfk5YuJQiMcSpSHHafO4/7oiLql/WCUWxbtjt
PHvmeC9gzf+hDwh7znxZPJk+rjx6DePHeWyj3zBHDgPv5DuJsO2xvBOJ5tupCtK0drfP1MBwmseY
8j3OD/IiD7M/LTESEtMDedcLs6cVHoXD1fgXLpCVTXuO7eA1Dp4LYh7IsObrryPbHOaLpiEcOPe6
hnBjKdq4ISxGra1yonoZ4x/ArpPdH/zxs5N+ryx/k3fZi4FzO0Qd7NEgBPSRBFEzZkPRX+WAlrxk
lDOcg0G0zmV81ijAgaYOFujtMdzj+SCht/L/6UAM8rnq7pyHIDHXmCiYIHevjubpQi2bgYB6lQT2
JOEP9jR6yNVpODEXkBMpf+kfe07AX9DGRNC6O4nFsAfgsDHZrf3YX+s201pfEsLKzBzh/WGnfxlQ
cHkS2qCDRBIp0zMVGUwiYCg4rQe/daeI6JBDuRjBk0NIzl4nUJrKBKUhJwAo7eKLc851mqZRY+RI
+MNPbJxff3R7PCNuN3fRPZciogho37mTrmpokxOANnxbKuEbkpS4H52FJTIpULDWm9K2wC4RJ7kN
3qE1/WauTWeNdWTkakkKpjxAGg5c7/X683bhR10MIOHLu88F/gsrdjB36Jo01EhUeKfXafuVSDKv
I1I3MSdFvzH9doS6RvrjRvU64n2nHFK7Q9CmQIthtwNEJLHyhICPPWJ33vUWBqut5OqVEm2VNCAq
JheXYuqLpOoyZ33bmBpB6qdi+KcD5eHO0rayPDcBzduvx+uGgNYymxGjDPs9fason1w6VBaK3WUY
hMmfAihdnvCJH+MmWEsVh1zFYKbCo05boBbeEuwVN3kCWYGjaF8iNNGzXowFrpnuJgRdr8svSwtB
cvD2DtmrxaIKvshf7B3Y29aXLU/AbWCHm9ARTMqmdGuguXABWW0wLXfzPNTkleMGiQo3vwAMi6/X
qhWB3khirjuF0tQJGDGNiAs31ELM0s2yXFkalF5H6X7gN0X1G5Ki/rliBFRGZxOqqkM8k8Qmge4r
HSFtjguITi1eY/6se4S51ejZTUaTpPdtE0KyKKozUpAA2+wHqeqIV7ItRjuGhFtR2B5dB7aTmQzk
w27D4PRBNaqamtouiurIKvd4PDwzyx0nI3TPxAPQFAKJox7md0J3/20Gi26PsObSoUrnaftMIjnm
aFl5cjRtzaKKrMv/7oLJCGkr2FoF0kiwT/222xIWVmhau3WPrCDeFfTzoRI48XpwJfdLLFthxngs
ZUcZ0N2aOYH8OR+oVJurOpLiBdDZlEG3BQc5XtKB+oo8tZuWFLcLqQmSNkATi+sl8hEva2mMLNP1
o1oRboeH+mwQtQiuN+E4znNwtW0czWnUNiWIbdLQT9GIlJ8cf233jPd0LIhVEfajX+Gs609kU5xr
XIhO1UuFgVmuuIfrqo2jHEp1x36OZ/6JqZ297tXEnz0X1iNfqIzLuK71z1fFHglfHB/fyzaoQxLP
clYZziUTJbtpOugr4O8q/G0VQ/644po6L+JDBomL+h7uUm4h9yxExXQu7mOO+qNzoVQRgzB6sxAZ
3aZ31+CxyIZNfEwKBhjQqwl09LmBhQeEbe4p/qOWP3Sq1vpy3d0GAG2BRYajnl5huQgEXhiJyb3u
0hhEv8aawngtBzpmAneYT+nbT42ZEt8dM++B5F1GlEP0RhAsof4c++exFYNj/2T76CI3dd2wJ4lw
RX6OdUQsjXbGHhFSvg4xzzsc4mVblw6IolkiOgNY8/c8I2zr6P1dcujNkL7XIZBLhekMGXsq079J
iWigpi7zBoNLaXWNfPmyeyqs4IKrlZZPeFgMPMh4WqlevroFUOEGWTTCQj41XXCAm0f38OaoPWSx
IqG/KHg+70hjeAT9znMoDQJ9A8y8IwpO3EoWEmkNF4i9YINLAzWE1zMhP1UytRMeawrPYRnr+veg
IM8HSZy3LaG20m0qZVLAFSm9UZWjI/v9mIdGHMPM80cborTn6gqQWrEcP9E3MXmFxfNh1/fuAcgQ
cLvC449YV8ZS6mHgnFYqijiKHvEuTZ1x3pt1Zerlf7OlSwq8GuR5KGA29q/z/xoL8xvbZ+QC2e57
ulqvpfOWAAGDjpX4aHIPt1nVHb1qGvh4BkCPBcOkrBjpTbjf8IkqX0qXq10QxFGyMHshvWxhHpnN
wuV8VBQS7qPOoWYChMDy+oEV2bIxQY53nn2STKWjngR0fcAy62jlx8k6hkPVpbO8tint+ji9ictK
Un+W5itd7v9hk4kmeoF0Wy6Xss2SmQEsue0FIgeKKQHf6MjFWEdzNqcOUhrhR0NUKbyGcAOXF1wP
aG+aO2+kESdnd+36xELEii8ppP6HDg9W0vwp4svNjw7oczRqTvfIXhb1lFUHwmTl5fihvEmY3EQl
xCfGNNm02YEE20dWujPqlGEluazVf/kqT+b3eTHEU+KDPs+RxQ2JVPIJgED3TsIxzREy87Jn7qNu
RypDh3ienBL7jKQsrMBOZeenijmBqQOumWI2ZmEze2w3RAcNPTAc2vZBXOhe8dzP03R99BUO5CF2
8kfIgdfaFKqm95GDWr31tKchWoKpJCLR452+D7/QBSj/+ipD9BbWL362BWQeZUU6ZK079jjkOVrO
rCD7ZHOozO5+WFoUOukKmoP4QJ9xzO//pT52e8vSEhlQNblTt6TDWWu/knXcUmiMK82WC6LmlT7P
8+xdVGDcrpHCtQ1QwoKbWkJHZZTYlBYhRDzxu6jTvYClwEUv8J3FtoGmXOAbBuWxa3YBHIK+fcMa
u4TWbxAIhphOANC4dCU1gBQu/ITB96FqxjwN5HJzqxLiKq4+Af9Jq7waGxRJoN//0qOhPV8w+95Q
nVchLe1Z2Guh2SR2s3auCiZ//KBdqijwRnfVV7/ddN7QY7VpYeSmiU8/Kw9J/VvOk1z3K+vBJshH
ewKXz7k8kIZevjrQW3wFYhZ4PxD2skRrbHthAd7vys5j6UFnBcX67KZDegenCRFFfckjfiZdJvqZ
+3ZZxoPdiRyWQGRV7/qy2ahDtHZWnsT3+ynjj0fFYTs3wfhIZcY6a2p1tEXopL0+ovus5boPhHIc
NrLsgtPesGB2El00yPYL11xmaoA2SlovvrLNdakWCNI7l5TOnv47PR56rcYSGnvIjHIvSABefefP
7g3qNp+Ys1gvM7LfI9UzkgIA9+e2VEzJYXcKCAYmuZS68BqqhlZ9hryFA4kJt+Aq8BncmVQYu2oq
9CwY8Klvr8uKnl9u4Y7eMdgg7JORSBG4UZc11exEp9XebOdzhln10zJnwTYH7FJ4S65/nyI9bIZ6
wUCuAOPy1hp6LkFnQ0qPSxBlWe6EXpKCZshoLoz+x+dfOMkLuIzBDzhxoOKokDkGnkH/NAv4j6gW
KTClyMl9U6VOZXw51Vbmjl4cYqYTwHz4OL2OjUuhDjG0mo8hjcs8PTzIp3QHjdoM3cwwaZbxcLle
4hF9/fBDRrW5VgE/EmPGV+QO6fXjVHBMm1F6+ZZUfFX85cdz4ZKE/f4mM3Kq04U7iW+gNceBrm0t
k6lgB2z8E66vRpQaqA2ZvMtq+Itqvi3ruGGadZPx1oQp7Yg7NHp1ThRSL1iUDdL14H4aMq8OoIN+
50IY0xNZMVD9IsocZjxktmC5v/XwKZCiVTGpqmVZCdDaTAKcg4SYM7aZRl22wTm50crPd5GKqYb2
zHyCPo+q0ezofLBXzgwxHnxDSOWIat2bXtIPEbCPBkr481W4f8VhwbZy0PHzYzvYgRPp7v0DE/59
YPOzHCqk8bef/GAKwqp2bSXVkyll1vAoTzGZh3jyIVypzG1jsoBSP0jQl5GOl2cfomA6E/RHpbBU
2Wb+XTEsJZHARXWQb80COzWq5rGG1fErLSqHT40C7o9VA23sv81vzJnGB/KHt9v92i+mJXMS8cIV
GvVjEcyrjeTk240qIb7ZZQVKar0lAOOnrY5Ueh3o1fUUTT4FUPPIF87JfQ0R/AddYeJ1n5QyouuJ
zlE59PPNZrTljhBDVtiqWUpFYz8kBwxG5YA1EIfNyz0F4DK4x0FiSQ1WAY85lpeG3vXfoctVYSSM
lJ6gAawiVslxO3hUxM2javeCcjhuF1KJ/2TionhJoSw7E61ccg5DJt0uBfkKTOssO5HgggP/pq4S
By929xGX3SL7u0uMv1XXd/+FDsXFLIeWV8OvEDRcZMwB5IQksvQcOFRjQsFt25fNq2Fpgk9VD7nn
rlm9ZrSvgx6aO5vVDxKa2LyZlecRsBWMaYifWYlpJLLMeT8Ka5u3DvzaUtTdvqy0ToZwf3ToDcTS
J+4rHRCKFIAYuD/Lc+ErpGI01wFL1fN+NP5G8HRTwi8xJn+SySOZYGNLFtxjtOuklzUF8kiM8UQe
gsGXFx7rDs6hMDk7U+rLMXOhU3IEHHDN5Sfyh7EPY/Nlo/hb05OI89GFoOQlyheHumH3mKRv3A9q
lIPTyA9kup0MF5VrHE83b6oZKg4uG4fs0Hq8jFH/L7SItkL7T5HGoo/tjMyV5oCsfAVQfDajAhEU
DNmQsYEmpjn+oB0m+N406LZ5+qUAdM+w4doFuaHOiVbo+eBAU7BIFr7Jn/GYFyjSjT5HCp//UHVc
F1BQCoeSZ7D3LJHuUCcqtzQg8vzFWgfk2jpLf/C29RLWDtAJlMCqxlFnIgkevFPwx+vZVIuT5TVX
Dv6QXH89sYmiFdOn99B0VaUb3yvyhYYKBBtIWiC+o+aAD2qSHFgMlWavssmQ69DAVxvzqJOQlw+t
N4z/KUauAmNbdzeBsHPubAg527cGLV2EvbL2EwfvwEmhmpzOdCJFES08BKhRu/FaRSzgjY/tMY9Q
7hqefq1/FRNxz+5rd1ZeUON6IcbVXHdoJ6TXUoMgZ0qmmCb1zP00i3pmK0V8Wp7e4Dd75FF35v1b
2WX2TGqtO8h/o7+gJeMkvgndBDFUYINmIOS+14foq7X3DpdORzdc1PLPFnqjWkf2rhAhUcNwjxYh
cU3atVCxnAvSQJtFMwQ/Aa6XmWI8n2fJKPtvE26T7RyhsEidIOBfAU0ahjQBgCRCMwodkR4Tj+NI
gh2ZtOb0d/szx983quvit2GPpljJ2smTZPe+DuJqhJmT+NDHzt0x8WA0l4gzmakxJ/oa5Hj3A3M7
jHOxdP2UOBUlp3LjsK3RZ+h0Kpu744HqLAxGIaQZJbZerHg+6AoHKJmvVmmr/BM/23JxDQ/idtmv
1DO8HLDtyklZPtcYeZuF5lr9JviDFqOiZ4NAsqqJcMae046KyHraQrwFWp6SOVRVsx/Y2uaco350
LEQzLUWIIqXWCherHgFaFvkn35WdcN7qSlgrP6p2K3joiA09iKk678Pn7Z/0FWmaU/Se4u0Mdr47
qBpaQiX2qhKUdiDbAexrzM/n3atItGqpUGSoCnwtR42J2Cg+jzIU2FiQMLEgNTezKnSw6HkILBXv
cu0fk+9LCSWDgGYP3RXdeIp/YGqvMcCx2zQCkhZWu/vHgEz+H+hs+89vJ9YT6Y+pAKtE14NXLtnY
URJ9NsGaTfZcKwilWXBeEzjinnEecvTnK164wiCROnvF1AD70mJCXgtW2H/4Z/p/KNYpirRBdCkl
imyt8eQcgvGDBXspNnV4APT7tpbnHvLQgUv7+Y4cYNxnyR0vg3z3ywrAU8r4KzW40Fw9rCxU5AMd
5UIeQIcJy0Uu5xP1pL4dRNndmwOWYmeVJWa+KsxwgsdFfm63cjnGL8ESlkgq65EdT7gOaeCuBy5v
fmz35cXSfuima89X79Z3VvGL/PV7tnoyEFobWuor4Yzpr1Aa4dR2OE7Wymb/cz365yWysSFW6Gej
IehlkqZc1WNiGMvoMdAiyGg18+mscRgiP232Rypt7ULmXJjsI0KD9sZX3KQT4b1Dyo6tkw4iIYix
yNdYrfp9XSdScnidshlGSuoFb64rn9F9nPLKLkxjqXcjczHFwIsNWvYuA4Mjp5jcJXqRitLJ2weF
o0TvW5Rny1VIEZzYyj7nIF1VDEc+rZsAxnm74cVpIzWCYmoDb4YJASL0iYv1f7nPi3FclS3WjFI3
0rxvr16HT9xmzMYRXxs7dMSYwUnjC5JEEEB3b/UxIFEpmA1pL0B5O/PfHVtATciIXOtj1yIfUJq6
n4Nc5x+mTY0YIa2tBOLflnG/2sdrCodBAcoyDYqPwWLoO9QYJwn4+6LgYFy/uoo+rs7snJyiRaKl
16Lp1wbHMxtSOJkmV/k6Kmvtjs2oykwcD8HVf4nmsW/OrkJ74onveuKLXAH/hzA8Q5lL/zQBI8Qg
I7QIG9itlxyiNg6Y3VGlaOaJ+dOpsJd/zvGN3k4aVk3WI/HdiKdAbHVrSyIG/AylWYm1D9gY3+Yo
y+CIak2tczZuUo/FUxmfpHNejUqXisLpRBAQnoKnxFeIEQvuOc+M7ViNBaYwH+d1GyAKncghl5sB
Bc9sSKpghNoqxCf10ekmV/QhXJQT3ieRQLrs02U4DLmlfWse9lV6OhsmCun2LnfPU7i9gF1v7+uD
VDaSXlLTQbZymJuoHwX8MNnSc6O1zv/TC3vSVHN9gLBCtlDY+jucadQzC7Xh2YryKw/RUl4ADbxN
NMuECjxuNC0wO+ud/peQwBZCHu56VDUdew7weUB1ahBL0f39lFRIntIoh7oAFQ/I+Kq1xKiH/sAy
58dTSpRqphc4WmQUJA0qCaV9oqHl48cjzAArqwYhxGVy09PL482betEictmjAjQJ85L/TYYXRKAK
CkTDoOCYJwm7E9aA4sr9DlCx74n1yIlwf3jGpOxoajbcBia4ozGrDics6S+BEiBr1qmvhioq+5oB
aunFju/cmmO2rji4jTd527OvhofBX/ba1CHg+ssxrL7lWm3qDJNoso23QwNxY8mdNRSZaHPoJuJr
ih7aTPYtZVqSA8zLlHP7Hl9Cf3nPHXtLw0bcN8RZp02rWcqvudho7jWX5T2YQfuTEwenYZN4QYHP
jjTE1lAMe2YLd4DS/jA3ONshXH+MNxad3uuSfx9PDoiS2fwro7xjDraCxn8G+W3QOsPNIFKhCqn0
1s209XmWXJBoWoGuusMMK8AZD7bmGRAjT+STQ+hANCEU2BKTGdNBsZiMaXtIRbSJ0tQnFVQYKR53
k407p9siQd/Bin1BfwLyNlT+JmQE1oGHlaJ9ydqK9wA84NzEGmuxrpYVHYaYY6ZKHD4uQsMvi6lK
42qOcRktbNeEmUd5YdEo7udSrDsRSV/tSPLl57c091XKxoipT1Sx381Snk0lhOpu3Iy+2s49rksx
JdCTKbu4bimMwyqCkiaziTl28AlvSnPCE1Rb3fZVgRITe0Kz5A0LsuX4lLJn1S908cHudywCfGQf
3q6ZEYoYuildj7IciAO2oWXR04oq40QLpC2yxi/JNiWSm9ztM7R96QyNno/BI/weme9ChLCrURHO
njk0jWRRqndQ50iH0oRT6yJU0pl3Kywq9Pm2tUf63nOQFplmVmX9ix8wqm1qDlBVOfcrZ60bLOgs
NBbM1JE+e1kzmehAfHA0Pe9HWE3V4ca2hy9dG9Yg39NhA97JoEbVRgFtDiCz2Zg9xgMo2cBmCWSx
UEiXyAN0tzFBJvg4uly2WFcR/lWskP22vlbB35IYJ/C2IdX/EdkHYeSzNC23a2nL8KAz1nFBGAAa
0OYbUzvUuJ33JGNAfy+M7T/2zgmRcrfTCvlt+lvzPOf2RC0N7MKDX30VehOKPz1ejhFCLGf94Aoi
9nQ3RmZbTkuRBN8Gi1bvpy0xTSVJPTQTbcb+nOLqhykhhalHY+OKoT2zFERllod/4xdNpLji1MfQ
pABmnTNu1hOSqZSD7Iy0toni5gIp2LhqSqnTUuVus1+acCOFoYwwQVZdUMPJ7S2SfYjnbtbNs0M+
nqMWuIKE7ZynQG0UvKJ7zeeCMr9CwO5sBUUAeEwB/cdRKNDJWwHx1PoK89aZZoJXSCYgNstiAAoG
UyMyR7S6Nie867pn/L9bfWPgooCuwCadwEY3E5h5Lif7g/4+cyzt3xPLr5cPcqm9ssSAO3ED5jyB
T+frBHvjztFq5QIV907S8A0shxX51RZClsUUbtqA3UO8A9gNt6R7bpySFaqgywWz2mmEIRgK/9DI
xDMICFwAep3dgs2q69Fu2Zek9DzY4hFIEWa7Va6S5TWO+jMwvYLcwuFqzwZUP9P7aChz2GGPFFSr
QEcg6MOuVby8h2NMQzSCDe5VndJ3Os60LBfn508u584Vu65C75dlwfw3puVp9cmgw/gWXDpyEauv
hE7QTWMKdYUmovxGL37bdPu9KFgMIkSQobGp58R7kv2ezFr613puHI5JvPFYYDNcOFDj9hlYhYvb
duak/YDX1ueNB5e8U+xlRqLwxbppFPq7ioZv2VI+xhGrfI77DFVkoBoaoRGV9KDqfvoA3RC/SQOR
XKfApAWIIlGhJq84/Uwq2Nkp56k6FsVy70JGOEMbWKS0PPVHiy9QJe+SJKkYPXZGXSp676gFxUiG
Ue+gghDAiEKCp4xSvqOwUTXfNzEax0m1WgmxOUFt/W39OHGQ+v2XcyypNgptg7K15m19v4I/QN2o
KFnH27Rrs+R38QfdGYI64XGHOuR7He6OijMeteOmiFsG06unhZot/J/qxow7YbRicdQrmz6154gR
pOJdo4ZJanMD6pTEpx4lRzYVDKBQtyOSNFl1kLLHAPvuYKFNvF37XWKjfMXbB4kI9UNoOAUp8dnp
UNTkcMRTgfzgEm5rsMQv5UlfKh7S+b0y6n9YOeGp0qOfKS5wB2Mr1JS4elckLOFdXt6sbh5936xo
6uVAkUSEJkjOwU4bkZWo5ZE/ht+VEgrb/rAGFUzzml2ePU/41IxxkRTLCPbJwrBGjW+BV7oYhdu2
geNTdfLcs2gNkI5/dvpHfZSFBM1JOlMCTefUCux3WmDjIe8EuYBKyvkwp7g/8AWal+N+aWDZbPZb
P9GGZwrBJ1VYsuthhyOhM506VRzx7TTjwP2vDi8h3a513F6B29YN7EnQRsqj65A0ZoiGnLOV2VSK
s6Hor3viyLdh0r+EdJ/B0dcSMjNid//WwZOIbS38d7fdUDNqWIMWHuHEvaYUFoPSc+/8BJ2pmVn8
9w8mAvlBEkhX0mI79vQjgb7Mwd0St8vlOX6g4MfE0KuvTkfJqY1QmiXvKuCIHCaHYNZ0sU3cppHt
o42Veh045eOe2d/69KBH29vDYNFJ3Nv1VzNJ0rFSOlm4GcP6L66rr0KniRQKOswSHsYvofIfScOr
m7xL5etEt7zykVXy1p6g95uluR2UHDTSeXM7j/oVaa02DqATIVDJdR1AwDlWJjt1AqQ0KCkLgkAg
w5+S2YGPL5EburEKOxORq3p2iUzlS4LCN1ZNHrvSy6knLt/g3jjL7aifpz6r97zP8hrhN6ORxFL/
tNkcPfx0B7DHHtp3EdyG4+pBk7Du/SmxMFxqDdCtoG5eB1bpnLBt+yFKKK0plyeWJh1CoCXbHSaT
g6ijg9LqpWecJm6dOy1OJE8PudVddADOawE9qsFRsINHW2s91xYaEa1RZq4YT8vnfet2nR9I+5ng
PxvMn6l+YvBH+jCHG50D3ltmQawWiypcu/bfEMO0lvwVhgK8yzHeWaETp2KXHatSx7twXFP0nZq2
JxrYFzbg5YaADOAo7P4FUmyzcQowbfv/4lXHGVc/sJZHYh1oGsZTtpZi3A7BMY1WO5x18rih/CgP
kywxnlnioDjwNAT1ZZxs9nrdPLlgu9xIeCu4r1lZe8x6jYfnsp9jnnN+9gpNhnGFbW6eyeVyWsMK
dmqcJJuVeKb7Pt5TyidBlL5sXNzFOChKeRzqaFdA9lWaih0p6oyMQ/fztdqi2VMQ9O6zFatXLRTX
QLeEZ0tTHeondsOEkEQy0rdlNiZO3wOqNLNtiUTTX11mC6b0xeQreX6NbJ6V7MOnXKIx0tpx4Kte
TAGRcYcsceYnoxmE5Ms+hTNEfiqjPmJ8+a7l+WaHyz0zMaOir4dlMaUO8xCNwlD/vMBPIutS73bo
RN9K1oRu8wIYJWO3QJD1kWcjXJvVDiCke3kLR7cI3RLbyBhYCyCgYkYt4cM9OFX6Tjui0JE31evv
Yt+arSrL7KEV5wejH3JJ5F9s3unSfQ9H8hR/WVIb+FXp0OzWmUPq7EaqETjxDHTThrjzPhjT26jK
s92Thr2yFzqGf2B9zZbYupy/jFPQXXLWRp4XBXX1zrlbF9vuRUZGRXqmnPfE2Zoj3CeqqMsgNjJA
2dwIq8jCzh4ZDcUnHrARzQEt3+ERP14z/UCpgIgFexbBjyYYpIRIkybtoHrNDh8idgEZEwmkE78r
+4j792jXaZqgXiZ/CKHyO8E78iwl1oQkLkSJxKOvqvj+DH4N3U5tk12omPOnsj7vWEQ0QRLaHYEo
N1o6bXuk0AuUoJtmRVvQ9l5wDuUGoOzvgHUngc7hsZZZLSRdvUzF1EtjA/5qIkGMeXdwspjtpp0X
ZZ5VZoyiTxYJrdjvUPxB5S5A8qmsZHFSrvmLGxGBJOiqLohSX3CZ2a89fS8+zSK/F2sIKaWK3nf7
at1apv0vXyK6z3hdjGI2yY0n+sJO4lNPs4KITL65bxilImyJZ194tT9OlduS7+QhE2yVsu9Ws59M
LWEABdGHK+iyz0fc/gAjoSqZpc6FI0fLN36xvrO3Xuw38okcVqXjCDLBJVSGp43OR8twsGWzVeZB
Rn8utq9eGKOqS4N4tiH0YTZpuBouLAry+flHB8oNxxWjXVZ4MiRhkDf/DGCTHU1x2ycGWFq6C0ef
5sOlh9dWdoMBHAISnO46yQp8eK5Oh9hBlIo/cXTuG69+Z0Lk7EpX4+ncB9Yqf9PKXVq+PmO33Q9F
DGYfjHfK9s0b1PX7crgUEBteWOmJz/s1DZZ8XK7c2+HhvAnXEcClob1byWqGx0GaruucfC8CkvlE
eP/6ApHxPYOCmAx2m+JgN7VrI/DFicVbI2FrZDWiQipIrURswvgFCpPnqOFFb3v75Lgm56g12DGX
B2YwD1YEHp0sEgi8UtYrLSRle1JSzOPPU9NkD/+GceeCkGdPIjXYON+yoh+Tk7bk89Sec4YarcWY
1EE9pggGTR5w8z5JLtiuV1skcOLbvofL76LEVje0UhXx9aP5W+9XRyJ8/wiJl2WLj+yVg2dqnPlD
oQtF5mAcc8dugGTqrdh+zR5j/D4+ATErgH6qyevD23B0ixDiOw/mRYZUyM7xOlZxSUynZG0FCjjF
eZkNE1JxYgfXHgANONq+ik+cwQbxhl2XhYk3MoSIoSNFqK7hLuPl3LCHgI0WimB5tsSg3nlXpU7q
O2fbGPNSPtUEKHYj20tefqfR8+tce4MiCMoqITwW2FBpbbTILrPplsjDv7MWPquuAshqUy0EqS2W
T6CAkaPfFqnzZ7RRFSUIgHvAgCKpYV9HHi09jpm1AnrzVsn3pRps0Fs7Fya/glrnOsXVZaw1eVcm
OVJvT2O4icbCYPYs9hneEdm/A/0x7RiXSL775WvbJURc7MdkUAAuGnd5RqCzaPdjM2FQRGX6CMWe
lxOK7M4NihTWmAlJXTDHSzD1L7NbmoJdAgqBL5lvhXEC/CsTsio2szi2ymQRwA4gzJo635PFSqjD
mXZAAARM/mgy96/QHcx8ZEk5YMjh4pWLnw9JhF6tuT3YPhk09ZBpi3hUmiaajYzKFyS+LcCc01uW
Ow7pTw5wr2XrK5mkvRT5Tl3kQ1LfYy2S6+H2PVZZSbQ1kSVR7r7/uQbIN+afF75NGpKX4ThAjvdm
1N+smFLoiem96HsPEF2W6c845+X5Zd3L9utT959ET7PXS0p0m71d1n9W+92EabcHkAIB1ujGdGng
k7B/MtmWVUIvy6fw2pqp50HZSnGYRODA6tjGQJs/rVWl10LXI63ndpWMMyhsqQBJdfBJSnl4DV5Y
9wetA+2N3GqWVnR4/UbCDvEgWtc7+gEFeoMSACKarxCHPutE4rOHO1Ym10Lxn7MCMwMcyoTF0iVB
A3q9H9haoH4Rxki0NDSA6ZNckyyVA9NBCSFH/lR3EHDm1j2A3nGCaTfWLFHBRe4btv4NxS/WdRCY
IGFENY6tmXoqbt6qvreQTWzaj8uf1/lLpd3MijW4ePPGl5yHP/4jOxXR3ycytxAVYhmGWAQZ1d1Z
ROd6oUmdcGC5MOHDEXHK/cVoFnDkx8zU+Zq1xDBwmCFMVtcSQb4GRSlj+jx3ySOC4izspC7mjljJ
JQN4sMf06lTm+aUGoCzO2X7i5kHvTc+yzTPJg/5e3Ra05kDkLtRhvz/g8vcmPhwjoOUwpFQZY9k6
o3bMRQtg0siCYvyUC+YaAGO7tDh0FwFcubxug5joS4W0qwu03VL1GTg2UG4oUQNBDYIfMQYK5ORI
pBFVFAy9J6+fO1xGKK9WijjM+D7zs9q7Bej0WAz29c7kcYOcQosTeWHpr9wd3iabdF1eUzIsjg/I
+laQSsChiaUwSiIpekWYZnvMqJKq72n+QwfopfvknIOIr5pp6Isj1FLxgD/H7H1zsNc5GJESPEue
mBfAA5hNWFuOdsUPp/q3zM5448QprDb2UxDm3pTc1RaGUlN1rNDyQC2CcpkLnDMgI3gZcN+1iSqX
jksONfmHzW4gn/TCts4Tt+c/mahLwE+kX3AU0r5vrTzDP0I7xbTg42zazbiaL2NY6mULdhLkNWHj
J4e8KujA2Nmi41pYg+xcRlotwVqj9bK4Efbb6V1NRUIbifEBTIi3G/sXlFAGp5w2GUpsNNbHRkNa
n5sCMzlbx613z71EG7fdTAyjE9hs/ABYxtJnLZufKy4nQJXtI6yE+y6QfJbBKpPEbUXHlixWdDaV
vSFUk1Xj4/ovbqJZuokLs0O42fTwAZ5CbEakTU8DTU8JTdCJP6kRDwyAJvnfM8vHm5xFBATG3mk2
dkG/p28vcIYU8zW6h1a1LTlv/IdvwLUfiaQKf3mp0Qko2wrCFt3BGHARxuiqzHrYueWJ87ypsNm2
HauA8kBk4ouRJmbe4pJNoLc5wJLDz+Liqijb2pWzByTbOox4PGAqJ41jrRAWfnwqUrd9fmwJzJt8
j3Q2nMkR3kP5qGSSdo5Z/5VH/YH6LT5RdRaGFTLpFXLYr28Ky03riZh+zX3EmFSsO+MxsC+qCVnX
WMknoUn4woDGt60W30yawiIGycInwyy/JB37YCmj9mwC2H0rgqR0XCG7AbUPDckofLzwyW2HQqP5
HcbYPlPfsvXpQOfkhkjL5McsRJeYJbxBZqEnTi2zQn77ODz0RyYBi2xY69U4WBJWFSB3+Btv2rkL
UMZYGDOs5yMubPXeuOl2P9lyawfVnMZ1hSdzF9v/fAAxcPcZcwEBkHpuRZsyEhe4PBFZvvJVx6h6
3mKje5PcJOssl143xnoL8L+gXBxuy/lw2CH1EqTKtniXxKM1PKjsZVo9/TGQ6vZHWS9+Qnxk0hwf
2ek9BfeztRBXQRTIMSDNarx8LN+yhgf39NoSGR4WDES5yu12/f2cjJ/oXvlfV3p1PCxe+OK2fa9r
ZWuOCIl/ZETSVLBWBFG76Q2lN17G8L3+L0ySNCtczXjcS1/gCl9LsoFHS3GSzb20Sf6Pd+TXBbo4
EkqUkBR8bHcYNH1H2wi6oVXN7sXFBT3KzvbW5zMcpAjB6q11sH+Gj1XQEf6NNYgx/4c6bMOfk1gj
Z/FImrhCJwDqANeJDH2pRzk1LSfqAmZsXsekKLXUDMvwXyzREG4+IwzY8soDzS4yeIcFHMBRMqIX
v8KgjA6kdzXwsP2Sr7xAtZMOD1g/65yCdBE/oCmD+FWak6LdIJNibns0uP/n1Pvp0AADec0cSVV0
vrSkXztxukDcX/kg8VnpQxTVCjD1qI4tbiFtMrsLbjj8neVLhW9szuPdNcwNuRlSwmKMeoy4FN4t
yYqi3tdtVAsoFRIai4jDFlDmCZ22+0VfLSjXwF0pwO/NZQBWob4ysgT1Yc0Ezpks3Wk+qhw68QK+
MTvlIKefB8OT25IiLBZpUR0wjgVrf5nxjETrCy+BdWCicMi1TQ5F8pJ0dIhfbvz4tRV3HcKJE1M9
d9TBt+jWPJvxGJMEDLy3vD2GsB0Bo1Td2veM5aL/5SEaxU6ru/OS09xpd/cGkaYPZaBk/2zanSNg
/WhCuZm3DAAy5JFUzEh8DbRXnenJAPes3NHVa5OEYe9UoK6ysq6cTqerwDbPNbqtEY70gjZntRKS
cgLMNPhestFZOXQeM5p8dXoh94Mn+52UTfa1vUrApfsD/coO2MDOovNYOodYf2RvplOfyCBiyUPL
Jp53/WD7eQ6sGmpFFhVof6y+/ov5sr4QgRd5Omw4Wq2cXhoat4NmoiSZLW6w5jOEPFKeuRZFaDWd
6lftUt3c1Nv1cNLpog8d5JIzLgPJmya9sws6wRkH8RhQjoBWA4nENbBOYnH0DEbGR2PLisg1Fgsv
0F4vMb+b4rXlBhTCEZjvp0wPriTMLmiJk+NqV6YlJ6KnGwWTfiYzc8hBP46GAd9FWjSMpNByD0ZP
/gEmJ28jSJnw2kSAcnN12Jt+f/DSkp7YFFYrY67DTR42X9t+P3+OIbzOQE3XtI3aNPaXehHOVTWo
7sgc5ym+prcB0Dc9LzdQnEYQbyd5pMEaOb88jKPXXuj+vse2UQo7tL0MkSfsovidtgBP72JK6cCZ
rE9RfzH0bIuJSTBKK/LV9E6rETQsVGfOtVgPniiptUToT+hfqGzG4fQKP94SSlG0wmpuBIv+YlV0
ruQ3+dDLFet1/jtnVJ4w0xPgVutT00RttayDQGETat52X16Fd+nPzXItn97t/Llx1BcVXuAF7ANq
lzCQWoU/A+LdLoraKRu3s0oMyf7JzyYCQNxrWxQWvNaeNLd8QwaBDf9HhQdHLp9teZQNH/fSA/MM
yxkScqrVvpoL6jtbY3nSnFAGiPdPRLVy+PwHgnX5YyWwJwMSzYhlDNloENLNPNe/yhqcPJLlhMAK
m0n7HP/tE6vf7ZGX7EgijdXCvmel7se/gZp9i7GSljzVfGkLIVL0OzrWDGzo/oHbWTRJyZm2tQ30
gZkwcTK02LuxlXLuwizikL64Biejc2YT1PxzcHc8O++otUgVZ18gFm1QvS4M8gZNHIboZYExdUUp
eKctTYeeVH2S563YmRJyp4Wo6C9X7Ih0y9PqayRvnKfSon6ek0z7N2J4ljAN+cRxSNpVh76SxHmR
o3Hn0KRP7GjkTufL9EwN+rAablwvVWOLfaB/I48Yz1veXTrEZ+9ieywLbP0EsXATth8dqQUmTyuV
dpi6tod+uGfRh1Y0P0csJ9dlmU5IF1zocNeEtl02wttbbJEQ4pvxpJrZGjGp6YttUdlDSdibyyBl
sYTXvKVZhgPicpbT8oVjxyat3mhgjav1WScZMLWY5hUIp9z4TFwVfTOe9hG1AM39ZHpJxFYgdQ7m
ypLHwfgZIYXr9UhpIKQ70Stm2dSaIGLNQUDIxkAuUyckNrQyOreHIHBUpd1Gp9mRS0PD+/uPBiDf
Tr3X4XeowmrIb+s02JOl+USVHi5q2jyEZ2DaKFX1bhsfcTOsphFcNq1Jb0gICTtQwRAKHvuX/ARy
2EF1eoqR3u1h7NZtir6dxJCTJ0ei+ZeLz38v77xUc5NY2qHKhX4IEZWGRIFYvxGlakg/qPN9SYsk
s8eg4Upnr0d4xX8KJXdvbge+U6JROO+w0Pdlj16jGpQTtk4n9GOOv7UbvG7urOvmcaa3s9jfF8Tm
aoyHOUxFuWFsHERgGnLjQi5cQ74i2Q6nCPyH3hqVx7/G38vsz8QVcMwWge7L8nSVEYKsK//GRsk/
f+3OzX8WXYfwHAuSloMc7B2txBRKo5X4FyyN6fuXYtDohGxW4pp7QQBmTwJgxWEvy/wxnC1pyZje
60arULEKgSYwCsDXeDax+CKvi/4s3YW7nrVFlp+TSehbiLHwh6oKHUPOHClGDvNUK2Zz+Icq6e5S
6Bazxqlgkd731OOs1PR23U3p8Yv7Hihh+iLqJsG/uxqSMoXpJvJ3bBNb4ybkgKse3hKhDe4Hv2Xg
w4ZzHaC7BHJNUokO5mOVMSTe9BZB2xmzJNGsPrKwkMpeXP01mgAa7k605lrlAVInDAUGm7PCXRl6
8t6WiBWe/rpDiRQy6BSdQwn9picsAUp33yuv+rFKHKeMQiuj874QkZ8ujafcHkytH2GntOYRVzz6
JtnyM1YqFivDWg/bB4Vu88DSO/r/THyM9d+Fng5r1o4IPNCr2cGYqL1UplAUHGdL5+PuMElEBWcu
wrvj9kD5b0MPvZXMgsgzHUcs/xxSoGHOh/TJMVoPxSTaL4INyFJ9Xek0ihJxJKTXrx29cpKIuJAB
8dUdWWTDHXAJ9ddwUJK29MwBXBpg1litQmnFgxA4vPz88EOzk73xySCeg5ZASBlnARtfUOPGdr41
cXy9dRxry5Bd6tcSpKUSVE25VUiT6o2/lgvYXDFfoAyGUi059TLr+j1YBctp6y73z7P3LPGwM174
ProV/halJqt5wLKCwwrmZnYB6cJT5y9kR+JiZgXm0gS9xB6lZoFiGh9qnshER0iK0fifyBYk6Az4
KfNwYymqU6Po0MEp5QaR+q8QSy/NhKCsEgHgIH4TxVsfQlOTOEFnCzfo8pbhbWKLOGLGfd9StNc7
JP0b1gopmQYScBAhY7sjcS1Lp2r9bzAc5Tr/M8OLhVJsWSUaIBNJOJTtVZQCO4aNiQmmD6DN+n8a
zi6lsIPX+/HiLT8BmBLcHq3LLEmGG2LxZ+EIxXdBPmQMFnOdBU/aZ9VsYszvKOStuE+Uhw9CCcl1
2QRiu/PeQyY1S57jXsDvj+B5LViXI4yqppWcv/BeFgjopBq2DNMP7OoCvVSjnVcseWRUStDY05zc
TXsmeXxLpYwfJHFdQVqj3gSjQAFiYWqJc5nXg30IKumesbiE0PfhnHjS1nOpY7rmVtto6MMacxZs
eS+LZuKMQSEy1mfRbjiE7DUUKujfDW9mvS4WT2gOLG2pLEFC9Vu1bC5fe+IsO0zWI1lJlE8CgLiM
ZLIuR04qtVEq2DOqZMoPiA1GCQTwUIK0dEogeTuZCWtzlCaWJOnkaoXLX7Og/GQphCB5/jpvZuAS
kPjt4Oc82WD10bEKTCFrGATuNSd+FIHvoF+BU0X0Z1b1mQIlhyR5LSmmgQHJKDvXMIjYylkzXCiy
tFmYhUcmx0UG49SxJAQ6ND/3HKYOY1ve9lnPjjZfhhsElPlWT5qGHijCLLAdmJhQsYdgG/zob9Vd
sFLh5gTtAT9nI8UfUmMYAqdvx8chh2RMQaJm4Z4ivtiq0p1F7UVRXkABBWIFMUwTEtNsbINI+PPx
K3BZQeCDcUZIt7Nvj7tdowvRdNVzjp7zoGnwtFHjGBWlbDRcw0o1wHWhhyHgJwX/zeaqHLb3aYiX
B832jpBqxoSfyJzthOsGstyy5xVi6M1HE+fLj8I0/VV0xvoXNIro9DbH/vlBAHlt4qqV3l2EamDc
+QI9lwn7hdBq24SEf57J9K8fGnJ27ZoJEFiRdWz0MNjwaHW/47/GiKVpN+AYhyGLHF63Pdw6msBJ
HDvjfUuZDuajOYL3z1gYt63iB/y1TttFxjiiG+ADV3EXwNWGur/mBlMdj757IgBKjQW9o3g5ga9f
MznLnI6PnL5Tuyh5Gt6Sghhpemqvcb9W9bcRnzjN5q3QaS1cFbPF1J7hcIbIb3rP6dMmX613ZSNV
hzTEW8NZ1j/1LLLsLDXuYzR4cr1TYmUYGCigwR1JlIzOw7lOq+qhVd6QdA17QZRA+I7PYvkwzQPB
NkhagKFG+IXKgB9BXWU6bNsvITI5wthVW/Wr5bkJYH9DCB+O3CeTk16pDZEZdPTgvnj1OzdZ6utf
yzFuVRmfOSPduOB1GirGZqGywl3ZSh/VxCM1G/U1w0C8rnVOGiqVqVk01p0t8ROWphx6GkKbZ8O+
HYFJvMLoVDOM+qWQBM0JMoU9gS+Z+lvPQKWFUZnXsxKcV2IFAfNSZwEupv0ZCnyaAf++SlI3H61u
tXIpP4Odk0RGZYioRBeBqIbXi16DEtZJMOWZ5gpHU03v79cevtFnEbYsl8++WRZLVC73uOAQqLJf
oUbXLpNu857F2Yo1QG0zZRPl59IQVaz8QvGpFLo0F9YKzniOA1F0OBNznkpqKDspiEiyj21SQ9Yc
mUmXaFF9wIJgUZQmthiW5oSYOlN+kxmYtyqK4RO98Q5FtYpVQSRAGlYzdZ7U8b9rh9m4vnfuwQwp
x2arcG+3shBL3HJtBKBZNbLo3IAl7/wZJSBU49Mzg3zH//Z4KVnqLD1cN2I/aUHaTB5rOKZFTc4k
6wzuse/zU+kJomKdslzNXmxf3bD+eWY+yGS7DtfcajHVsF1f2jA51lgsG0qlj3YIoCDZQO8rmVg0
ItuagFr748tixP8pFb6sbzI/lL8075LjonBLfs0Exu0EIKdxCH63sjSmJHsTNa5XTxsm27VeCK91
KxSd/vmNxVjZ9gSZT3HlZeqbWMHZPGf6ISKpAZOTMPA5LD9+jSclxNazE+mTCe/iyiJdvSAd2AmW
ujAhnfEldITruPMHyH1WmesEpD/B44Mae4KN3ti/iPZ85D7A0494oheUQ+ZXZhn0Jw0N+LdDhGe4
io5M3h3JBStNf2D1XI1xWWC4WMov/zZwjjsgJi33GsBH0Bq+6YhLYtTeNXsbs290CsmLDi8Kl4Wx
nxNvNwvPs0KqGRvNN/YGXza5T7XpH/SAwgJVKMuPuw0y1/4hU/X8qxxB6IxEh7tq8qv9uw6OAjQY
MIeddIQyirdo/dL0X5l6J8Xj/dVqA6OyPWKNp5qDhKI3PYr1QtM5oeHAUkGssaawZ5h9kRtydUJo
raDx060CcqtlfCwRHACX2IwbMeVRS48Rd99OWrqZa5ZjicjQ8JeJ2OKRrligyCbs6s5kQn2l2YvZ
1o9sqfTPhuX/z6hTJRxZ1FRnuhl833An4RsrG9vtCVHF+1fbRXjvyMtoe27s/9i0m3sYxit9SgWa
2gUTGx4zZTL7QAZlfFjNl/+AbUg/jrIBWpVZ3pFqYM3+O1Vlfz16ii/tUHd/D3MjZd3tGmc1MWxQ
psn0tFucgqWaVTRP8/GtisbcYSa+QwX9YQApSOAplLuTKHs8GaMzT+m0PWY3v2L4WRmsWV7FKXKP
f2+fRvhKFt2iACkuHskmElO/6vyeazuOEZCLaCuQKz9xqbJt5AQRSm7YMtuVen5mCzZrr1PI3if6
m9FkcQtqFnAAaV8Vu57LslPhhhU6c02QmSvUwPfxW+dsl1kkkIYddevMUdJrMimfyPjrvlLxpGwz
7K+5zlKtgKfd7dtSDWFBB+g2LtX4y2UpAyrGiAdDAb0EjjatDFMg/hkbIZthjvaq8nj3AXDaeHDZ
3GR6+LCKrvG6CRzVmNpGJ4U05YvCbiNruy1EwfqAbsKy3XfElIgqKHWW809dvHoO1unB93TCvOuM
j5LZej8QJUn6OejezheQt1t42UsYA8nW1WrVT4V8NUoDMw9m1eziDVKjffIrMpF9r3Ptir40lsOm
jm4VqZRGfZ2owtm/Sg+RwkgJ7fKkaG26D8Uw4+pttjDjVmadV65MTQLUQmYgr4ohJE7VhH8TSFDn
RSR/Lo8JFHBopsC2Cm97W4KulFi/jYxEPauEGptZ+QNdpOndhDvVbER7P17xJId+TgfYuTPNjmRk
19u1hHnDcWNjqertVyCP5owEHBBaXzuQEc/XnFXYfk9b5uqH/ZrEl88MWLbAbkfdQEc6YLv+Mnu8
lL1/UzEs+s1ly8TWFZN/BFjcUJ4XyyReA10XmhqVf21KaXwHpzdoNdc6jCuLk9wU7o3dtc1wdsUL
ACl6hoEwKt59iRWobGy9E4gKRUicLJOIPUCosAe1IBvKWSwNRafLuy4qwplxGHgBIuYsrm4kTmFc
vC0WbWIRcCsra4xTdVZWQIRBhSKTOfjnqSx2F0KXlTa2xOQwpyD2C4lRZ0C5Q76O45Gt0oNcf+C5
uYoMub0TkOWNuR2DJcNSXePsVcWWdX8nNZg7YlLRYK8r4uHfcRomT5x+Onz+llRPKy68UPIdrMsq
XKxKxo1LKFXY503gVdbhkyfcxY6FHqPnhtS8uGVXisfp5C4ussH5aRPqv8DPBD8JMPWRI3JeR7YA
eCMH898n7N/kb5Ue/Npv6+Zlq2VAy8lAuFsSoSdBHtBcz1ETy+fKknvNuwbtYHyMGhbuscP7H8mV
M/yrtySZGyHnOLpq3oNObfrQg3OP6NlFEhfAoFkBI4aUmhLRRg31N4rLxKpqgS63RraSWrhFnFT6
3K3ZtU8kAev5MF7761TICCZNlTmxO1gWoaczCRijzy+3WvhGuTSh5qmNoddPWGpBD2dBWofNNZvg
nRP8l5tHvIxSQeBJWrB3PqgSL/gm7P4Yo9sEdfQYhaBgn8EZxe7Bw1Tlx1n8ZKX+HzWthizncIjg
SBqrLi0fyI251ytEOG8kJvrOZYBILyK7HUpgE6w/SIjjAQx9dsZwybDm1QkIpcZFTeG6f/uBnnww
3laSW/pVvWjJsQQF1j3/lpORAP00d/xBz85IgM576GPg4oMXGKUJ3165bPKFNW1xqJHHIxOB4p/h
a1Q6FTTVD3SUOigRZmmK6rI+knxnnOz86ekrMjYgC4q5y1zeq52DCUIadPctW+jALO3gAhXFQmrj
EmP9WDVMust8r+fcC+vl5g8Mh/YJE6R45krRTAxFRK6g6c10I/hTgaq4v4aOnKNW+PsoQ2XEfaoI
zay/gM3fXtWrA8HJi0MMqQiD/SrxTkrtEqaEg+vJK5lkQsojO0x5Hclw7wFcgKVwiZ2z22MzvxZv
fA7s4tTzLeDwv4+dWn1Uaaeqzs3Fyveuz/kd/EWrWG9OGtQtz40uGjwxNqYDd5AgLK/lzLLHCaKQ
gGEc6qpxYB1o11ZZzK0Mw4uLaZzeere+E7ruIXaBgo/Wv6cAN5vMSGjTFX18UwDS8vagHojOMsgu
a3qKb6lIpOeOmkdxWu5qkzpHs7h+WX6i2ORuS+kpZigCbJZ3+0YbXDWm72tzaSRsARhTwdMKUNrK
N9AP6B7yBYF1aHmIw/6/8X32oaFtD4rlb8GJD6upe7s6211bfu+GhbQ4M5qlhUCWrQUWxKhdLPLL
FeVxwbG1Rqif1nv49H3/w2b7DRlf1wYOgQJwzVqOGWymmtqOmTyMBJMXruVczvcoJVehQBOKmLSI
jp38S9JO7PCaqm/DtjMos4pZYB9p04OM+ZbSy21pS6e/qVcTMB7gz5hl+5RnAUbiQtWq+xyRAjSS
NeP4Hju1fCen/I3olb42umXXnLXT7HgND+wiQwsfCmFyZagYlLQkQK3Lfga1MY0b91Qps9tdcLPl
JmZ3Nl7tn/N28Lt3zSDuI/3z923rK3yris3j/h3UBsSMTr1Vj/gsFz8TehdCJWV6mMhDBD4nmDTb
NqBvgoJRlUkQPkPJNVqiveqwE2WLaoZn5WV3wWaOXmNpjKXZCrR5C68Fo8O/437fU98ZAt0zVaCa
LuR4U6q5XnHTEPyxe56B10iB4csUUyKEFEX4GgNq8iZdtcLCG0ScSFZ9/1M3VdH1AwoiC46vWJBL
mhJSdWAgUsRcQ61i4OY1CDER425DatYMYhBEtr7kLYAxcpUovd+XEY5JwY+rhu3fD1BcsdIy85Kd
mM+h1gcp/OD9Q3Z1i6YeWHPw2j/Y1aff/4Y5VEI8SdGOm+px1wY7LqOXE5Y++FdlA5V7LE1bV6tM
JLgGmfS1VWeHtdXQv4EfLuZ2Iz2eQmWUhp125wyGzPP72oxdbkZkJI0yiJp5yOM5rImH0L/Olo3u
xJYKPHjbSptrKfcKIHgNWIQD/PSuU3ZRoHFXvmcl+elgs4ZCUGWD6Ty5JJYq9r/OkT9Z/S6yEjRB
46zbRKNWP5cTgIoRs/NlaHxq48ZbF1karYXWCiGkyYRC+T6sxleKFxcYIAoGVCeE/lDdUCG/mj+B
WO7BRHE1mWs+FnWL9E25GL1N/tP58q6a8YaQJ9RcBc3uR4U7YEXsmqr1mTvWO3h5RIAP4M25zPbc
gECSxQtBOo80frN3Z4jU4P8jKKXvcWqXId4bMGyIIVhdEp2C9N3QTivOv0RVF2Q6NJ5r9KQZdHAS
JNFWGhvvdKu41N+ZbyURa/Y8D48PeAHD2xOW5VSoPbdER675e0xVG8jcpOI4LnT2AtyUtzqGjeQF
F3+u6XlMtFZR2R140Y+X9T+9A/TrGPrctEP/cTQBn37P2uUCOQ+eD/Ier9JqDkc3+WDQB9UlMiGH
smDiwYFUVWmVuEkzQ5QY6v5AGd/ijhLkdjmB1RBBdUjduMGenSutmcq5RaAt8gIUbvMco5PojoZt
Kw519SCnWugxsxvySHF346J05NpX5+5oPDkFoa/PBIkjahsRCNOkQaiYELmcV7eTMbZdFlUGiJvK
XiyFnEnQW7zGkM6TrvYXsbgymFE98j1FXxKaQf6jokaSqSG5onGeNpEKNbZiW7xDtqu59uJl6tck
25PDwh4QoYccah+TAfOyAkN1jMCsBrC+qjZkLE7qfhH03kGB65o2rw7szoQZU4SNN9NjASPP3BN2
n9G+BZR60IpajaIp5klqJw77wnw9AYlZ2OGiBTrtVprI85tO8iA5ANdpiO1ioKQ+qCEqfVL5HTXk
hGTljJND7WjL0F4wkfJa1pT8PDm+oTEEjZyjOEOboM6Odk9Qw5CMmkzvDSR7Z/DIhgiOZPux4w1F
RS4YtG0D4MdnVDR0r8MA5bDo8GrRBDCK9ktGudRhaTxQb9IcFiwPuCD7atp5BeIvx/XcYkTAoA9d
qG+KO4AaaCLfj05we3/XenAGyWmivUvPMFiQ/CBcOZyvg6hGVz5F5UGCEhRUvCbdA+vLKxemN4AR
bXLEUatH/8GfZDH0cISHyvjfhE7nmJjVDO456AF1n6+Q+tgz9BRfDww0Bwlaz2srBfWNa87Kw/ic
vPtsgiQEvVEHSVXuDnD6E0kS38gzX3U35kEf1h9cH/PlaMqy9NTvrwZKHnhWR6jZQCxsCJiVf5AA
qzeEmUBJtVzbqhkbyZGBXnp8O+yQQaARp/gSOhfP5s0CtsEVDILZl8yPktzZIlDQ3/nR/Twa9ok7
3V8e3l3h3hSy2RkDpkC2QHZ1NjVztZopvHxjo/DRMum9m79eDMiXGDngG9ANSF7UwLf9uSg3pwQ+
Ved7kGz0B1C62G5cU1IQ7jDUzu5Jt1vgZonEwMgu6EYTp+SC1SohBSpkE8ObIhVVOKDN7N7IxEsf
y72cFM8VamjYmyBBpj0+z9irg/MnKem0VJcSIDv/XnLZPFc0cOiQBv5oR5OBqoF+jo81H9s0FdNt
phx+cbor08RAzq5pAqLOcEqImFCmf18exBy0YhMxXg3dnbTnxZKYVNT9aeM6x02F8E3qE0V057zV
QGV40gwoYVtPCg70ncIMH6RFW/a/ftebuCFY6M3RdPn6g2mwSGJvZwEk/tiO1j3jOrUwCG1KLzpK
vTWu4p36DJg9hoNPsPoIsFrfxnDKBTFmJJ7OGmfK6gd8VPJJhOnpQ5Q3R6qjpiBO+pDRRUK+syYs
pbXAktP1tlzqlHDrX0QyGUPhB0GjmOAlxVYc3UG17itXSG63wZg1fyKMlRupJuMJeyVkVA3wFxXf
dJAQcQxbDEJ0YMJtS3uue0VZkd2JkkE0AyyQQFQe6p3XFDi+G0Pe8Y2eNQFOBQQuCbDi1ZxQSduN
V2FllhtECtBXR9LgsxqRwfUgQq/30FJuduIugBaMkH4ojH9AbDKDVCSdjJYZg6H8TsjGdMd8RSJT
EHE3ektHY0tzKJ5S0wYH/iW9M93y6Zdz50Cvtcg5dj9AZszqAmXCU8yMBUHvxPtcf4bU+6Es3Urp
uRjgp8Opi10acGLMoFbc0QByv0xGE+qzK9BsSgJPJJXoyLLfNXx7MrwhjrZ516cf0Wdm0qvnFLiP
l836YH9NVADMet+ymVPFes5s1fWlq+aw1CUEpfqsnyyexEOA/hscJPlsSnb1zAzU9JFI0h4TeubA
uJFJIuuO1NJzd8TpkLbJBW/pUvyr932dLqaexkMJpogXwIwWr/itYo1IQO+aKfbXK/ab1lKcW/Xx
rA8nFruYdej71lw3TMUvvV7U3//Ga2NcwV0YFtnWwstueYM3xzYO1iwV/9756OTdTCfMBmEKaD99
c/vNEjke/hc5U9UT9QVLn3+/Kl6+IY2cVP4HIZhlshp5PTGKVe3dS3wiJe9Fs0Cq3a+7O/jI+35p
zryz+gQDWFH//UPq3VB7OkodDJ/fDP58huaZbDKmhVYcCAT2uHViorFsyovr+fUhILwcPAPPIAxK
TQLmPys78lctYZQ9IQCoQZm7ATCFAmsfK8wx2otXYWY/dV4RFWRCmHwpop7C+s4yy2DYOv5QE3BP
X25YviAQi55YuTyyHuowmoAv77C/V5eikL6csdbgQDYaNxAgi20zELLWnjUAhyrxZvDgKDrbGryD
CUTyLf4kOrZ41Bwj8+fMqveRJEQDxvfbpKCXZw0leBEZz+FXGDmy9Z8McHW2S1eYzHSuRw8XAMkN
OpNr92yrhDa4gri8HcovyWg4aePze6VCuLQ5GmCV0md33NAvq4SScoF8aJI5gKLG7TPX85+SQyma
gILIgo6vAb0OBZCe8OfqyI6Q08ZtYZrd+V9Q9rgYeYk6aj+IRtIrN76WddDTCZURAI6YWAoyBt0Q
SYsKFb7zoaRmEamOxNRooZmwLDbJwxZPy/WaOzjlcNbtcgecvkKwEOdkDfKOHO/v8Aufkafe2srr
n7mSwbYhrOHhrrobzpvYLJJJG230iGGiRalN9DQe43VNN/2fQZZoHYKFGD5zMWEbcVa9QOCFHdLw
kmwYiHq4JJJcTWYtbK82SXUnA27aSSADi+xGGo3KFtloE9qV8r/nb6a44rkpWHna9ZXj8UvVf1yI
cdNP51uAcpX6APoMj8B3pXh4NGhRl9LqBRGUM0kBYCUq94PvgWh081WvD2xinL3CeNWuTJT0mJSD
Yf2/yl5ZdB5ZgI/W2Ky4+3vJ0APh7qiTzsjTRXgvU+Y0zqW590wyqpJhyCp9wNtEi8p0xM3Bi/WM
Eh7zyvhtSBEUbOKkF/GhJbkT4kjScZMcM1O+YFTsq/El4F33XW7MuZQlWnERh9dp80uJImzYs1li
+X1hSKISedwhjsuUldEl7qlVpl840LouLzW/0z8PU2kvVv9jNLtwIDk8KEjvFvXN3sGMpSzQDVOc
/k0VIQnOZA9EF1uLcSawdZKo4yWwngpYoY0D7YNNCUU6pSGK9Tixa368tvbBAXqDCz0BmQB/eSVk
dE1hld1rgFrEX18c8rLgwqbTeL085u6/rYsOrfhy5NYiYs4OmGRDBMI0lAkLwe5mNbw05oZNcszz
AIASxh4dtj+2ZGkrQGss23UGH6T4mhmRKKGgF6mtuw2nHEsudHJYjCVNhbdisznm/kHEpdlW0bcH
3HplTe/YWtH1Vw2vvqxFFLqY5lXX+20prkJ9FpiGE2XfBV6a8lNv6vGzayeVtMRDocHnX2+74sav
QB/XG8yvbUVFVBChegty1+78G0ppAkcgpmTboAHFFUKm4GNgMyZoy0/0AoSvEA+5qBxflu6uuWRY
dImz+mGcyPjsRzU6/GlfMushXOAtTDI+dZa7eM9V7pRaFY9lBtCEOIKq2YethzoTZm1bi6T3PWKa
qQjG84rsev+CP6Lb43xz5keLYbqVGr7tbNbwhyOh20C6KXwvi1L166V9m/m6xY9PlMku1VYBcDP8
PieS4ZFihVUBmD+O2W0+zTmszdO8YQlSl0aM6gjactNPzCzMMx9JJ7RrJ8Ga3K/0tlYxPnIpOdp1
6H/D0qgmaK4NJHgtGFWUuiA9ca/nclivq/k02WGNjy5wIDQWTXlZ94N+bJI+LkvYG4UgX2VhaEg1
Ilc/TqLDxN82G+XV+Vnyft480TTp8DqJ98hxEmFXUC4W2JSGy1ikBXGGS9hLbRzR1ZTn/nMQjwju
rdYOZwjeYP+7zK8Jgtp74YblBxP+QHowOOYxeZZGJ65pqgEJp75CuT83mKvYWFH4gbz1S9JapB4u
NomXZtgFUeKN+KfQvC27SEj3M1Mg1/q4MSqAX7q/aUpSVUr/4t2eN2WzDD+F4HY9FKS2+qQWK6PH
fGLTev5+grxONvS35TwVxf+7/1Dg+oIUJ0g5C2+lGbWV7FVG/U71Eh7F2RIl8+NCe27R/kKckJMj
w286zIcWX7tB3z6h/NXfxr4jL9pvTlcFpSqiTVbrR7nZ5A4oulrquK5ScjvC3ZYQF50/GB/XA/g9
8SicKQqjjKTQeI9h3TOWY9ZaxMg5KZxUR5CPMqCaO537qEuCslr4XsZGoBGuyWAMIfDJhuKL6N1b
N/sdLj40ybDVOW5o4OYoFKAU2foQXq4X1KedbxHiRgneeFNZbZsur2goy9B20f5FPMBdnR9+3SN9
XhTO7Ft0VNpLi5oq6Fw2vC39IlHDOSXyX3jC8wLV+ZWikQ+s4GagUtSTPgzC6SQNzNuhqbkQQWK4
mtYrrsrJoi1pd0fAaI/zM9lustN18ZrbXllgMhMUOuK3Bm+5uA6AwP9ROtCkchm+nfB7vjeqbNyp
PJdIF0zmesEwJvr3I78T0sYs/ynqrvNm3Zpd1gEwwxikW84AEcZQWS4oiZJBKqkJkVqiYnOZNP2q
1OT75GO7tlw11kbMf4aYIh6pGq8tXGPugbaO2PMRiXxiTd79atM7VuoykzTISjDDArXX0UlkeUWR
woG/EMAMz5jidlXvEygxMYiOci6Ldcb56oICkRDSoHLpyW/cBr3c73dCAA/xbijOnciRx0NNuGkV
xa7AbKeJChwmmQCiH2bleCLS8L0W0crSt345ivUHCVq5S0lAArhiz4eBoX8P/HjlM5g354xQAyhZ
/GUkgqESJqJhD8V+6BVMXqzvG8LvqmESzVFy/Kbcs8ZSLNBxtvyjkfF3QaY8pPqEuYgAoEvMt2Zb
6UBbp7XBaZ46cv8izNEkxy90Snp9aeHXU+7mlCPWec0tPxMXVvdB+diKy7xvPLdmCPn/eG+rdlEq
y6/Xd3VFamSzh+EJ2QUfyIUL5UwtAyf6FLCvOZ00c/qzYU6ocgysL/uG5pSBFLCtoSM1ev6CSrfC
KQDVGT6sZP1Ft/HanG2TzCFaB64Z7TZdyc6NPsUBkegTbnoRrqtOb5c05iGk+ObZkgHWCNDigW5C
EJ05gYoINekotGeV4JQb420uvwuRs8FPwXnUFD8vZndfq/6zsBQ57SLN+UWfC2/yj4mRk/rn3VHD
TWPKSshk8qiBpYIkbf2bt0Jk7BptyuxsW0F7jfSm53iqRYt+ILnK4m/Kx0Oq1Z69X4YCTumkJJR5
xbgHzaVZb2tfhy3dizhw/3GwyQHtm2lFtJkbAXOkkzj9yAh5nuk93FxVVaGZTJ8V4fO8IYRY9Lrg
PilDqPnav5xyHQi6JypiEC3r+gMd0unvaPTlBHHhvdZIf4pro9vnDi4XfzRQ19oHUE/4Nie2Va0K
9bOnoAY9wlqAN4f114EyUIv3qGF/DcOQwncI0s3dGeBxTOp3AnIP+QvQ/mQkT9jFdbKjAYiCNAmG
e4R1yX70tLFDP7zh2wtev+/oQz3dplRxp9hIPI+BvSYdLFP3iFmVNxGsvE1vMT4IlntMU8FdNT9l
zVTPacJbYKLAhkoBSxG4yMHy1FHQtZ/mqcKdnI+XyP1/5c4Aopko78/Nr1U2DcWIUjvyKe2W134B
vPApFEa++D1IbwpsN4rmquBF+H6bGKsBjZdlEZ7EyBp3NkDt4UU4z9zBERQB9Kbd0zMpqQ75iVku
4rVfoOIx20fbrC9IWIZaWBPCLLpIxc/gjRS+f2HDg6f1Igx8C79oP+T6pw2k9VQGwaOE0r+f+SnE
PhWeDgrvUSXlaXoqS3ZRd/y1K3J8CvHnKnnFMX9mzNJxY1aTXX/s1fy7DJdsCsHsWya/leVG2sxD
3VoaHH7nLATdHBe55/Dx3Ya7VQ/TM3J2LzUnoaPfmjpoCupa8Xt+0rUHTuYBusWu05w3JZ5kKt6G
gvcs2voVyihICbLdr90tUIn3fdhHzqXfoSYvEdZ0ujG+QhPxmL71bT3jq6jGoYVS1hNEdAl7y48E
3JNnbDaFlPrZnOCE3wIV+Jak7rpqXwU9/KnrP0S5OYMyKvHyaQNdq2tXhsmIJVnAC27iRjKZydsk
T/bF9kDCpUl/80ouHIXyRIP5QisOgjY6U8y+LTxEhZCb99qOK6vIfq9y3Nl8Vvb+5Bvx3VnH5pqi
rNvjye5oR7atwyxuwhNpoHpdHgU1cy2xSypO+raGMeVgRSJ6eAwOhXoIh0OoYk0YwHQ7MDg14bVh
xXC026kpyHHkZF5XE/mYTPsrZ4fr3Hta2kt5a2bgDwJy+d5dUfxEkESL6FGDpG2g/O7JdtXHAbcq
bo1ZiFaB2ddyTmaFIBbGp2tkVHDvMb9joiFq1wzas+X2BsY5KudG6i0WFvYxsM4WEuaTAhTHILa7
CFXmcBo3cQSpqOx+F6SUorBpMaYUxvcx4KZnhZ0xmLpmeCYZauvbfg0a13c/Z2h5iXQ862zUXb7c
SRyJgnBbZMXvRiVAggkd3eoOJlyw24hWhwq1VpJcUzZ42dvVwUFZyhvCGCvr/LPtqykYY7Rw9y4v
gKnG9oLMaiaBceBXVT+QsdvGCIz4lAW2GGPkoYnWZN1HnI2l+EY42hCCD/xiK3QoRaeuk6v8amT5
374G6o1mndsezaqltfBH6ScdwwZoakCywIlrtVLK6sYkn5HDh+lmC1DOuy74I0zcbfjLtWtyDELt
QAazG1xxwvNdaBdgFaXajP27nhPnzrETzNW9WA6AwFICI+zfOASkJFlpLIVyfZDzCQoN8d+5K+Xp
dzSwYo9WFTb6/nxM/1crH939sSLySKQMvh2nlFx9jYTSq/VOsEnIojpIDbHcc0JXSqYGmtS9bCqP
NTHfhiBwcPCOngZGMI4Dl2mx6ZA9yrnVaaKb/I1xtflPpcKypC56GlpL2bXz98FWbKjWis924i7g
rIqckuNlDY1ZVCNAZHSFx7e4/V4e9FDZrUvTXhzCk5/BAwECz/iSdjyc/3RLCKE1kwSwFeUJECEW
UOStum+lz4lNuvrFYZz8rh15KSvvzatxgj5MaB6YndtbNGr55crr0hxAVweV8bFm3VXTcDMPGCeU
9qRx36RtWrkEzvcEU3JhNMJ1vylgdvYgFpkbMAeBfcNyJyVbgTYAi4xZfeeN0Eb3XlCO/s76ljpI
CfBiocEY5w5boyrnzecae0yUKbFOOsvOUl0dpoHEDPMjG5fKyG2MCGwz2N92xRCSHyuwKncFGTwt
WYmRl83Noy3U3YRUR1G6jlCPQiDP+9V0LnflxfC4QiOEUTx4GIv1stRdNEPh1ZuZJ60hRlkOFu6u
oJvGIZM5ygwPCXJyx5RYKOP87JEp/zsNIYI3s0Q2nj4MzDBANmWzPh3r19ktUq4HFyLBalX5RMND
8/zpeqhHGsODO3huZLFTDBKkYRFy4R1TZp28poURb3OZKyHpjMKTYqziPVWdmmnben4Yefv5+uEi
9ZPlw7GbOBonNYcES2xO9YTfYD0vDdnQhSwFdmzuY5affNm+BAe9ZCB+H3ZsuUysX+12gN5wIP5t
GHj1gDOjeIvoEntRqBydPSfnfa+1+9yhaenlms8PDgS+oQ+H3aqnowQYCs9QMmM/WhT3nR5V9hLq
cy9jEpIlciL15ADKiqPPuSqp4FSf2E3NZLVhogExOSMRw5ZBUeSzyw9Lf72E9lfS+aMKQNdBE/9X
9ws+itV9i0fVmER0f+znaw4F1/O/im8r7W59+qAh9NaCSR/lVXhtG/9yixT4+1eROM0Zm4qLnYpS
xVhxd99vbe560wZp4PWIhRrMU4HoU8FtXQsEA1f0F8TNmj0t1r9L0pt90kLycAMP1OFCp9xqTQ0v
X0+ctB+ZjXaOsLo7bUSmdh395YSVRL/ofAJ9vKlA7Gq1nBya3HZRpu3QphXBzrrZfUYbD6YUl8xQ
fypZdq9QlIHX6n6tOMEkiY4nEsRqgAdvHv7JYG4kHMNA876BffJ8aAzDnJ2ZdmAY2BxzcJ1cgufL
Mh1HTvrHZ3PG259hmWpg6+5yZ/fXq88Dl6T5AOVKtlBkNaANTZU/jZDkqLm9M832cz+x09+5cTRb
wVk9AQAEUxTiJM7lv0YUOndiPWaX0J8VrW36Hak3UK6dgWfeSpx2UrGugANeCgY62JvcqS4jBZRJ
sPRmBr+4VVujgPHS7nroLO+Hn9AEtzJBuJ79nKbxkERt+sQjT5fWU95/LZH+FU9S1b6bk+rBgPvs
tzpErIXC2XxschBVR6UfO8by7TUuXW5hMbG32+ECbXRM1mCAeGUuxyxjOX8NzIMgTF5r0PLxFu3y
EtgUjy/8ZRFSmy3MR7bOYv/q8fB4osH+XVW5ScBcObPIY+jMbsxEbmZX4tDE/jBUkJaMy/0DUXeA
XVRyMzfE6SUSzo1FmD2/6wR8dfaAn+YA94ha/clrsEU+ADMBg8dG2qCFe/TbkqzZZVpb4YBijBMd
r9Rxt+9vSCocPF6tjNEhfcPNFK09TCb6hXi82zhAdtlKlNJ6jCmIx0Y7J9wagJ3SLU4No0j6ylCk
2STBzTmdR1zBNk2WY77/GoOCHUsxZGscJTDvkValHgGqFhVjyrSFjwlW8sAWDXrHBwkMpsVqcH93
Hfeedmn8mFAmVOsgSZ50n9kXIKJ40nVu/v5bcLm3ByXvLjwiwzZ+vnNEwqk5dRwJlqzmqkwkJNsM
sxvFfTLBDM/qLZx29HRu+GvAatvOjnxne30pIo65k/nYzHiaUrH+VwtSsaKZX+rBhSEG4J29Q8hv
098YmLYBObNzToCfZvt+cEzzx8MvMJL6K1ZbPqYSJoFGs7yYAhgm43aUROG2+f0JC5ERpQmuhD2U
3xi+zIik7FjrUilph7R8hVBPjbf1Ub9WcZxPyjzmsdZ6J1xvmF+cyO1WgjUvg4koGfITRyfsYLcV
71sEwkRdPZSsFFA8N2fFlf0jdNqnzQP5E0HBQ4HTJ9q3XMTnUdaNl6twxVeRTvcV5hIBFCMjeqWp
LiKrpuDfHXK0Ojzj3gyld9U0ghNjwg2UPA9Yc2VnnvWK0ngb/ykXwTtil3gIuDUlyd2DMXArJe90
G8tnin1CQhaPYoNxZRXZOW1eXoYxd6MVZTQIvAZys8Br7HOKOElFQFTUpYsc7A3M6rzKS0GZ5Zyb
cconcVqXhz4fRLiqHf5VG1f6SBVxYu27uZaaXs66tLI1ixUjOpt7YAbDFT4l2V9FC/HjLFQ4XmQN
9GgC5h3o2b7ysQeguNVfvzTEp/KU2HpTWGeL+0EVcpdkfBgj5gVOhBLdgcxJ/oid/R6dG+k0f38z
vNvW+yrRzxiXoz6u4G02Gmt23k6K+vu0cH8fh3J4AcZd7/EcHqPXEmd56ukvXdXFM4RvWSa6xGpG
YUiBLEJG0d4AUaComTD0abVDkW2jHLCwOlpJGWS9YKLZqOSB+zJPKLsoX2XGrfu01iBd5w4JSW2o
3lnSqnDwE4nagHdu3M60H9DBkM5k4i0tlAVsApQGAjyAoPGkJnJBxayoP7E4lGHwo/KU5/TncwRI
LYiCtZcx9ChnHTu+53UP4iT/Ce7pG3aq+208SgkfJIfVRVCaQHHJ3fdgYyVw6bbcLz6LG8KFIX+M
PVnvonPwmcNWr9patVwXqCZKQsnmNfGqkq5kE/6r4LXtlfGcV/lRcYqXVYCoOxviv/0N5ADS5UiJ
5b2hr8F3EQlw5mbkjGnUPyF1+XDF8JFckGNIT3sh1g7/QMBHK/IUpd+2hBovPFoNFG9ZBACyq/LW
i4iUwyv3O8fUmIpY99lGi+jiQXOsl6idXnTpUB8zcXnMrbAygSnG6sNplp6Dw8aZnNhAnMrla02t
Bg3WX8ooqTotmMx/MtvsX3VP5OBowTqk7d8eORobBNEKornluroaZGr3optD3YBR0bLO8EkRsbLp
saiHtSJkJSIwQHNcKkGVzXAkiOUEhagCzPGD92wc1G13B9+iSU0gVgEQCqzFIANMFRZrbQWN/cf2
7XoJvSEVWUWS8BIXZ908aJaqEAsdz7ua8eN3Tpi3EyrCpwQR18Cz/cB4FuEbxt+AHL771cJ+30GE
BLziaftxYZW4E6F9whzjmzKAu1VN7DZ01AsFu4njYphaO/CmhynC2qnRC4F6EOAxJBMgucxgEGFV
ePmxZMBxj9koRrchvxqPp3fL7ak2LX+r8XlAVEZvOT5Q2AynHxK0cKYOFUao0sdde7Kfy9KirKbW
0LW6pHwaIn4HJOe/GT4O+izPLVuMsPOdeY1W401KHMEpwbQwdkJyzhkU7THi13jMtIeo7IU8JBZB
Mc0cDm20PGgPvBoe/vX4laRrSEuP+jmuTmlQOs9qAG/paJUkY+Nvou1Uxe+rZxDISpDty2g2dZ1H
7G01Am8hxIGKfmZXT6YXhw2P17pJLWsVSyeQv1vPFxA16KUAG4Zmr4xxOErTwm+pQnvLM244MVS/
FlNFdxZiFNZV6QkF2PoVLXtfcKRBj8Uzl2Y0+XoRdAb28jMsdgmjC1vsWobTS2MNabaW7qKb0Fr1
V7JTnX/15LlGnw+edjcUcsdc4hvfwGwkJOZQ9rXVVDC886WuOTJIthJ73p4mWUKXZLkUxice2r7i
iMIxAsMhWhTa1yJUP25gj39n627dsEDqxeVxBRPQdzfuOZ/7qpcbzknQzJ6JQYQq8yhmkaVU4N3d
gS8+knPHMKCidEVBOt3QG+w4m3L6ZGhsen1u9LHoFyz0EP6AYbnueTEiJqRJ4+iJi2+3qjGsqUh6
N3EcRYpA8jy2j6fJgnjGm4LuyVTllmuQtdi2kvEV6/k5AgtbFxIWxDudLYJXHqoraGA4EcODq38x
sUtRJ/NqstLvxrs+6K8NfEwqV16ZNqpEamxatGjm8Fg/Nel2hZywaUsV6OSFJ6GIztNkAixzTggx
x+KL9yFVqd89s8ZIO/O4zsSWY8yznCa0ur/978jldQmGuaKEXkiTrvhEnDQFXrjmnD5qaY/Jfc0r
OrVjqK7JmdN6FA5IE14m4Oh30x+6l8hliblYLgyQhLSc8PDftMI16bkf1+PDNCUhsouVIKYCZoxE
1zR5Hh4okVSt/YkZPtdYqsAK+ywKEhVroW0RSp6CI/cjSJPi30SsWcHy5/tycJFDJlNvZP2lT2j1
y3NdsqCLjA+QaYpOqQwgLAKxyEEqhE6pe/6JxWmvGBKGoPGHoAOyPmo5SEdC5wS6XaKVE9FGpSUx
4C9GJXImlYCHD45aAKR0KRKgDer7mQeHYLjgRK3cfrVNo0CtHT10Ox1sDVpuG65678+EYnn5rtRS
2T0gk1DrSVfrfBuhllHaFcgC1c6k+8Bd7nUjOeiRtr2j8qN3CYgqHymPfo7tO71Wcd6bKs6TU209
MmU37mHLyN5bNlp259dc8EST0ih/CEFrV8q0rotvAbmcWOID79UX7ghOGmaS3OuG4QXJbU9aHei4
RuJIh5EkwQJ1e+0pYRYBqbkFp7WIu0v2jp1jQdGOoN5N6ZY90MsFKVAYgzk5Msh1nb96ECUPzpfu
Q4qVd19HyYLdrkjFuG0Zr2Nw0twav+mi0+mcVA5KrHl3O21eTGhvnqSOhfSrGgav65hqezjnoO/y
5PZP1fHz439UNQIOfZyO0lRs3xrH4eIkhRigisuPBQrEJiPZx+BZCAJKqVliPMWk3U6F7fWT7Zno
2RYFqRfdvi/peXtkigV+P2Dh0srUu5/vDEtGRCus1l6iKdBHsMYPMEstRYwTlO9+Wef/3ayELVFA
r8c4BDGJjo+Bp3sIO0bxKjt5hwUboFTAvgD+eU0xMsNSO9+mN6M2RmBjo1FGjUQIuJdMPXuptT9E
XyB4hdl9P/HKRwMGuKCVvY6xxXk4PYR+S7XNj/VmFZPYxYQyJh+yej1vxobszTA053Yka7h/L5it
OSACk6LOCRGjoFsJcc9s65dxczG/8JPf2AyZo1Im85NfhMfRdgBM4zLIz0hpyzPv4tYiCdle/oul
LXvbEpw1GXjD8DABJ69+gIq1JzIfH4XZbpxqFwJifA4yT3ClWI+8XwSSAjYCBWx5dzR7qnWwYq3H
v8pulSkiqje/yCUrQRB9Gi9+Xo6ccfVQvREYQYZhOgleJl+2gP7ys2NIkTnsfsoEqE4qTpQh+Zk3
L7c2gYVOMFIfpAeqlHk436BhUoMB+MDj7CFaoZmxUe4fTVzJ39P5Om4gSxJjUBveWgBqh2RjZ5X+
mMB131yZZVSoj5bkqKv9bLfJJXg7zik9TP2Lpn3sXz+r/mN/qcrJNsSnjXYucsBGghD6rG9k2hmj
G+fothWy1x1hgL9H7NgHuRJJ1Jm+k52eNWTrIqAUxKI2v9vGbXtxYCKukbKLYsVJdbK8dSXw5Buy
UTEXuAp0zhYXKBvpAwS9UiiPnhAih0+BOma8ZtKFocsRAqfi1OtNoxvoAuWSDA9MbRhERUmvuf2X
qIjNN7sgL4y9skdFXCy8GPxUnBXPH46casnyUf4VaLmgEGbkNtorFjJxpnGVqtancc38cyFLRc26
QVZBfmgw3FX6K0aLwIBgljyIi6cNnOs82cKhWtu8azrFGYVXZjRva4M46Bsy63DHgtPL4hilBYu2
eOXxpA22TH/r+DJ9JPfZTEAWRRYSuLirkjCpof8n+TDSnpxsRp9aSlHTv6FxYy7bMzqVkefSYQyH
UiSSwFLYmiZG3LE5PFi0vzTxqNP96+IEik9L36I1Wulo4Pl6eD/u+p4OHhBVca3edTuoL1zBQa+J
Q7D7En7we4JIbODCs3L+lasWs79d8skuKAQm3yqrw+npHq7tXNeMEdt4kVrJ8KC+618l1JEIqHF3
LiCPMhk3aQ6rNUSArbXOmy/toC0i9LBemKKEz4aD5Be5g8erkopQSRRGGeRG9y85rEy6yC0Rdea4
0gzV/VT+PYhh2I7yE0edlw+NbbjFdY+7MC37SJ6ec9wLiiZiyTuzFPlhGK/5VdA1wR7oRGiGVfA7
5jSD0H5UGPz+1jrJWowAk6Mc+ykqMlEAp9Np7ag1TnLi7TI6q63w7zHRPXrcSzSMcTrgtVeLiwDS
xbBOKDEfvILdIUEVnd54NoY8H4SAOmnuiRfLpZ860VemxTPDfYsanm0Hj2er8tfpZlnE7c2gpLdv
Q5w0ileG0BGkjc1Kf6lW60sGO8H7OulmWuEBWJeJ/FdXt/N1hF58V5emzgQslDiJJo6DecMUZ5kd
5ZAcPBKZmvw2nVN/pXG9+GrReVwkosXuTqZnB2oto1ZQy/0EGC4MEY/LQG9x++E6rjzAcHFIlhG6
cGUg6mxrkPxgHsAsi+sjzNsWuVdCbeGcvrasir8Pv+5GzIDg+0Xl/XRx7GmiwXlapyqGdNAYO5hu
2khsHX7k8cQTDjiMSB1Bz/SNnSt8krx8wyWV4ozrR5MeHTVRiEPQnDurJhqQV3gNW0NrlkPp0V0S
xEaHBYn48y9+ZCjAQGlcPGMLOFhpmzDoePb26jqSIifSHNWGAf0YMiw9MsLcaZRgYcKcjraBpyqd
uHRBIkgRO/28x6Djck30oQCI1/oihqkvAEW9Z8J2Z0Zn7ZQaU70FS57lO1joxpYwaRo4E/D5Hcf1
2IjvL0VdTg0xeknDDlYnyyy4YSqVVw8ECwtNS6AfAoOKC2rFrzIp7dEFp7lM92nbNGlprZl6UTUY
5AjpVmh9v1if4lvHv8ePImi3+cyBYL71y+EQvJxqdR4OiPiJRsJHB/1nXVNTetbrKOUIjOSVS370
wGVXigguhhRwKnZFPye61Hvqv9ysubquJ34Hp4/exXrCXR+56Oc/O6ceFgg+trV5PTwHiC6qMHI3
O5S7GqA4XuD6w4Ojptw+QfODWv0bEFi44z/CqNMw8FbPeV9EYJs2yfD7HZLQ7D+p1u9u5xi1OuV6
zm6UrHG6TpnLgpiS2fLeWYlqk4q39dljsQQvWti4aL4DJde2+YpTSDGGt7EFSoqxbmTSWFW9zFKP
V1ryKAxc46LtntKwcLeiYReVpMHMDVolYeVNosVAgtQqdmW4f9SWTtAT/niBR3q+jpJP9c2nJiIh
t/oMe7JSvbIODvpPTuWP3a6uFkBnxpN44T0ewL10tZaxEqAiejcBx1QTW1Tl5P0UKgTUi4dyEb7p
C9lrAClpPUuiTR9BApebXlLqfnnw7eJTlWW8F4kfOBotdE1o3JYUGToVzwvLnuCQFYCcSdM5Omoz
4A0nOMgAjgT3Wr/pJVtdyhF9sWcEaxSLmO+07/R7umAh8FaGRHMOSZvfMLZIrCAYjSLnaQ14InMh
eCSpbgN9CuT1UKMQw8PCKDiq/WBnS+//fp4Y1/JSvfbAwfIbKmSYXKRFMJsnTD4NZ3jVJAWzArYw
axIGbGe5RQgDLQHVTIt9C16ZEs2LRpt6N7xzTPgMdtz5rvYc8FIP6MR/ITBnx6m4oTHgNynGbXLn
iBuw5DDsFkZ+Vj3D5D7QvZAiusSIxXoIcsErwWmlOqJd98+5Pop1cPWNuW4qGY6iy1M5CLPNIeW9
ERbmck7sCkxPx3XNzl5q7bM4cfovt3ze4wzgCX6nJ44CrrLFdaRZSk9SAGQbeRtdg1BryAmN8PPM
4G77ipxLXDIhLiGuFiX2/Y/ISwVyGXBOuFOuPHHzEozM4CM6SKQzIyWS9b7p6L5izq6E7t/fJf/y
cpesGToi3jQf08V/Co0Bzz9im2JewN3ZM97NaLVonKqdje/QMLjqTJXns68BqT5R+dPJ0flzdVMb
/m9xdPFAohZNX8Ga6vtgzesYDvoL01Z98Onoa+fcPmopOCFWvbWZEj25B7rVSTn7tuLwQeZ0aCNV
OhLxZRVB/ijOipwDu2mYODm8EWKQUQc0QbX96a1LP3gvg368vQE6aT9a9krWU0W1LTAZ932cuv7y
wc79xFPKKoGp0X8xannsP3p2DmYuggwNa0O9uJQs3nj4m7kduyJ/GnKTT+2CQv10ptMw5r+IqU4f
XHcyvo/sQwdTy5JGWLChCHQ8/2SdbPMHEUsA0Rcj8MguaAqz/6UnMvqWPbGaxQViOOA5K0WXU2Z4
mB0w3YkHTwOhSEtCR1HKl/ObF02CKawA8M22vVc+8zo9vP8Jd7BsXrLdmJNL5S8YTuOi9MvBaszQ
V4a2fTA+DZxuZM95Brh+5jKebZDBlycb5WxBpyKGLTJHkTx0ZvwuObgZ4lNwISncYXtTmCgk/UDG
CfZ7lVwcUVtfBj6g6Gi8dK2Gx9LDwSgKRF1tuM/g7x3gBJz7ZZBmrKVry5dPvg1pQPsg01gOs2h7
jhHG/ppApwD7dIv8LSHQp6ttyT+doIgSmPprb0/lZ8ZCAb7wOmaRyO1YbuCyBqNfr0VvZmqSzDCc
u4Q2rcyLRgMofD3aus6QQRIB39KIcYy1DLUndWpK7anpQd227fa2+27jgkBYKoAWup0WuuEPfaSF
2B0XzAiLgFkAtPPr3RZmLZnt6BsJecA/MDgIMcTxFt7PCd9IPW492xze3nCkDPPMp/fm6HazNTRo
s5z2OaFHAENyDDeDIYFGnzXpHIiJ9EqIBjw0OyeZ4aiZ7rJ7zovSbcAnpkuzncUVLxL4DCKqSGTN
ny8VHJhlFmjftr1z3emBAjDYEysRmG0Z1W+iPzrXw1QfSKpdHL1wDmTKYaqr3FciRv69sbSWVPGS
CGOn865+IBEZzJ+iVMojoQAE87Ama1Jx6RIMez/ChIkpgoRoKiJ9Qa4AmtiLB950/YIgE8S+kwmQ
5o0ismiK27kJEHGJj67Wnt9Pqn74eiJsLu1gQN/xI83KhTlWBPheg4wOXNzXj5xBGX2UbBXo+XHH
lGhcCCHnvgLJZ+vLNoObq1QXk1NN/sJ1+KIBU67HVlmvWCYtXitvsgcYwDS2lZfDLJcS8+NuJlDN
oNBJzB2zJqVSPFhn3IRwzG8rzg2H3iNuQRzHHacz++8YXTiPnCfzfl++58Su5Yzr2A4jmfaLPWCs
Gg/XYOOaKCd1jOMUff9fHwvvClnljF/XIlF58MZUugVrv5RmXiKjYIejD3+Rp6lWMkRev5JSrC3m
my+oD52Y6cUTyCShkAmMNx6QAJZq5//sZ8gZBSlRpa9eCSVbwdyyunfXdMa2Q3+jHClyN9rouam7
YZSzeNBxSB5h0xmaCPYkhe21Bt+wqzuXrkQGvYipRry/OxPXQGu/bnBzCIO67jA55VPJw6x4ZKEB
p27r7GxJ2rliVHbjJPoa+d9Sv63a6J5G4p2gPuWUPkkHGewhqjye3qpAInOIaDF0S7DT2f9IQDG/
qMcffe4WL9AjIqxjVWUmzA3QS7Tn/v5V9Uj1C7FuV/1UVlv4gknZzufBtM1k2LdQ5U6wkU7ZEs1X
pA4F5mV/+QfhVECpIN0H68s3kMar4R3QLXr+Q8I5Dj8wzZa0B0ZUI9ibT6/2H2kginoyNTaceTEb
3JMXqck3gnyv5dmu1IUKASj/6Gn0AQ3PUUhl0faVNNmyAS2gTrbuvdmxb2ipTznuKloJztLAG9Qi
hKlqYf46rH6orhkh8hVZqgdzF7ZKSKj37X+dBPWgBMDHFAVYNFx3vIZk82d118ouuzCSpscCR5g1
hsPdHVTPJ05wwa1GUxFoZS99KISWNLKGCgY49svHw8XN02u01fmfWgouHc+Yu9FS06q7IK8mBbPk
e/nFEmZLT875+negIiR/HnXUBfSoSCkzigKcwzz+dvYMCFN/RINqU//OfLa3XsGCRSIXQqW4NwyF
Xr3+oh9obZe754ECYEZHgmOpOKKqDyMwVqJ/r2TibL+07OXR8ElJXbXDqSPJlWIy/hybJVotp4zM
JvY/9itZw5qoPzM5NolJrLA0DOgAcPuCdCM1sUrA6PcC9cAqrS6mxJPJkzmhRpNm8GSNdF9/qc4/
XR5HxU9MVuIA6XD20ulgnnzoqUrA3nrX1Mh7Z6DYAEilF1mQV5XeF+IO9duLVBuAemoiQV8WC+n9
m8yyxDKFEFigY324n9IuPwux0e/G+NT24PMzBz/2Ghlm0J2D/3j6j8/EQjEtf05+/4WmxEr6ST3X
WyAIWtNUzZRJOfZ/nygAuT9znRC/0RSQwuucgzPu9KetoNC7ax/J5som/GwIgj6ix7tnKsqbcDKH
ITcVh8asSOxB+Z5xkFd1i57bnlaJlrd6VioNXXqqtwwzF0lbD2+o5AHlxSQjtr6F9M1a+pzApGkG
0aMQodVjPSNi3hVw2d1GscIYQUY12ZwzSqgsGqqMolsccCxU/4cj+g0f/7ZmjTXrwCC9zoH3lyP0
iAbEuZT1NhpmI0PwaYXvV4uQSPaBVS1eME/Z4iTWdvKwcf5vU9hPP/beZgBAxEZBQ7bex4TzcQDN
tyva0/kxRSXhd25x4h/mMWjDdTbWSypYoBBwWS/OPwubff+PxsZu9EFXAWUDOd5NfAUz4z2czHmx
uDyWJqGOcy6QewLCFXwcXZSqvkfkBiw8zUofkWRejTdzsCiMx+v7p772mGGocjF32V+Q34YMXYDl
SIGg1uzSjzodnl+n8y5ACDf2FfbB6oi2h/A2sVfpLhEZxHBzEICViIySLaJOqnCkixkraqOjXeL7
tuHtUi6IhnwQ1mHNQ5G9D67+H5if8aklFs1a5pe8oJOuigpwcFsDMLgltZs7I+9wQG7o6OIIWpR9
fyUh5r95HdZVfLj5yaevmBbnIp70yqxJZQiWYF4OlzyO8uSVktsCu1RuFodb2y7Fp4w4uO/0wuEv
oNIfZOa531rp261KItGhGOmKinTdObCssK5/TKPbLW7Hj2Jy6ltyZHnmwOSBcgB2X6EnaxDy2qSf
Z2Zygz/mq3932YO1h1DABLjIr5aerYmv87YbXdq5iacO7tpLf+7E8y73XkAbyRSdWKn8aySLvBPY
9hBWU/mcA3KjXrjme4/XZY4+TshIJQx64L/LwZoBN0aYuUs/d38N0lYQNYcW4pqNCLLXGgM4vlyG
DwF+uBMHylOnimdtBvmuTueoLT1FfcYGEyJe6AtCGyJMR7o54CZ68ECX/M2kTSZvofZMxvVUlggG
3BdG4gRU++etEvZpaUu4Vl7KfhrvSFFwcJTTF5AR7K/ANO9pW/0g5F+NKY6cWMNSwwVQanahWDSv
2LaokAbomXbXTjBqJmGRrFT8jiqhZsprrScyyoQJIhnkSUufk+l/TM6PIvi6lVzA6rKnKCydVlf5
qU/2J1kzfee6H6szLPXF9vtmtU6BiUzqQ7F9vQ3KL1CN2GQG37z67FNAO4q555JArbhH5avTpaH3
vG+iwQew+zL4PyvsWKM7GQKwQAHTpGz+oiWR6QFHriu87uQBykulRwmu5Jj2Tkc+wRP8Nf0oKbTN
VdxFR7k5V9JxdefmG81j3t9e/W6hBdCkrEvChxGEw9S6m71Rr6jy5Cl/aZvwJgX/kR7DSDi8uX4d
SDMklH2TZpyv/L2NED+hPcuU1SPynqgjMBpPOMaL6lUYrp4VXVSWLFV4i64G4Ha4GDunU1B/3Qug
ObOJ9uwvXXhPeFEnXXnBN4oLBXADJ9Cif/1Jr+WlvkNh0pzLylD5kd4n/4Os8N0cTFmcSrqPF9Cp
s+ful37YloKknUOR92uZnnkHy+PFLdcaAhwp3jFckCDOAOzZ5Tg0MsPVp9d5xaoCUol8avojXN1m
5c7939L1M1dxmBBpZHZhH99LmphmLMlDFE6NHQMGKSQaQ7xbpVT5iNn0YwNhDFLD1tfEAzheV+gw
odKEQ5p8STH+Sxz76vN1qnL0gSuFdMs276rMXVKS2p/Ns9ZWtDjjEUo9XP6dfEmLmCYhXyxWZn/4
hpfJQOPpK1V8Tvd/o7rkIpcAWLDy75YoB9sc/hMhv3QTCZ3xptdNcRXtM7sMDXOt2lWtQdEZWlkC
xpOFjvw+cJZ+P2yYnWOIAOCjOTaRHkgLioa/TwbH1IyfuBuFJ16hkVUWOtnw4w5+ov5lVDTKaiAV
qByXFs+mos1qBlMo3AaLerxwiewV96ypCvQia1NHu6rnhvifi5JC+uP8NpPtHgdCxzXeJz6l5dZH
1/tJtFDQzeJIpQTLAQuyJ/z+cq2tCCoLd8GQNvVzd2MjqD3h64FRiVCTUp4Rj9Uxe5VFH130ufTa
fKqNDRVifvIEwM9PJKfjDQNyNhd4qdBBIiDMFUAgEkXezBirzB0VwjnN5hCGXeMoxTSEj1cOjyrE
lUOBU/MbVaxJwAZzGbfsTjFZr8oxd06zKpIlgtpZ7lTQDnCczFfNb6xDORu0Yw0GZjT/YZ5dm/6g
gMMt0T2vUSPTh842PPA0pFFyYdW6fYVwgE83Qgwiox7nsmKTaaUAhTUCGAL4yJOl+j+xmh9Xpynv
Hh8ghnCrdpmKSID9fqpmeoP34yxMlBHFBTDwQwBoiFWAmGTQdUkBksdBXlpnBlUAYjAyqVfvm1El
vm3xyt9s+wNMXNeFBmqKxBX5owFArZ14eExU9Vo+uuEs9w6ygm3FhSTbPZRyYXGKkAsIUrU5FUGB
oLYYhzZapQbTUczdiBJIqyZ7rpeE4KDZo6BdmAJKXnt7vtGmeiyl4xwj7AjNRTO3GLcCNo3J1Nxg
bxhZ1xDDbGBZQhBzpuY8ODJH1yikkArkNZoQi8z/knkDEfDTySTDLIbmf1HZ4SnwbqvIfGbBAg3V
rKzvtFgDKNLi+azJXQOwjUJoP3HaaEX64I7UNPHUYUe/H2Egit4bJLZdHFHvAqABJVYrAtbCe224
0CErwgK6FJCqGDJous9PGOwUwK/bYYirxtnh5jMMjpXN8qvDvj/vDl3Q8chhZUmVMEfLvtSFkO61
CjwPmwd9CiRSWGbm22RKhWnUZ4eR7jkJoiuQnENvRhSL3MLExN+IkhnufNDXgErw04N2PNL0jGoK
cUP+g33mQK0RvxuFOSvSZR1twKeKQ3I+o86YlcgUNoMvrEITv2r+qrhUJWHTtDwxG+IAj/ByNsjU
o99NCmWCwqTp+2jBaSyXyCj7+3N8TijYILIMluyfk6ckmb6wfYbIq36cEXsQPiYZaAQwZBeA18YT
5xdiPwLPGPV8mpLSH77aeMhAb+0NFoRH3un/5mhBn3ljSCwQPQUAmXgOutzNnDYcpbptdENh4QCG
CHM84cpIww3F/pgXOesY+gnRCv7pAwVQg0X/uXJm9OEO2kwFoF30530DrqUzsVaD+0k2uDlTQ+1p
3oj2eTll9S4loS8QWbAYYze8OJ+GMGVKSWT3fqlGXsXlRlDEaYGQNXzkhijpYB6IT1gp31k+ESWM
lWN4QOulnDaNrB/bjOWf4L83p2sjwFgL2qgH1Rx7PXuAu4YueqdWU5YhDqoGvH8fYK8abtGr/5Va
hN9BRFlWNYApASHQoaAXGjLE9RiWIYTMJHNRAM3AMfDRIN2RaJ37E4L0du0Ve9s49gD3UEfANzSp
gbDyCvmiU4DKnpM2BlMpHFrG8HHns4zFdmUxXz6s0ZQjnMOQNow9c9WAeYJRKIIjW3jThJymqGbd
NX7cxrxxUFCCZ4xJ6Rt/hW6mSsDgjD2x7gdD0q3tIksmjkhBxDxnrpaWuD/x95jSlt7KVYEmRA/L
bkgWQ/ify5vr6p7X+sMPUJByBpYkOtofQ0Mc7YeOU2vLirkuMdSWS80GHC08iTGD1kf5+vDkrizc
JdUWtv3QnNTdJhqIwxy9CQWMEsHDrMEG6TYTt2/NkR5Fx9/Nc4vhFK4bhL7Y10ofsKGMHZYh5vm3
4jOqkY14QI8jtWf5Q4USBTAisyt01fcq/oVyqFAtvaRX5rvFEJdAePRtPiyKOcw1mOab5kJK6Y1g
OJLbDqje1zDAQUHNl19ZUXS3t+qgpgmKSM9vIVV8Vs4MQOyVWFGm5j6Rz0J35bo+OQXpWbMnBhup
jry+OtgFQV8BNwxCd2fdr5E+1tH6lRC3EUpDFbWIRKLzgZ+I1w3NjWC8wjQuqkHvCa6TW9GaFV9d
kAmVn1vMh8HwaAOmaHKCpDJSiBXfUAXmBOj9KWCaQYX1l5FOxd84hgmJl1O5k4TnBDvX4e5zAHbJ
eBYmlVe8F5kW2uPtQgqHEXM9QVkuBN+zq/Iujkod/zYyDZP2EfZEzHrDbUcER4pYl3Hwx7e7osYb
qPBf29cmz4dMGRU/ZQV9BMKDl/qwJ28danPrqLjm46owx2g8/7R07Nk290AMU/9SDfrSbIiN/4ZG
HSiYeBNRSROYue4Xjn0HGSb/q2GgXHUMJaIfQbtqrMDqbIj+CPKzMEhKZt8SyzK1fXHygZDLMgee
vaPWR52WeTY8p214DZM1u8ge920bQcVBcPnCqeDaEIXvoJG8IpTaObiS7KO3wK9myKfT9RMNSwoa
57SekT30VlautfDs6BzLl8viCPKLc+A+LwqTyMZQPRImp0oz/ulgMH+ghU1+okAf/OEGGLsBYLUD
QsbbYkDJX9jTpPIUImM5oQdtWOV3bFLJ61CFZQkYdwDWBU3eGA6bYGNi/GHVcpCvPK661o4OlIz4
W027fot1gqyNBVpd1iNH4CuBYfQDH8OhlDOqqc3c3N8xnnwdybMu6oiAvUPRhszXP6pNK6vs0gqh
By2p5Ogfg4iHxWrdGVcBHGOGWszgo+aO4fAtTqfb43YKDnb1P8BMaapkAOwQ3mXZzNNey+YZ4/jV
Rfkh/wNmhSMMdadfH8VydtIzCfE4XfOnqZXK9qepMPdqwVmYsgVeYyqnLnKs/7EJNvfgTK2aFwa/
2wZKCAd3McNVLhw3bFLvgkQxOwQxiEPYAwAk90+Mtok6AvRa1ganQhEWTrzr3OxXBxEnMNp1HX7B
cAVIcxQ7nuNAqcwc7PzYP+TlwPgLctl8l1QzkvOCDZVxQx4JoOz8G8WXq6aaI70fe2vbAieTYw5S
sYe5F/3j1ktCkDeZCuwGLzRm3fYaIDYlGncIdo5KBavRRXrEDEXgPpBNZHydfAh0XJ6cQhNgyYr5
bP8huamlplCKeWaOkucx8U/jBIF1TAxkxRPQZqssqqgUPKxW2c5FSuMPtEojjhleSuKiODphghEq
6LpaoTGM0pYCxg7dPXb10B2kLkE+lRd5XzQ2Gbrqe4aYmAtt7kv+JFVkVjagi2OHPNp8N4cnuAjS
o7mcRFh0zcgQPIvOfJm35erx2Nk0rR2fqjSQS0X7XvoW2LKTd+ue64iPpJzK+yJh7qqDi2qjVw5s
EAzkkqmigMDvmOPE8H+yyFLdrEqYcGgUKNmnrBydUPLtdrB89wdVlW/eko5P0+zO/L0dRLmUU5a9
EJxrAl5UdnX4jIsO3ooNCMa58AJavx83LGngsoTOsWAGodmdi9YOcItERorWOWeIs1VZ94BQ2EWK
7IJLsmhaySw6bpC658wIMZ8dSiEPOzWhtsStjyEpXIgaPBJqjerMuoy4adR6dDSol5mqe/E/AiGi
GPJDoFhpbt/bfqoNY/D9Xh4y9tvl2q0NKHvOmywjBYSURIWByeB1UziPp/jIuHdehM4w3cWzLAln
fZLAUW2lisCxrW8OzVUmQmAyHOQSoJEeWWnS2IKFcuF/FRGZ8e7s6sbRFW+84oZTBaFM80WTAttI
tBVPciO1UVqcolt49E9MIVDJzxlXRH2xPJhsdXHmeFEfvtUG/wc1tSj60wM+cJcrP11fOFrNtuKM
7nU93PBjzn91DWuUPt7fsyhtKIEj9YTyk8Zx5CzyW3IWxD9qFQrOjEqL/Jk1Vhzc4Xgzfy5NnP6l
wRfUPEGQbSuCttxCwcySo0IPeUVQIqVErWLeqdoAqLPh2Xyf3/sbq9jJ7pXs0n79u30PeAdPOwev
V8hyXtbD0nj8Ou97hRDEvGw2DnTHr8xuwJcTdhxMn+9xY+fk0y5dHQ6M6DrpO+ryEXkNmvwfsvWq
0gW6hdStYoPU8HHUM5jgmYwc1cXgglhVE1Dnc/WKlu4Hy8d+CsQPPmBG+ilR/VGH6KzsW1nzVIGs
XSJpmid0tAJwj+9mZqJDavsovgBg96jXHbo7fLHgmaGk3ttBfchiSRwzUuSi6Iz8BrNj+wNzdUvD
8GBKueZ/59s9furYCP740cwIzcvC7SvDEaWI1cUaQ0yGGycqV0DiTl1YS7s5TX5ZuxgW9zNBaaw1
oFkY0dQDaoEO86k3swVZWHiJw8FDQvwu9QkzpnAH8MK4GMa7Yv2p6/rMfYUYjWpQVFVPLn92/E8N
hUuJ6Xpap6MNZN5TzYG6KRe5NX5MdtpWxx+cJCcT6y13fp6jTuMJpw9wz5F1MnnTd/S1XMCUrnvv
uPsnr1ATHLwQ6Dp2nOJV6uFwRHHtlPb+/ccbcpwmN7het1PQsjwdUoO8Tp7B/6XKxdIcDMVFchM9
Sj64o2te5eyPxVDfWEDVx65mHFoLuU3Sumy5VsGlLNJ2PL/x7qmUuc40e2dgoZZT7wQauNkyiXuA
LT7g3psnj3NLGTwq4ktGg9YoJE+NxiQ0/bRMzrvFrG3DeR0nC5lhPJjcggbksaJb7CeMk2RWbZtr
og99ZkfgBXrJFuvQ8fYLuNuvwnGh/r0q8NJ3H5OFS9KlhtDh6o8eTAyJ3Lnk96lJ1B0ebNTuhH3p
/3CykU56VzNZZYBqhmHJ+sI4Ky/i8rbfNZ/AVtqnsmo2IizJKMiQu75NY6mtAq8ukDHvGbiDMYZd
lM/84PIuGxWNmmqHz4P9CaBZX0f6mFGECN1rpZsLXf1B9AfM9d2LIVM/NksK5r6vBkxIBhmPDauP
BBzREhkbe8EKa3reVgY/5zQc82SJjIFj9nkVC3W2HzbQ5y4gq4Zqiitr7D6vIlx2EXDgGshQDhPP
FMJ/XkNFYzJRSG0PsGmysdlQXf5024fUaJz9VjwzmZb8rxxtJy+AB0uATnlnvPWJ0jlQdJjtCk95
19ic+7LdWDtz7juvTGZ4+zAHKbfJB9JK9Vg5Zqc0isW0J2JnPXHolqm78WIy9UgHzQdSaa68I/xu
K72PLFziNOopr92iosLde9uj0+ozplXDjEbx6GbtzjcLi9xyeihlYmMEq5R7vOHSLlKJhEqsxCfr
92gJRaGgF2Qt5sKOU8F41f9qlMwENpbyP2I4K4guvs7MqHQmGO/CSCgetVJPUXOaNIpjVFrMFm00
2MIRUBgLcytiJItAHK6y7J9A8gBUXyIl7h+ShfePTsRvG59+kIbW2z8Pg/1XU7crgEUI8Cz45G9M
FrtweFEmhm7F6NYSbg52yKcub6zN9l+a604nIyGLqYyIjmuUCHAzXC5KXPrS9DdE9iLp1NDJN8+u
Yi3OeeMynC61imwPSEc9TfYtlOnkRWS9FDy14AmArU3sq19WUWge66eq5nVjTqvybAvrg8W6tK7r
XW6UF6eX6nzwzX5VDU7pRL98WiAZU5fRFw3D7e2tPhC4MDAaRGUCgDxiIDc+SBfqZqITYW5wlWRA
BhXm1oXnhmn9M65AZuQNPqXWsFUiIPDZ4vfaOeKfachmi8yVbcCQfRSIMf8eYuThwSDz77fkFGbl
dqYNwVbqz86UCgRFjpUEKx9Ui6uDpfZM+DPUTlOrUCcc++0O1cH734W5OXkQqcPa/Qk+6hG9K3nT
D15G0ATndls4/qH2BfTyUkdKFjBtsILfvIaWGtvNkJ9n/XXe3tR+9DsRfzXlsAce4lACA1drqxnu
iyDEWXO+kmfwbdXhajNnu+jTRj6BBY+XXIICZKIWVtBFI+kUx1JCRKQRTcAgHoXDE3DQEg07tDz3
5EDUg+Ye3J1smOH9UG6dMdH4dUitdShFwOX45Mx1FDSDrH3cZu+++Oi/emm7Sl0Ux3QhhJyRrKNF
uPULW+4VKOmi9DHeLr2VFmoduWxHZFb2U18WoAa/VT0ZRUf9cvg8DUI8IvnU9yQOqGHxB7IPHFkq
wF0a5WY5lk4k0oAbh3WFifC2fytX9a88347bAhDzK4ZgDWT/3FngWybUV4HhKUhVPWo/n90aq4Y1
ZR7RPDrhoDkxRShctB3yuYaCKow53NwLrX0q1dWcnu296TCaMvBW2gFehHsVbYBjmDDvRpDwL3xa
glcktHjdSzkIHpSpMhHMGqEVXlRLvSWCDhyNr8JzjjyA3ROd8UfC1vnDCPzco/lGKHCfxC+K7ZU/
eJvi5GIa8JOxG0/EHVmpxynBiT8Ddr97AENohw74kYa6lVTUwf/I5OnFxpVP/RAd6jrKz9NxVj6e
pbb0ECPDC3yXHW2z3JYszl0xTW1c3omzM+wRzDqeF89KpcPZs4Ora8vFHohE0wxlPwTEgnbmgykX
8FwoY3k+nmj9ez4ThS4OBCSkRW+SFxcsI20U3NIzxiK2pjLalgPVxyCCv9ZkEMQHN7fW8mnJ6E4R
U8tBCKTaAiYq5OnoMy8cnXzWj2ih+2d9Qu1EpgqGPLzULf+mBZRxUVf7LF8cDfRWwlsCw5BFsqFx
dZjOoViQNToB3FJ8SKYWx0pxERdJI7dz0JBOEWTRlsDiYMM9cZBFapKjqFovEYIFJ0hgfbu9GRuP
TVNr3O94O5qeNIf/9OuqoMshZ329RAu3MidZm+BINtyrTaaDCaL61a0C+AGZo2F7MgCjlTlycM5Q
en5VB6JAu+gnVv7tCdenqKYdhi2B0WWrP4ze1SaIKfD0s3pl5pJC7Vql8z8X4LVKYS5qzMO9tLnt
8TZhtPkfhXliytdBtaTI1CZHGFcFNfa7tb8DLFAZDC9k5UsDpMKHfTlrt/cDzwDHcvH3JdX8QSNF
jmzG3TU2avE8FTmuWkLBSupGdD0Ohrrm4OdXLKUOK6NjtFaGEow1FTioF3B26cicYL2/u8iZ2sKu
Si/GdvK10S5VJTA2A4AlgNd+/HdTJPRLnNWKWIfTb4/+boDV0g/m6VKUNwD1py7oG7xL7auiw2QW
LDTHslFNWUtk7Jm+MsTFlTV3XFemJRTgkBMU8pbp4oPRWjKEGcldrx9cTrVsIxeWl1Hw/1BHnBVW
KfFuB/lOZ7lgKHnhjGLga+e7HA3ElyJAlflUvgXYZGJqFCJJM7CrdHKHnbAQKl17qWDwBqgm2DcS
fXWss7pwJgrE6IAb+jEbUqzeqLaqEYgKxeWDNJi/42B0Vus2AGzf2SvV29tIVDSoADutMgT/MlRZ
U7jm0uwwSAseg0AgJi0sr0uc26XXrznMklv+k/S0ptcW42BY09dWZ2nqzHqD6NL23d5CikcTwKvD
QryejG0m9YIxptf1ndlOPJlAQjPuM+SDlZOefTnJztwdAu8Ws06uxA8sgMAfqHTdQhm8ioHTLwWN
4xVuhWDWP3rfd9J1E1wbXaKWX3GRLsJbaTmcw5wwMeI3elyxI0Pn9eaen0AmtKrha0VlWzf3R04A
8j99Djf3HOCNGDfhNIOw9jRivwT/pGcJYl7HrXbTdeirk1no3d++nhhDpBA5BZXswUa48eQMVkkX
c4ex1wfEfEhc3taf9E0v7Np84nAmheJyQ13qZPT7pz0EFVYzAx+EiapjJnS1yw1MzqhUhoqHMysL
8BFbGo1r5WAZN26BrwECa1W+zesSrlHCeaHD4g0AdgcsttJlEpjCA2q3GODGMkkXUGSYQMBHtuxM
ZGQg3Hm11PzjccKTUELH5imwjhyhklvryufdHlnbsWdd9mqyyBCrqWJTla8IGyucCFt62RRXw4st
o3e8CQLkp3YWS6Hd3HGWiO4qOoXXCHBgdyOx2JRW5NDD6yFnekLv557tuqjSo9BnomwUqinlPFhK
C0fHrRprLj3bZ7+W3Kl2mYxAZlOcMQaw2m8hu6EYXdyRE/8VkdpKFK5XHPeVwTlfVd+LNxTXD4Ek
mFaiArmT3U+4AKEP8HYKGZtVJakxc3azKVEMluRdD/3CzUDtuiVthYoNrSeOGSDQ0x1VTLDpOxvi
6XHoYphhYf7kZjOy8KkUZGiCTZhBi3J1ZbLHwUtaIUU+iCW+kSEQumEshlarTvsvFKXIKMyOf/GI
jz9vtFYsIwqOvDbIoilew2oBP9oVWUqAxGAepeGWqbwpPBaoclRTsv5UCNw2VF+aazbH5oyH1xng
ae1ORTaC4B6P0ZB7HwgYR7S3wUkOPesZ7OVnPZ/SHXJX1KdfOolAwk5ccmiJep13NZLSAlncmhaS
wWYZUGKk5iei835wMXIcFHV3F1InYpRTfgXqWmpxDfRvCcAxErmYhBORi75nFou6ZtYtMehm79JR
Z53yQ9FoXVaEXOMDhbQBWJGG7DfZ0L0YpTfsbkx/y3rk9in+dzMudt79upxTnwLSXLu0Db/isZzN
jxMEllBF0xcBDHKms7u75srE9WnDSew4G9cUbT1NHQR5vD+SKLDHMUEmGpCIdGhhD4pBsoie4qdk
m+yegjgcscmDbDj6vTiakejt6tjjDMzjK6UXdmjh3AntZnZEleg5wle/KIACPJNes3IGXp5Gcla6
vc36tNWUzC+flUz2IrmwI7e3Vr2mZoVjYymLv716Z786gv4DhT6Nn76HJUDvCLVDtKWd/q2uLUF6
xJXt8+SpXMCodtJAoQ7Vb8hJy7D+FdluJF5t4Wcn+GQrEVerRRCHeVU6YHIVGnHG+suRc3W3HCcK
gfgBFYOY2PLgEHfIJpWLiVfLswVLZzV2k46eyU2y376rXK1SrKYwwyUmpfL9toRIoPOG+U8+xDWm
lxSc60diYxCf5LlHZeJ4LVeWkF8Gafe574TkiE9G0cjvtOcNFavaprxyiwyan44AlJIdhVyIUd62
1ERUoLStu5WVtszhs9D2SmgGnts0qj41UMnWMd7YMsJb52km7H03KmNrtR91eMxmjSTQv1BE1itH
av8pZpBcT44aUYdifrnEI0PLlRunkHW02cvkfHXvEWn9KNo1rLoU54mfy1zPD1t3OMdhTstX4+Vq
Yums3RTY8yO2/yDSFQm9wo4c5FXleC/CaO+lGujgtpe0HpRa49e4h5mPnToDn4qnH2/yUJsol+5O
RlGPWXKDqeMWake9bCmXhjNtcxcQZmKZo+eqdYdgFyKSW7LkMFzdZF7MQHtI6LJhYTHW2hCnGN+I
ZLeG8yHkS5+4I3YkDXcNXk4k1syhzEwBcLoFFQDooLLcMx2UovvfY3/yvUX4sdj0iFVVAs2APY9R
3/Vb5hbPgT0Klm+dLqtVE6ObVt6aEIKS6hVLGw6J9KtxUj1sLIMl0a5w5Y6K3UbSrXjV+4BBpmGK
qCe82+FCS8uOHHVOEHvMhOPZ1ICXT6rJuD/NBirCdaEcio/CMjz1yN6VLIkwQwCbFrGXCun04iAM
ixyh3k1ZU0wNSs1/gDwJGJFEuyEzxKqirm5IYgHh6xbSLNUMpeCB4xz0sG9lNZq8+wr5EA+bZHz+
ccxvUqF2uyVTMD6eItGbUN86TNrigWR1XOOKV2hhXQ7Yo2OL14oEFRpnkzRKv/Tj7a/b1WP/LK30
GXbCDb51Ua5hoG15bM5WxtmHubgGDBApnV3CdFQX3FwZq1FaWvK3Xv3wz7+1G/IauiYvMbno72eA
aiAzZEJ+lacbvMENRMaSCvhMKCNyd/ZulxB7wOJ8bMA3hKWtpSpeg8j86MYWJv78NbhEpcme2BqE
8vNVmcjRuwXIfrj9fS2Lk46p6y3qbekFEhbRClvpB9c9VHpV4qLcN8pu9Vb1a+fy4Fi8Z9QBJPE/
wfOFOvteQsv0dgbLAywc0COAaWxFIqsBihxFxJEpnbIl3clDXE579UbfjCjNGAiPrVT6T0Ba6ztf
no1jxAPWSWADJAT5GdaX00sgAMWU4IEqidA30ZidBC8xSzPnMEji7N9GpUQiT7ZpZjszypoVY4de
TKKrDj/Q2+9rPjqg4CxZyRuXQutUhp1rBV+rv408fRpaZTNsGveUnsP8NIY/itAqMhZC6z6L56BR
aWIEYKC+VaD4OwRDIxG1xVeKLTTT+ItiR73YYQSpV9FnK1xDjC8zFjKTU3aVjvOBnHJ5zgz1TN23
ZIQeJUuoJ9Ab8TRUgYxlLcS7a88FK/XtZ6yHMdt937jlVkpBvIArGY+mf8cPDhAMNM/tuygFLTi5
4QvgHyxMKqRgFSl5EaxAYqIG0EJyrPibUsQ9gkxXUc2um+x1xAbJTE3IPZRqD5R4ksk+hnkS8ozx
av3YnsfX7b8DX4vX9kiq9uv/cTfXnosHJj6vqJSVhVviRvS7V5iJbGIfMStzwlOwPnpP4R0h997s
+wJxZEmFo17pkvY4/Mj3WHx8oRiu1ghd42jyNo93/yz8Nl/VNMgt+W47grFWGXTjPAiZs7Xf185r
lkKGUgALjiY5BRbU2iCCb29RGCjGoo0QspU8Ik8kMXT7kJW7hhLodvuo+OJ8fd6uvkclFXpP+14p
geNxwkN+BSu5DQdNKGj7w5B6Nq1nzt4lCHPubyOWDYBdKOncz0I/HhUjzCU53sL5TtifaqA/uhy8
VbrSHSRIZAa16uc+1YBVOHdhtCdapOtgwqhSBaC4c4anatrhFhdLfaJT+aqmqQJBc0Msk6kpfx6t
3b4PP5G6QV2Rsa9eRgL90rEqqw/4uwqfg8l+L6BXNkLMQfTeuLphP3Pqw9nUX8hlDi7i2WPvAcLF
hpgckMSld4pJ9pVy4XvaxDosRqBH3Qd0qZ3fI9QD6bRkMwr2zdrZsXdk6iobrMPYk4KQj9WZHOpL
26sIFbGtxfyrLofHHehSU5++cWKMn01DltDgXuSsqgFa82iUuJqJJ+Hh6LBtcXj+CxwavUoX0HzM
/hzDNWDGPVyrunOzz/ysThQ/lUjvcAN9qCJ2YqxeyjFjQUORqeIs49MyzQBLm8ZmNywgulPy9DDt
U5DMuA5YQ23ahkKOcsz/9TB0nukQfgJvJ3Sd/rdc/QjnAR00QQxdq0oxvdkk+C/mG5nJOUv4QC2p
s7RKYxiVIMcoe8Zd3VAVU83akvM6uOzBBMERm5gjGIhnnXT9wLNyXkJZlq4UvIPdHDUEmkYleNFq
euN2Qo2P2T1BB7nY184nh2RKapH368RSClIK1LuMtkIbLEAWDEnjoD4b0wDkEdn/d6aLcR9PGxlb
qQ/qlBlWg4pDeT2mLd0pb3wx0qw/qh0bAehs7PmxNMPZxNjSxVPOmRbZLjHX7z2RbUqGH8mw0QLi
H+vTigYKpmLdADWEZb3d1iNV/8VNR1T5dKtPFB2RJ0GZai6KtddtoVfQRyE0AdQc2YWRjNhrzL8e
dSjV1gOAoNEzYGe4sMwwtMwxqiAB/hGSUodf+fCRPMUTpQITsL+jX/uE9X6UzPpbvC9YCgIZm4IU
l5RcZoRYJSu5/MwMPlczklGS95VplCywd2oXmW4yZB3KRpPnjQJMZ934yxEk6aoA5Je3t/4IgX2d
0uuH38bOSzlmx40001WzLZo5jImX9qj6XJvZp9KOSXb/0SHTdN7yoeOJrJqWL+Li4HxVO/Y2MEAF
32rOxLwIuBmnPQzJOABsW3/mEyolzFEp37BrVgizKCQIlobcptQhGfizSwlpIpzzhZobCmXGEU5f
eWq2i07jsoFenIcTv+7YjMXAVH5KFoa0Gw7BT1Qf1QL671EnNua0OgGy1QB8UuXfiMtbLpOF0g7q
Hz4kWz0cYXxgCAAJx22wNZDN0buhKTI+SmfWuFwThUaPn9WtoxDJxlFXfljRi4rysZ07iBCrHky/
tXZX9+uR4ed5rH+hL1pLG4MQxW7Ed+BGJL/PfWxbN7MOf+vlUGuotIzhtmAAy+hZFalrA4q7di/a
gSreeLTLov4fVAXosU8kwzCCor2UFArS1NZjPTzIirAepPuhAdY0rsqR4YNef7JdfrUyetAPwbhp
KYGb67sZI94ZdHn59lgJoRTYJoAkJjUHUhOtpxye25K0esCXm56Kqr1DUgKRXmdE7cqBH02Adv5K
0JSuNTCReXrHA3grjICLqPBnABNzCZkiIh2RO1FJLIpiGQE1Pyj2Ac8cXJBf58/dQIt/+AuVc5iy
3sNfmI+6f+eZoFchkJeKMvUKdfDn9R+Ii8qDGBbOxEH0IFz4EN5rNxXzX0Ts5UF2D8+ayXxJz3jB
xPxvL1QKlvL26nJmDVLmAcCTf7o8JChDl5FzqlvjBPzLeB4KIQoFvS6QOGtIdyfjVu/OXq+s5Oxh
1eaXpRSs7XeN4gOfTEd1dv51JhzhV5CAJsyFwO/q2/AOVzo2W4vnpSdc6fSf8tYmxjMjvAjSNrvV
2hKAsRXMrbc0x8wAPhKLFeG2LdNqNE09VFgvJGxWR6uma1WMZfjQzbu6gXQ9AA1z6qS8jvNvIV7U
Y7VlHed8YMZGS6oXMObsY06lBk2BUD8Z8szYA7xSGzHBkehS5lsxAVGTKymOpFCmGPopF7w8TaTr
qkvBLZkSfQxRWUfgsGTiQPwCO3K+LHC+C4D8ng83Ko8MmjbeOaW9rbrNFRnFAHJ/GFPRuvkYMs9p
MMdV+lsistUe2oHj4TJ5xVtPtHdn/Q29CV4jH27l4FbHayyemPj6KFaNBKvklfiz/z0Nlc82ah6C
YrMW1Y49/EnZl9syWxAyMvQ+C29ZCM2fnWlj0qx1OjXSlMxoT4cTJZip1ZALwVFUFR8/DJFgFfcM
/krmG3oJAsS0p6kRJSNG0I3bl576xAKfl792dwADylU4OBEuSKmsfGd+j+zdLGOv4QIu1ymUpsv4
J3ZfAeBTO5IihvOowjHULueQJy91UsenAyBEOoqsaLTCP/Ja6l+Y2ZFHhaUbqkyr8OxF3rozhyQj
ztVqlCZxS/cTQRIRtAqeMoePetyG7JuKS0k/Na8D3A58qghmrgQE/lAF0PrmA+/UVDLGqf3ekrd1
4tHTozauzlF8s7GZsthVBmG0p70z4AsWMeihTeR3bC8pVKyksUxSKDqctwn4r0SgYqgE1dOYKgsX
Dhny4xG3qlAfa7T0AINR87vcYZq0R1tzCgnJNVFizW31VqiXcbjprc4gEphoxu/mtBBVAmoHy6nh
k4xFq43hP6WtDsTEyqFC73IGOlKn9f+/cpbviudVjoRRvYdn2tqL5VJrg6gYlXQn6tCAo5JcDL5Y
84J5UljENDSYImd/G91ZfvrMwmQhpI7l3681itojI6KANEnaDl++HnoYaoLRgk1aPhgJdbhlvwlE
CvzvaLl875qJm2TBXKlt8aempZOyDnS1Xab6rB32ky6UoXFeJaTJRztvPzCPsgmRDcIS680VI0KW
C6rkPWr9oz69AX+zm+2zOSt5PWEkAfIlyYFhFBSWvBiGXopyDbplzMLK4AmI15C7W7vXRY24nRPI
rXnUUd0kKcU69/jjxCSI4Fjm5zvvcdGlC9XvaeKbOhl2hYUNvpjukpjwdPg6XLRtSzgoE89+Lb+U
x+TT6mXy/lzzfCdDbLEjIx8Vp1OET/SdPnWei6O1vMXuYLWfhtEC2CwkuG8eJcD74lIAFAtN/XCD
/yB9R2y2Y3Uq2Uh4JtOoCxpk1Tq/Si2afHSdWtncREbdhDbtPus3MXwLLOFzFwgRDqo/otitI9cZ
EYukPTj3sJtSlyJAvGh3ccW4p5hxphxpHsMNy/dsjkolvpE7jfD3mnbpMKphg8SYsmEFTmmEIGqP
r2gVw2eh7i1OAanV4B1d8Jdtx0GT5IxPk9FN9BDpLJFMNdfOipP+UkxdaK12+olNpyIV560zb3ho
LZ778b4eTuw2EJU78GWa5UEGOAGYEgFQEr2L0RlTx4tH4yAtNvfeoNNa0XFALT5IG3vgQOcNp/Bx
LlAk83oE77n2UFcUokwEHFCuyGsOJEWeYAgwnO+s244KR6/fGFdnaVXdhBYKKBdhedGvPri7dCr8
atkvTw4g955lXQ7ZdEvL2wmkJxJan4MFQXBOIVXYiclWlx+VTMgJiLe/cMCRhBh2/l00kjpDZ7gK
kkzzIYVGnsIbrzjTAdPuofM+dtv7Bn+Yk01eaZ1uzP9JmsuVnMFhpsulbKLSRW9tkUVas3nGadRU
De7sUs1LC40jBcuuf4Q/H1hWEYkIzDNRXqEh0UAXd/IuYAytupPQswUymc974EQUdZau2OPfoGbC
wNDpBC1zE9o2H+MUC7bhHl6SKS0l43Rx21sX38YgDzVsItuvWxc0BjeMzpP2gC02f42wV5615cN6
JiflF72EoBr1STwZVgJJBYmhlV3oKBuPvAXunjvk27xPydr5u37dpM46WtE5kI8A3xF10dsW0FQG
q8RRbLa7vYr/gKpueRYCId0abt1Zoge3WIBKumDIpf2tblUSR85uK6AOa4APMqmCAJbpTitNQYVc
A9y04cjU+JIAJYspSn4VXEFfxRD/IXeYaS/6mjccMmEZlRerVYlwf9Z1WenUstDnm/RUJQzTCybT
Z3wP1TbpO6vxy7lXmbFRFU+jLEFmLkcM6fGlRT/iBTqGicsGqVlcX1DSs2Kq+PivkvKmzGoiznaJ
YXDUcG5q7Lt0LywpnyPc2l3NSaS4uXCZvgPjRx0W7X8Ogz8y7lxCE4sTWSvqZc2Z4UVr0uLqX7PW
D2m+WEyU7Q2mjRktuQSJfl+QNSfZzx2GI1c4Qmx33O8JMCLU9aanLUUAUDPuMVOe7QRBAt2h6uZp
qmP9qovV0+1gSio79pFrMQPMZcJ/pZiPMJQiz9wC0soK8/aWDe7jFYZpFwzPWsPK3vOY0RZaQBX9
I4MHl3cxZjj34XnsqnUDAizguood3BP/qc130EqHFLM2Bz8IgeSpk2fdefV5lzPiJ+0i9MLI03s0
84KdviPaeZmJ1T1vdLc0DD5QJwq/jS4QmsMO5Cr1kUGJrKNmfzWiNCZ+YLSIqe+2tmSAkswXXKkw
BBi0/UYkNJuVfOenmZBHYVk697RWxtTnPoBl3xOTBNLzUFMQ0zAKSW/ZYwlroFX9TN1Ofrh/6/Ic
35YyCJ+S5OiQ4gv9RvGtHSuNrVtxydl4x0OpVtcH3z5y5Yi3XrY7kOB/f+6edTKyl61zUBkcEuDm
Zorg6wE+adMq2n3EY3wMUqHXd4hCxohmPtV0edtyF0VwIEjwyTAIoEjh6elHWDFeRa81a2O3l5zq
MLe0qTERZncNHP7oWWFxSd+w3qKsv9zZzQ7ViXYRM5+Z2IPAZz7IwGoZK25HDrW11P+nF/s3+VuL
y6auqLerTe9e46wSHZ/FrBXMwBcbC9IVlWk3ySItcXq/SyfyJ8yBYOU5vDGGPbxlRXmo+/5IrqM/
lk36iSJxoHnYyZW2BUvHkYCrIvdtsGslgS8L6gw6DeVop2hgJqSTE0DERK2sxkir3AmcNRSpTFKN
LIEUr+7J2WXDv+EP4bK8l+CbRjx1LDSxi93bjiN3Z15FDyvDCcjWkDZhDBCjuXr0/BYGnql0IPGL
pLVVyJsPF1LYA8yTSOjtPHRCcv69UOaGoj0rIhjNgj4QJhh3wce32JvH8fmF2GWZdtkxgf6i2gj3
6xSB32vwUPCo9WbPASRJgHPeU7hKZfNiU3aTuRlWqh1TqOlqdf8SSC/w/LZBAPY7v+g7Uwg18I4e
7MMr42dkJDsJOdL6kbQGofRR6SEyQtGid2qh53anbESAMimZ3EVonEen+Mk7HGNIGET0t9p7JUq5
6kN/jL07R8LhVhERVIHCDcXHlMiMy7UAx4f5q1RvsJ6zcwoWRyn61MLpA+U0yvymWnmsS/eAhkFN
mWB4i3AMAnBsDMpN2Z3cSERgMx3na9koLQPe3WKf1T+bi3+l48zGdUox2oJdtq2lnxsGLOrnScSo
F7cjbhB/lbpc/W1kGWu+a1cYNbtV09iUQbw5Sk6YY6YHdbPBKOcASYSumEbVCYw9WxrqKueST4kg
tJA9/NfLQ1us/NPrmmGFyr2Jg7v7g8Ce+k8lNQqY+ZDONSh3VH44objhybLg+YBGAL3VafgFOiJq
ps1xPZ8hT6T3lC7PR2Ciyn7GosH9Q+fP0mbvuPq3dlUmjDS7ItHpdQymLmkHyTZmOtFyQkhz4PZ8
2e7tiwTtTaptWF2NdhtEbgCRW1+M9j7Y/hDsGu7pHJ18KPbgj/OTj7oQlGrpiMOsy8GXfJf2wl7O
l70m03/Ntl9IAzJ2VDIhztdgbvPAIWXnawoZi38FSvyFOW00S4Ss0jmm1nppDE9mgw7D38aHKmZA
VJ0od2M56XW+ti5kFpDAbtvJ5SoTV8d0KhuqHPhIPMhPL2CULMr2kDHiktZDc5B9iZwBozEermKw
AiVXXYEAlAtXYgSpMAkUy6sdUlYlNPWp9ya7+3hDjlkC1A+tGm99E6BqywV7uSzK3zQiaPgIQocz
mV+THnuYiD/oT605yp6qKPDGzY7IsZZXdJ278w2fnCVSJFX6Gzl+2RnTivzz3qSa83oxOmeVPnvc
PoU2ZJ7Q04v66wbxtpA/qH6a/tgaHG/7UbRemAbPnoPCrDaDKWyVkwkQU5OzFD4uSC1YfZWBP5Dm
SdQiR3EnGSLgjFeO7zTyQGVCEkBZ1rZM9z3rdHYWxWJHII2atD42hyIvRlyvCuLbYGPifgKqE9Dd
XIA7p+sGXkmZ7L7qKcK13K133S1noVp8+Nu1xWUd+D7CbXWv2e3EHKRYvKXCxBHxf9iTujUrYRlw
Z+9LKRj7x6E6e1e96O0RhmXgw6rfzt5YBdCWDGqtRyi9DVlD2mIp5DesZAnTJ7gaxuLN+BTRG24m
F0SgrDDuJrcpOpYN49CwDX4SBtNyU8MR2Vb4OBbIpnNnBxmz+cx02nUbyILrcF5MbaoSCwZM/uYd
jSQvHiVrLfBqTOLmzR3JxxBMOOqGXi/H9M1/nRwUd8cGnA5OvImu3WenmgfEAZ/bR8otRU1MTv08
kda7+AKoTR5Jh7fsa3bHJw9NgczFYexQSBW+lSe+T4OZlXTq6SuyxmZ5hkmV6ilkyIRhcChgrZ6L
hH2hPE8oHLaL5hcalFJBsBltdGRV6jsO7h7syqUEsEIXH7w0nQBF6Gu7gprgBGierLPW/GBg6WOb
Jvk6t/h196un5Q8fRlrHoGtnyHymYxqcqxbm6RabsgPyY3bHSJTea+o+vwFzdq4YqZxjMNwZaLPn
oCcwa+e75/EIMkyaXLxlvMRfBTR0bWa8omtrS5U/emSc8Mj7EMMvqv4aByQoHYjeWduWUuq9v3cD
t7RZREK9Y1m0kgBtavM1ccxEwoo1YdTg8SUqDZtE6LcdSixgB0E4O0SsagLsQyjJqWZV5CZa2SKo
CkOGn62zbR30WuxOB9EjjVDizVTMu3LFOAYRS2aw/JddwaJDnLc7zXHzQIRQdNyMcTRL1L8bOlgc
0KABRJR4nmox5pzoHJVIfTJpvZCzTFBSxXZXBUTmTqcYfIvos4Dh3mJR/gmA8Te78b2k63fbOWvp
N6+xX+XxLHdhmw9qAsERFXPglDLtStZ5hHby6CCw/iMGkir+xDm2zFBvksu1w/oEePm6P7dH8+C1
JXcLYVGnzJd22lx+kCfdBsCjzOKkF4RMA9aDmAHWpZk6qx+t1nioe0//GUWI7/t9WP9e7bndv0vC
r2it+hx9XixnIeBIYJROcutn/2FZPEfxitbWN7azSSeD5t9Y+Q54mA1PAdBmOPhFdK4iZQydbHF9
ovtayH/z8E/AKXRFVsCzj6fdR8Z7Xw079p7UXHyKKDthjzhsPIwaFxOhiCgGVDPfuhZzBzkUeNj+
GE7TE6FWEFjUBFvITis4hnsw5Y26OocidLzqRKPa6yHyu8IAk+b6HcqseZUh7kR0yW259xWCqUhy
3/OX6s/KdwwNFY0pXuD+TcXuyCg2LjwN3GZWoxq56O+pVQL/cmH9Nk/Sc+8xTT9yCpJ7lSpqFk09
kcVtNWQx3LOqboUjxnAo0JQt/tXDAlnwnXmhDuzOf3MhxxpcK6mGh0pBkoLVZTtCfbfT2xNPEjLj
jpMHu2sxhp/CPTnRPMk5Hd9IhpIBPL/i0H/0NNFJ4tuRA98WHbigoTolJE0kd/4hKEcyEDZwQnr9
UByccXnlR3P7xDg2EG+BHRuxhKGIOANIlV/p2UhuZk0+mUNc1hULd7p4AI+1LQfMPEYhp7+y20C2
NxUMC041qEBE7CJYv42OnlG1cPXwRnxUmxvgsQRoLnz2wxKe58sX3FOjkfu9FOWLoP5n6Rrh6ZQc
sgrZt3DI8kGPrgSNt2JAxOuCS29ajAHXQgodBt+ma8nZWeWt3q1fG7fFb1/SiMdwqYioe4VL2tZS
xrIN1dEWwAz9J9HQIbtFGG18Zb9MpZK4DGGFN+Ct2MlYIbJ6sPGhUkieBnY0Aem9NuceZQdXndsZ
+lFwVahCqJAYD9KyaCRDGyhs1UnJYE5e7MPUY1uf+NhoWgGOxEygYJ7almICQa2DxbEmsxaFaLRs
E0319kSPhkMzePSyOWHYgNtr+Upa5THlAjpNC5HpFXCsBI5g37LJvYoD65Ez6FYXwlknMEMGcSHy
jobzaPOHW17cUE5m61EwR3NzMcwU3TNPkYyU3GMZzl2cxL7vnMGBN2DzHjTaFN8wSHZk+khQwyNB
D9rpMt5CWOmkflYKBmgM8ZRQmeLmj+yA+9U9GyZYll4K3OB1U24yFhJNL8r++D2ApGpXWYKs12xo
kqFi+EPJh4CXVGygl3F3KBx/vdGOzc0ozgX8KkhFB+LIcVGk8lS9JlSISkaVtHbufBK2WnhwtLsl
CX1PP5YRFBsAYB//b+a9swYhQ9FT9jNkemAQ1j1m0B81usX0SBqf+Flx3zH59R3/B+m3gTQMwahw
uSvk/jFBdMr2AopC63WKOUIg2sBkozFoYTagzWcbqjkaF5UVLtf+5HS53bEptDraarrh90iNrkMJ
cEoxt1JgqPy7CJiY3k8Lpo2u5/Tk2CT7gN8m/0OAHe6oqqz2gpt7hcb2y2OdcvxxDlWzAPckBbnr
OAgKqx+qfYwB38i/fi0olO5fw5nal5P7fYslJGzhsmkEGtLs6agX7TV2RjgVwPW1OuqxzmgidnsL
S6XNjrAZU04x8I8tNV81YewWSKKfvvRJKiaIsx+kEyhgnntTL41nkfZwbXQJ7T942hmDarmttwhT
hJw70PrwBT7q8Di/E+uPF3qU47raCUR05obUoEdKRAJBGAUeEzrOhxVVyKfl1xzjahDE8kyReYIo
PuYc3DtCL4agi2XYiy3zLqX+EcuaTmgsSEmxZuvVx0McnBXWRuwke4qlgBjbBzHHD5Jtb8j42f2m
KdOkZU+f3e46HFbpdDN4Hz1UG5O0havPlZ0OLfyfkQ+Qkg/KmOQCtxZgNdSze17H57rqFzoRNbiZ
mXJWCD+b0VIGYld2nsXqpRtulNXeRDy71txv9FxDTINgXsgTSNcvgKezdcEgO1zduTKNd2Afwmgq
KY8Ac/tcHDfA//mHJATtrxtaQLfO4BQbjZlZqz/WvjXPrrfOSch38UUVD0ESt9VQLzP/5jwCE1YP
AGII6KLnkN8KFSAMz7WuSq+AjaqU0sAmFJlndXjixWGGkjNPmq+SKGe+9UuK63LYK+Uh+/MXVJhG
74wdUHTC8a+im32x/tIRH6ZwONKLuzuP2HIUzpV4x7fm5/Iv4VUtzqDGJQMRNbJhqDz58pXl40fR
mJSsMUBVE7xpfgmwUE+DEEn+OkETjx6cNCKuAV9ve0jyW0k/ARLB/bxbcxtxXfqRUgCRuxSWTQ1G
985QDebFOJFj/fIFYY0fDemZlPTOAPST7u8CZPugDrPJxmLRVkGsRnLd4A1YtzamSy9X9ncMO6Og
eEkKMWvNhcZd9+lxUxleifn89CHQFaSOGPBgCSLbVsjcGj7OfTYMj2pTjWo8Mdjh4XwQ9IsSI1k5
AazdORPIys+MFN+OQR4eoWQ1oEuda2S1foYMtNQfz9eg4Mi2ljC0XW4EA0Avz99WSsd+sESEJLEX
5QV2O6JmsOJY3ZQsosWC6rsnMC6KWEVlM0opWSVmx/X8ezhve2C9xsgyclOZTaBd3gWCgjKDtsCD
psM6uivMqskW7NwzBKvfknN45uKmBgFWQFLgqNl0hgYGSf41m1sp/rEw9j+F6TxSqd7oprl5RKDW
pHg923+nUSH2xyT3CnXM3jydVQF6RG5Gqtn3jL0bv8bHii4ExUPiSC1dRAs8IOPS1LVuFujCA3hy
C525LxNjb5l4hvfUSemSsdt6oWvWnoeJ+YvsOVVrjQ/gGLLuVoly4DCPZXMS3HxYxIZmEd03rt1/
Zq04RhGOeNwwRmJcs83HWVrqC7QLZnwZo+2E2VzmC3a+536x6ZCX5v81RsuC2rspDg9QSZJSex9C
l2lftREbGijnHi3O9NrTfCtXgydwIyaXuM2UzOouZa9keeohiSo2YOIo+lS6ZXshMOhIHSwFjbdX
AzZuOhRLB4hnVP0PSEiSEHIj5nHDLjye5/EUIG6mB8rBHNjqdsBAbS8+sGodzftPnJCGzbbsRpiT
D0fdoueQ85mf8EY8gAHDkSkm9smjtsIBlvZaL/Bf0rgza2298uhkSh9JpGPW1PMhWTyh8E31KvCh
9TgfVQcuVp2Q8l4omOthJA8DlLALfci3odSKhceWMNon37PDczBdBer0/uTLzWSpUSkmzB4CPz81
2FepmlS4PA/lnGnC/qbAbkV5yXSDCy4LwuiD03ZHNbf7YbqMmO2+ERItvefb98hwR6KbT0CUo2FY
J8u+A+Mhu60iob2ebRuiMlTONG+lDp/iBtT5exzHj3kLZpJD2d8jom750n/gwVDm1I0tZUReICzv
B/RtBxLiwpWRNPipcIyWBg2kfzKe8bEg1lq9utW4wZIuJ/N7QFJWt2yub7OkyS06HTb8QxiTy9qe
bDjG8LNj3RhMHGkg++xT5MZOGMWK7OXTHcXJmZm3O9RjTMU6ZLvNNbpC/Q3VIbUZtF6D0HO+FeON
PSc159So8asB0WdeoE12aKLqHVkTlEeLG665CnIQ7wSpkHXy/pH5z2pQcbC6Fs0UG7SIqo1swZr2
voteIC6oPLtNZw4fajlNndMi8anonS4l7LpuxUup30UMaITEi1uhVBcgfggQD4mYO9CD1vTpNrGw
EsXeGezvA64L2Dw9i/elcheU+RY2W77uzA4cc++y4QDcVpH8HEC6rgnMkmqMAQ1aIiLdszSGGvoO
6T0QlS2HqktLd/ttRGl6Z96Rc+w/LEGRzvmXJP9mgk2bUoW9jvrLIr2EbFxlA2Jq27O6eXGkneSG
tMhy3STpeAmYXEkRmIh9weHyV7+r5MfqiUlELfwoLgIiGMYaDcRsN1oKDYhlBsDctLIUyNfEGnKM
YBOw3osDBwtOzrc52ruIiz9i26Mwb354v3QDCnD9F0ePkuLiLxx1b31t8FyyG9dPZz59bVBVeOcf
oKqQtA1FYEe6AhRGweNLQMg9kgHZZ5fGZRDQBwX4vXkTpzW7en0CP01ES/NVwnoCVTuvXDLEZ6I4
MYaH9PyuzylwKqkKml75T70pVl/S3qeaMQk0O9rvUrYDJ0IDMog64SJreWSPi9s+ay+1nO4d3Vdm
RQ/06pr/8sYrbj6QYoyY7ntSkDcnoJqtPerI9I+xc0KJS9aCcEyXnfpRAy9qZboZ6tgM7gV5M6D5
HpWF/GLRZTr0pp0QH50TisdGmnWG0PnI78QvZHDgDX5q9RzEJsYSR25LkmkxI5vBOc8eLaVx3TRA
5pEUPhP3T3T/TYlSBqXgQCSilBNmpXgFSC2vqaIYkU1476K8PEPPA5r7XJOT8C3IsZEDqXM9hUnb
LPgtPPXGWHL+Z/ysKoPNi8AaJ9kuAFM++IaICq1QJySiCNCeM0LE1DhviVBem4Tn7mVSSkS9/WsA
cIRP6Gf7m9Nq7BDwuak8iL7PIiGJ0xxF9qCGgz6UOLfEpKbV5O2gwImLi13Zh0Arj7w8ZGDdMQU2
2N40d9xAY6tW0h+R3qDlaCMDBgbHHDt36Ws4On5fB75hYd+B1NUzrgytZ2GDQUFQvKOo/bW2M9YZ
zfS3oLkWtxdvV08+RbnZhT6O3eBjt6lrptmcjQHUDOSNw9KcIdpRn6+b/cjZKEdWGyo1JzSOdbvU
BQDMsf4XduI4/JzGwoq3SMmKJSQajCen0voSB//sur62P6eGXkWJUd3IFqxxNcU+uBiK1/6BmK77
x6uglOFqSiLt0EE1gnR2iYDhLykVI/yaEh8vMSng67vs3Nb6/U0ToUZ2InY5/6BM2F9CKc4i7osb
1dkmks5gLCZKFPhPTtlXw33vVHvvp4msddfnMezc7CUy6+Rq62qS06O09td54MhuxIVYITkYlWfX
kTg9BLosEFG0WpLJPyZ7HmEqcpZx+Q7iO+fOaavaHQqfiDrd4MlQy5R4zYYeN4N2OE6nDXWii+EO
gYUbZZZk7KP24vSY1IfDBcgv9g+jHWlUCiTfyUa2B97a7Vdji9DGhtzAOsgK802DXNdxvyb7btmN
qoItL+guI9lQZJSeHpRZsxYR2Ki9Pkrpnf3znVro7T5VxWS1p8Q5hOwIXoBKTeregKHdVP9GP71J
ukLR0k9hLYnkCUq1wYnbMg+q9QkBB337y92ORG78dGNg741mcjqQxQIRYSZMD108Ed4l2/uDAReb
J68IwVBUJilJeCabDPWEIvmKJbMlhXiScoDTVFp5c8HfokPK9gorPii9CxcDa0wY2XlkqrkbDUTu
LCRwoMj5q3/Ter7w5xWG+iCgf+9H/v1ux7h+MyDQz1ZtDBO+IFv0VHSIjBiIZti/E7hJsgNJ+y25
uJbVMWv75j/w2zwp5IlZSIp1mSWh6HQHSeoj6N969JoodRd3Aeh9kWl6RmjmNlTiD2B21rqx3pG2
fKmyqVpWVauEpNrUU+5cPoep09k6+maNwobQX5vH/TQrL5gHCUlmS0famHso545jRI0fV95PMbnk
M2itS5pW0nZ2ji6nC2u7BsKsMFnRR5mTvDyTh4FcN6HK2ADSvKCNF4yVw82d5+B9/e4xM5wS/CSG
a5RCuzNHTlIGpik6gWNMhCfr21qCb6fKAItR1RZtLpIceuSPcM0gtQJeXdAn+QK2zudoCFwxa/MI
mPu4ZuuCGMjt77Szf2K41nwPD5thP5gjOC1IQeZpI9u8XADEvR6ekgjj+enApQFp6+ajcs/QQMPm
EPRGHpu0kp5v2o7tAM0ViKYXV8+mXn917AFGtxcf449bUcRwfxVfa3XesRefqIFLdyppaZpuBdoH
HGt8Z6mB2ggiNpUYdKKFllzULXYtaMa2xRKW/rMvw4cs2Qk8Q4ol8Kq4Uz7c0jtYXsEMH2JT+TTC
oDWtO/ptpKbAOf5FKtAGW5tIUXKEOWBEOp3RnBQVgQaRODVetNtDb15ggtG+zCeBfGFOTNnM79wY
//mrQ3sLRqpOYn8YlDXMYeB73WvbhKapUzYc8J23MUwT9gHiuOPWgwQMxq+cf7M7SQFhMM/27jAU
5ubTgCmioqHhJc+Lc4PAQivEmEkEW1nafnFZu6dPUYpWUWHn/FoQlM64QCFekDRkdh2OikXsh8BU
aJg/pJQY2rjHEcCUifqHn+gqY2w+IX19FHgwLHO7ovSndDBovW6oKCJey2thjAS1115fdgSXFvzO
0zUcTa2B4QJ5OMyFGMooTB5ABCL9wRqPX+03y5+RHQZD1XbX4e584OeIXF45ec+JxXeV6h6vSyd/
T4GKmekoD53+GXy+qJsq9GoG4aiEb2IZdrBgMvY5aAa+ng+AF+UqOFEpRoHNlU38pqXfmT0/orW6
c3JasTU7M9Pi9PmpAZFJFKrj0nEiUwLPXjx3hYJj9gVc9Ei4ldBY6+XM90WkMH/lqb3mLIHZ9adb
m4IfQICD6D3kBP1KW7fY6d51IIHNtShAdcRAy8/xFj7R9aIm8OJCBNcOjrFJUxpaa6y3v285Fbu8
qou38kR3zafsdmuXt7WBMLr1e7+dNU58VU0LHYkfJcj2DkngPZPqK/OOUt6QEFvd4rNRbEHvSYOF
A+OxCrVMAXvDzjiJYR13EiO8Fv/r3VYYfg/7tj/xnze1G6p3SzqA/H3xsi4dxSA9Jjs33Im/AEI6
4rTNqF/Ty/2lbC3jRzSD2I7QAA4ZWBNxMbQNRaHPxrPnrqRbYIJSJjX5m0/rzqXuUH2Yau0VFdeZ
yWSILkcsQrfRHYih7mBK9UjkrDpVnUmhshh9aB0CW4vfPFTTznrH/zMgefJfAXU/Pi1YqZiYcITb
gXRHuT5364XBf4+J1xjkXmtmqa/3ojCxD9/Fj/g9xjaE7pU9IruNIqrKTAoqFKALHUXSD18YZTM3
UHt9/0Ju4UWJVR//6Bx95xM41nUnuKsglLLwMgqUD83EuPDAihrm7bOgYZIowGbNGl6iDfED+oGD
3EZZ1X6tB3Rfk230ktDp0ohyrCzwCDMwXmlbHTEcyKxuDi4MHSa+f/qBJq0QZXOD6/5X/ybZZbQr
ZjNwn/Ntwo55BNr8lzny5mulKhTa938jxNbh/NNq/GrBBvgHvTMiLdZIcC0yn5+fbVAqljyII8xP
bPH8aWHqWqjemnFdPse4rhv4nrUz06BVTvAyq5p+PXmNDPJZl/6nOE67IMldsdpn11CerM7EIu2h
cUzIBKCvtiLXqPCIKDxUD5Uu+aw/pBdscBjQRvJ9riKsRmAbCoAseiMIt16X2unPQ6ILjgheMA8e
a4GhQTJ3mhTY0pZF/yZwdEDL2M3OpsikZudbIRaFy2oDiF0O23PbpDcUnmQ6B3KRfqHcaMporxuD
PB/PQWrAXucLGkP0ASsgrH/EbNdtauoVPOgAeodLcVoQ96sRnL9mHxhIxLBrFQR1nzEcnlZd2N8c
UpUoRPULJXOPGCGjNDNQPgcxixiBCT6w7K/oMIY4lAJNhPW8nTPWJXUvUS6uAxmJ05CeeUevJ6/o
eLl0nNfTrmIk2ldCjAh4as+cLn1FYZWOq9yi1YmR/13Dsb1eMbzIn4l4iZ/N1SIdAVUtWi8ey7pp
UvyBZdE2SRFdmwQcZo79P4iY2cSeO3kJuBqAaesdRL3sbYAeeWrBulzt5D/VhFNvYp4pslyId+z1
Gn422gB35DD+1RBsaB6cptwwO+9kCyOQeGs3j0GoGuA7wFd+GxQzD6SYqbKhNjpF3cM96T1/9XsJ
Su9X9Lf0MsRR9rmCdmbQ27s51J1B32pf0mY3G8CBx0bmPFXlqGwn1cULU34RvCJbQ/NBWW5qxtku
Q5n9TMmRCG12l1Ny7oXkEzoCDPL9If4eM4X/OcZttwnIbUYOSQtgYg/ljVgeEGlbLlj64aSYztiY
EAEDNtSf8SR88WR61pIHiVKrC6ZjLlbntItAyAqo8d2a0ES61rAXCM4gfk++IEwXkabzci6EA+ue
xQ79irCp9vgqahTk+HusiLVLeIYLVFogua9JVtirxE/TX4rdAHy94e3yDapaVTtIz06MslSKbD/u
DwmQeXuKNrILUitE7s9hAweQ1Ix4pNQoy/oijpZaTs3R4+qTEPCoSj4tCBQuGlhXHTsgEKNDKCkW
lz3i8YAC5hGa3XI6+yuNWEK5sXkRw41XiPKWNTkvvER0k+l0hN1/KnU5QHX9zl6QHYOIMXnvSrcD
bg7xhT1Xxx10KMT06Ak3OYjdyBwx3LGfME5yS+ODzeTBsXsRslwFZCqG6ExOO02MlFtOvjekHT1S
n7kEk2x0I+616fxcNVqTSmGPELq85+MyfzFG4LCeiMRSTZAguHIUDgq1PTx1YK2MC7Rd0fX9iqsW
5OyP/4tgC5NY8qtySycxodKJpsE5jB2vBovaDTvT5aM0HyHFKzaXdWy+EZSBKTZwmgwQavb+vUQK
uj8BWPVl40jPpFfIzNkyx3ynUo15ER56NBzsriJ72I2b8Yp31NSyz3xllN6Jb55j17hFQZSoEl1E
fkmkbHy8rqqgHREPjCTPuzfkE3ZKDkGlUuwEgRhcAED97+CUEYB1bIKDwFt2VWlMYgKcdVTgqZ0h
5nTBcJ6aevTCYZctqrMIW4z/CmlbCuRcVA0GYQLrhSwJ9wA9nPBzVsI4PSCzWy6wKu6XpK6lfOSW
lVR+qmXg6aRW8gVzpJZyV35fe/eX5LNhtKQ8GPji5R3EuY5CQjjuU8H768lkPgmviAUdOXGWgQn0
v6hxNT/7fyKAwQB3wCCjMP88sOAwbqNsnxT0Z/zk9CzPGgx9UdY56KJHyQQoPbY+gvjnlUc86z5D
uxLddpmu2oxquNjFQLru6m4MB0NMah9AmgFQOMQ6J5nI0KYoqzXM7OMLui1AYQP8NTCnOKnJfs6Z
DStMmgiTMP6LjXRzCHIv0b2cAYv9odqo3/zPHKVIP/ZVKK7YJP4Wy9GvOu1MoO/AlU/tvKTeCqUD
GGz9yxve38rOUGHYdUAh86kHbpLn1l0xaw+Ni38lyZa3bpXiNnvAeKCvysI+3kwFWpDehpPtY0Kz
q6M5zdaRsfxEIN7/anghgeCWiv0o065jj48XLZxU8t7ABQQ2SVkoXyahLUSOdTm8B8dHiIa5Xi9R
D9sSBQxq/evyEgKDf3IHj0ndmFXZUiH95guqOG5+Ms6zd9byNiCRGyD78jr/ncdNqTWx9cNkvjwS
OkRSoPU5FgyhHasJJeso/Lk5RYR6ZsfshmgFT5cJgWZaig4rG/cMnRLTcJzfceLtf1RCIvKAMPjk
Kr/xqyYv9O5vSB8xWGQukmzxu+3xx8Z9N+u99tkFcnZkYOiap0s9h4OeeYMxnPHuT0CTyl1oeyWs
9trRpvLb5XleN+OUxwgr1Dg7U0VkypjJHYdX7WiMy+qKlDyWRSPzLKT5GRp+hdmjnvto6TfK9ETj
SN6bFOA9HvtdJNwb5JFMYoJK57a4uo9fOi+4JCs/sU3DWLKsF0d6BiVu/DJsGAxjdF5Hxnsu5s+F
GEYiBBH8Jw4839W8UK2kfaCmiMIicZYPmN12MYUAtiRhWpTs07ilSTFSgvYyC+7W7oNZUb2qvc5w
TXJtzMYGkfZ0TOrpIpDCXFh4FSDBZM6AQ1Ohk+upsj5vlg36M+3TR3ryxI387t8rBnDN3bHw8FJ/
HJZ4qx2lHfbYLsT7sYaUCt2oYjMArtWN/lI/Hm6QSg8s+I9OjZD14qv9LIK2wsPzB1QqfbOvPXaJ
M7Of+v2rbB8Sj/IASE95XLo8e+90rzeVx+p8s33wI6AQQ2nMm/bLvdliaA3k6UvxPRR48UdR1p6h
+WSg14EWQ+e3DwoDcmzBt45IiShjzX8/BMCQT2T+bIBgz7GKFGmEOvRhzt/Q1+3TwOFAmvZFfsgz
mq/i6rm/CvXVHGO9QhdEaSAxEQs13Omo1JRk21043iWN6U9/F3aCbZ2+eTdQZjK37NamyW9et2o0
AAOOoLETplJyylIoJeIKMao+9NbFxv3aIXOyqC5OrZeP/eyYx2ax6oZun5OmwaGmzvbj/8iXNTWM
2kSgJ2yRIxQOzm1K+zNlpSC09+6rGkBx33MaR0wbLiRwTMc+QBbGWVj6Vb5GgSdcZn4RPJniGLid
ctUt8IPb1t5yUfLlfxea7i/KLfMAPNqjKF7qIHCg+EcwLJN4EkvCWgPOC5mVy6ijI9wEyYviZnF6
U6fULrCBl+Rw1wiDozOqA7hmrK7FXPNUYzFaDp3COzk304tfC+UEZoCcNaIMQPjGMxXbZQswZufn
+DK9hJp+RV3oPml65LO9qCOoddmfZpj/FPiyoZG215UOgN6CicsFQ5yVkbAcl17UjTUkxclpbyw6
yQxZj2KBQaNxMCyKXylhWn8smX+CVNFZh1jt/JZ5HULfOGgWwH9OaBX11fgWPVmkUbvIh8IROyP1
HkCrBVLAHkLyBz/UhWOU02lklk0iZ0qTVRE9UBudXLUgR1W/9ZLnmcsYk7IJeXhREygjn3baBGIN
PfB8IQpuE1P01a8wMnIlhvKWfmVLrztFNPwXqFhtO97o+ULf0zmDgCKwGTaThr64ABnL6z4t4mKd
RGdXWwq6I/dAR5W3F3thQC/bb84TqOUBIpgF2Civdh1EJn3YR0xdyFH95UT1w9DnVuGDZA9gLBzn
qK5RRM0O/t75WmUOrRYPvpKJjzj5b1MaN/u0ZRiDFc/x0mT5vfOBC8gssAKo4Ru59mbse+jvmMJc
hdwraFE+wx81PknsX/govFMh02qRnWlEPmaEcSNN2F0s0NcZfh5975yOkMFsevNDglM2TSCbTQGq
408dLS9nzoKF9HSaW5isrbcDAhlWYN48OpiAfcO0EjhXQQd6KD3Y7phA+hkGZ03UcNilfASW2fuc
UnsBGwgaM8ch8MPWHmT5PK04evUwPnpEki83lFoG2252ZEDATcUPhYB+R5ZFr4+/xEOr/z11RlnP
kJJ1QQMx2rLWYo029KviR0y+A6ys36i7+iScjM85jqbtZEtvSoZM29hcsiQcYjO7BJ5zeTFfh1qC
cgFWdR6k0+BfE21KNgXt3tT8N3Gv45x3K/hMYA6FAjqGOYG8vOix80ZjSIeqLd8Lf9ZS8FmMKlxC
QtVwa6ESbZinAH298XKQ/3H9JZQf3dYxr3SEfDvImMtjbGvknGWS0bOQubHIm2WdBBjTaO+PYdas
ciXkR7Cxs8DTwb4b7SlOPF/vxv4MS0UGhjimaibGEvpqNWci6excLJKsvh79HktlCKdWkNTFvzrF
qBPIm+KhgrwodZWUcqWB7leaizZbP6k+wYtByuXB9TLjDvyaSmH+I3fH1gDFtFLV5XFeDQIziow4
DGIuooQGWOHwTH2shqdyeWHvjX+dpItfdjFbH0YM7Y1hDT7X5C/ZoIRzTne2leh3UTsMPngeQLpq
CD1QSdI6XCBDaNpMnZ2+P/S408K+7atgA8y6Fl6L/PIhQ7Ff1/COOSc6YcL9fhUTNDbPDCmguiNb
mOLt+1NSqoj42ZB0Mz8EvkXrpbZL4bqQGyP9qiWIALAFltQlPfIM4KseQAn7gr96R8IgWqybpgI1
Y6WAfp0YV5CxDJrcOL2bQNmVNvfQbB6LWxOqF1jEpH2gWQ3oavSnjFqXucj6apSCYzkBJ31aOn7d
0HIEOTWZwTds97nnC1WzUpc8mcnaY10QX+BLst1ztWh44gt8Gxw5O9oJcn4lGjeGyEUibFYp8dFr
1b7poQjVeUsfW4i1Utk5dqvkVYxY64WAwTOs5va1TNeCS7290Lb0pFItj5gL0KwtyrKi31Oy+YGD
V66348Ip487GwvaGoSL+lBm8wShti/iS4gdod2FmMbFAx6laY/2xedSBDRse2hAd4oNkmEo9MJ86
v1LLx9zUExfZceNHHkilwBTIXTBnreL5fHEkR9y8TTEi1AENgY7BkBAOMt0Eme+uUyDAOGYP7oLP
KnFo4cFYTk4oMXoEtVtWJyOHpfVJrBaj7sLSRltitiDvoxfCvW9mk7wDvahQB2eVrsrVVwsI9sX/
2yrOZ8lUlNoJBJrvJgMO8N1dv01PNNlFa0TsU7+Simik/NOASM9QBhueFgedYKhCyP2xGr3A+rac
x2sDejiZzmu2FfI77kkjmRwe0WI2v57qn9BeObK8tQE4iZBMysKj2EkS0rNJHxCDV9Nz6ly/ca0f
29SUnTAiZIqxxDhg1Sf45WA6F5ZG5oadzqgIrMMLq1gXD8juRBV4QysaUYlVRr4b9mu8GD8Mt1yS
b+2JsD2fFcpzw3VJ7FzWx2iDNCFahQMThLUhLusM1+HkXulKsr75/RnhpI/MO0bePoNZ4t437Edh
/aqcGIC+wm0dEDgnbho4uxS6nNFthZJ0epWywpZ6Duqk/3TZlW5KuUwrIRKVfMKcR9SGpH8etPrX
XDrCLjqUGqiKNWRw2PGpEKV5hQnBzyyJYZTWvE5snk2c9y0rJeoLeeA2pf2kjIgZJqnb5j4xyF9a
in8ukP93ckn8mLzjIb7L2S5Un1fIYDWubbJ3Osxys36Ze3yT/sbXr0fvmLX/HK6JLOfBbZtTImBm
9DZB8IqJUxgRBN2/IjkW1Vfe4vwLi2uj0x7H7bijPKne5tuBPpZ7hjuKw9Bz5oEUMIa6tF9IFkRY
pRk3Ehk8glZ4Rxq1IFyOb3IyvtheyFuhBRpRL4X2zSUNo7kZ/z8ymxYm34KL8Vfj6vrHHW2PsuLj
MgIRplH3Dhs+l232yaxNt+wgn1LSs01EmE1b3Zj8WxAuosEPwmnBiOPNXpf4uj08Qf6wVhgqn08A
BFI23fO5nxYMYD+0qqck/XjaLQlFgG7tcYKeFpJXF4hWdUYvskX64MOzysZMp0zf/8N+eLAlQXyq
D4pgiMQq3hopS4GSxZvCcUHeNyZWc0qbTirhbpgNpRVUo+1nYu45qhSaKf277LdGw0Q72YE21HE6
6SnnAY2byWBrODmJlEo5qRQtay5qgqyStA9ekShCkK2tqRNCs1nzydT2StQesLi6MAWRxVA/Z2fv
05zWBHyhzO0YHVHl2H91W1SCMYIZTYJDqAB9A8YUc0bGL39vjcyWI/5P0QI+lh+WSwsjrxOO5Qqt
nga/ArabHvB7U/nJ7k+t4T5G+Q1KULo4nIRTG0o+C1NH9rqTJGG8M99on4Qt4SLu4AvAAALdo1q2
JYL4C9HrH0DddeqgfMQWlKbSHGudCc4P5c8Op/dmTSet4/eVm721wTL0V8LURX1FpqpQOJgHzDJz
IB1Und2YtVcbQRVSNp9Lv2iY03lwATqIn0cvHHRYmdzbP6cM8c/ZghRdNEa7aKuj3ln9p6BiRTRZ
VUS92TQrLjXbx9EpsKYXfrQtH1e0gwA6ruUJozXITJXc8/grUrwxPdVS0CZD6Y7J3Orj9qay9XpC
CfpCyJAuSJgjZe+BnyijS5IdEzvZ+z4BkIZN5EFtZpiBj1qAE8CpGQsheoo6X32cb2HyGSLS3qGQ
2laoqstFaSwNXX8yR5CEyZzQGCSCJCfh3aGtOs3XRq0Q+3LQOOFu+4+yVxjypTifVtW4C151f/iM
BDhCJDgxWtIu3B8IpcUIDrOz+NpsM76vGNDCiymdxxHGSUEr6jHa/cvU1mQ6n9hnLShVfUglt1U1
CEaQnZJi7aph+mhhqaV0o7zPIc01/pkqmNdaS6IPucbViXLjKDnPCxHk3Nm2ZZzHcrh+lg7v17A0
/Q8u0LnLNhX2V8xmIHykbPlJa45CqkE5fRnLNnaR+lPWM7GeGKpism80HOTc5feSv8tIg8FRzAwc
Eq620ummlPCujAIaNMngDIUm4AlmEyfs0Yq5LbT8ueIDPHAZreO7MnKZgklHM7nbofLmN70C+wQV
odbvi2PcbwvpmIqJ1hll2V3DupVYLm+9vnqzZBmk/TW9eG1KY1CvOWaBSBKNdWdEMibm2QMVfwxB
yz9PLh3t1wFrkGA+jfFDEXqJP5tgo2KSLxpN3V8SK5Bj6kH4rO8fm9FcBjCOvRYkKMbbGopmJQ+3
o1v/58ecUQvX/4HrNWsDHNY5ZBfNUpm9nXbh4yJ9ypgoXWh81uNSBS4wJx8KQgdvABJRCXCOAYps
xZwit3GohIjhmgAGm1I7dB6GxXi3DDL7cEL9claEt6BVmVm95SRRH/2V3pTuuVK7oyVhQ2ntXBz9
NixzPRA91vl+IL2d+ddpKjp/2/+YaBKr6JqrDnSvEm5FWqp2rXAw9Agcxz7+f/w0duJnUGHhIRaU
fqA7m8vlgy8V/xVMhm8Gh2mgHJ48xd/jlHpTeSAQQOcmq5dg2IlqDqGu2pfoPctiyE/ushSFlEcS
WysPXIJujcrA4jWMG03sCzBiBFAqbTW1tSp8KiXcLPoqNRn91HIwXiBuV31AKhIVLY5veZheWVU/
towt+b8f8ygKwsFSt7e85LIw32WAKZYQsqa07C+NaeXqbc/6rHcj8jUbg3dte0XXcTS9i/SEyzEz
4MdKOPEhtswmM6ypvFLL/cRpK6Eh+FGbdDsUTytKiA3z8kxL435sVxWhE9YEhANfCqFDsqt1qWU1
79Kx/qPBrRJ16iMQJWDqIbLA6/iLwoLNJRp5QwfD+5AwvqWhSGF7fjoZ6MV9aJN89gns9lmcU+ky
fvs9iEI1iisaTCGV4XLOYBbDzuta/jnRUbG54naMprM9yCFJHdNNbgHctxecepff8BgRrwMV/K5W
Gb0N4pqc35CrK56KZn/HjIcHfdnsEcuNOdOH2hEPUCszgimiqtKUXmSA1xbYlk3dN8kURuMYosWw
ZBfdyaKCqp/MJVbtQnheSxx2sOchPhlLGHWNt4OIsdw+c0JJlXnMlwQY/JEzuw11yke666sVL3id
5bhGbuOhCwa2ibBWuGP3L6Mnpk/3Vru0MLom5amcz8ji/jaCGmuvVL8qqu9ZtMjqqG2/LO0RgYXT
vawTiLhzGlzYy6s/E0q53pNDLDcq9CJmxe6UmGySXx6HVXJ9kXBUecCI9yeUG5hCKowox5Q0J/i5
uGyaWHkpslGdx2JcWhbiDGY1M7PP+yt/LmoNRbroM+zuQ9KngnC8w/csEgpdBAx4EmZA8ATzGgY5
ddRVJ2Vz9LfNlNTU/bm+ao5oZHUSGYT4vtZqWYjNF8eggWcNxxZ+RTV/k95X/VSRSOmEkzDiWb4t
/Kh03UlzIQFWkW57s+/XCgFUe8WsC1GgRstjMROcncz3P6mkHZAdoJBlbFioAxMW+XxpxcZOKmtN
y8zZcmcyZvNYD4f2IWn2Gnr340BLqj4XPJxQv1AGUP4Ui5J+7b/IDJ4iPVB38xZMLiGFiDgIkJy5
Kz1Uq3uHPXXvmKki6dNOvyqtCpOy8R7LOtz6MGm8Ai5ZGTgBlpJZsy8aYLi841WB2jw4PlNeXtoy
h3gr499wnIyjd/LlJ58MuDuuG7w1Py1vJ7dFwgNmoniWSq8dEx77G2Gu7+RMvxBQyZu790ucuFnc
HZKV7hg//ub7R9oAjjyI+cYe5q+7dIvteOd8O8sWCIO0/U0H3GRtx33nadB+5l9a7HQT1U1xBlUP
jTLHFirrgqcgjeQyRhNhJPlAbV+Atj6hYbslf20s2SlAQmcvjb7XpG92R/TB46A1qyAEmfMFgS2s
2p+STeKmAft3DfugldTFrQYr5zoNeGHi979a0hlJ1zRxczrZ33JPsupcBp06HQ7NcbPFthdvh2GR
R3eVslrJfPozER2LcWgx8I5q8APwZY2DhznKHI7ZpIG8r0Vy1boQbCCiUap8FszNhf9BFn2ZUdRB
QKaL3tAc58DBw7w40I2ovQTHeC02zJqBJjw8AjljE65d8OVZo3bTG0W82/eHxqnS6a0QhCen6QVC
jyM13oGbC9Y/EjUpJIcCikQB2tjPNpqk5gmzW2mBh4eBrDv0bfAeujA7EAI3dUBqlz4sUNQ3wllx
PJUQC5WkEmEQuhAKtEnhbZ/O0khs/1pnbCptq3nwRP9yBsNWxk1HSi0VYGa/eMdKmnqgrmjyGt+c
Dgf6fK88AEBOaVB+xGntQT6b3Qiqx9Ad93bWwZFFYwVTnx6qGYLt1P4ELoFksibkto3///3Ek5wG
ujl8Qk2QLYg43GZaYqWiZ7abiTYY7EWNW8kyKBSMJ7p0pN0qyFChykhT+AgYbqrNJ39bIeeYRlxr
MReT5r18pQcmF70nI9L+31yLD++XB0Oc1W+s2zmBltkmIYnyvj6EmyUEWA5oZ1LnskZxJMMf4ISi
GFRJtDyQ9bdRBICb/WbQg41anawh/HMa2qWqrLOKY3DsZNJiu1xGYCJqiu5wV6F1ds3SKZgBGHVR
zFyqhZiUCd6rvtX30O3tD23z/heBolqWx5HlLiT4Az7OPgwRmY7kiA3WP+o5WDq9CUgGmGoN2Crw
F0ClJmHnbO1DVt7lnr9X7CsVQLnylF9hfaJNdvZB42XqF0pvjfRX3l7jPtr1A5mShsmsBLoTWlmD
UrzNDlG5FXD2Ke1Rnx89Y/70q8oUj8hV42ivl9EhVGu+EMl6h9G/O7ehIEMMmcxlnbY8u67kFaUQ
IZoSZoAc4y01Clyq4mLECAPOQJuPyHJ9Ca+6PkdGGb9TQYwEZcmiz/Jk1FyrP59Q80sl71eCUbRp
uLLqDN3m87uBvCfwWhbMozoTsEi9TLnLf3KiF1sTL4zoD3ZNUDMcfptRq2TwHLZ+neGDiInb0URg
+GKsS8B+xx0lQtt9hTdmcR3DJe0i30/WwnqW+0CW4UoM9Yxey+wuSS6pvbp0b/fAWZaLrUMp5utV
v0wzDWCXbJiXsAGv+thcqBXoyDLhAzj7AgvC5N0NIlBOLRKyuiAmIV+ydpVVIr5HLnPyWzwuP2Vl
sAvekpzTdmslEJO3sOfv8BKAWHklQAOq4rC2X5LNefj8pqDSk79WA3MfDU74MQ+HzuFj+atDWapZ
mPBA9Eg2asT3pxiIjNOrM5U3KuvUVLkHTf2Q5dzaSme5h0IgVQaRJhNbX3YYnlOVuAZsQnViSiQr
4ydAXSLRCQWrG9nN5paQZPStWXZ7lmxR+h+UVtRjoSXZ1qJ96EG6IWHcWBMQsmK5Dw374n/KCza8
n3RMHwykUBAwzEaspOWPKVDd9klgV1lLYcFw9p4tEqI68zgloM+tkHmZGyArYGTV9ZMCG4ftkEIO
fFl0X2yfULoCoDdh8V0o/iVjQ4Is8fDsjdF9SqgOz9y08i6awIcaDtzc0z+WqHybnIZ7801pSj3D
4rVclfhUjvnhTNyJ7jHdRgFpPxWVE1erLdKDLd3wV/6FhjLSYBCfjKXEnZLMPFYvaGDTuzC/473I
/1Y4IxAG2aiCeX52SiuNwDitDUS6UuXVTPDLo6QRyhm/3EXOVElYYynHnBxXVa6Zr+U4TyQDXmbp
woed89eeBDMeTyWtALThH9JmFqtNDWugdmk1Glk73H78J0jIT64RIwm6GmkLyJGP6pjtclcC7Jz5
vZdwTyyJyE9Yhb/gvtesjfRb9dfW84QKFDJTny+Yz7lz8qOiWMXq19iKEOXkCnmxjsgfRdq4A+ZT
8GTqpI0OdGWsePpIQGIeawMYL1QDlK24FIGkoVjhyykC7pW65cop6g1Q+Sdbt+zVaCSq9bSpu3Rm
viMbnemaq3otPdJvGryDSC7XzisaHwheYC8IDBjiPNj7nqf+AD3A9jPqafnDNIvBoE+WgOvemEMk
X/NcfxIbLNdUOoLKUp0TIWY3QvLlrJeQrJpexURNow3AlT+nw43LHXNAtoQS5QzrIIMR5DTKRrKY
O/Bi1jTnaQCJBj/n1Jh62pfUCjLvWMcnO53QXYd6IeEnze3fN8vfaksof+FrsxTVss4fEpH5Z8Jn
yc6KT7d3jdOHJtyvTBRHME07JIBf0Ylf7dQ5P3NejWnAMxP5qfuvaJFDau5xrqdCtwSl5/e8kKZb
8P5YAk7Fm9ZnN4qRiVYsIxAvy6zhLpNDkruYjs/SZkbs6AXSjaaZXU0LGG7g7K+lW5twbFUD5CUF
HIdA0eQCBtagQtpzrNh4zu2nylbaaZkzb+vD03rIyWu2Jezhk+ntZZ7+G6B2Zq2a4LTozJS4gEU/
fHejhfMPmHYBEnqHz1rFD8iYWesqoXboHui3k2OxBMXUwhWw2UVhojuTpqO3o7Zz2gr7Ek8gKYsg
kiKEMV6298VI1aatX2W+nxjpvEA0OwRR+jMlb84OWP0YtY/LvFwD9sBnNl62+P/W3MC5gdJosZYh
M1/hgTXsiAJq0To4jQqnZWGXMvfACNEIFcUVp8JNuN0mfNsuo9ZrvY0oKfbzcIEP5ZQ/tR+8BSQm
oi7bySgYF0yzzjGGCXzjYmwLAXzGx9DuxyRrOiDEV69CFxB+PasSxQSvYjr/RGMdeHeZ/S4298IG
UxnjGguLGauUhhvgcQp7Bc0NmWLbpcowqRe5L4adJRdYnPaG2nhTI+l9qRcXlRKGH8ClqkHprlxS
F5mAeXy5xc0PGSKsOIaPKnZgqvoLXTm+aQC4EiM0XT7opd23ec2+gg9Z9O7I2+nq4G5jbdMI+goB
8z8hqIl0bEWanbdEBI7MEpsKSxcb2T5AfOfGY1A0LT2KMt1vkgU8nltvgcLO8Znu8gxJRtmXq+N5
hIHorBhsffVD1XFtm2OJtKFIN0pcNsmzTv2tU4sHDcteEiftm6URqvn3xJ0hWtzde3WoB4C1Z/xM
uk9xAn6ZC0CVUcXhPELJ+dEddfPKRtomnUD7HOOnYalF4PK8XWpxwAMgBlU70Nqou/4yzxiMws43
Q/iithHJmAA8MZ22edOW8SZcg+I9bBQgp/Z5E26dBm1zW111x78NtDEjM1Vhle9/t1nekAE1MyPU
/yrm3H1kGhpDwRzAY5fJ8pCAeFiMBPT3HED+8WoH9s2yO/dDRZ+omSz7IJRM/qj3LaBR5la1m7+j
i6UaTK0KhlYN8XPk5XCSU9eY9B3RxrDUYMo3v44O3zAkzVIZ2ykst4nRxHL3kUUB3VJXCBU+64Kn
yJkIW5kcFq/8AzyUeQL8uMszHkmyFQWFKrW+lo1cJiX+FnAJbkh8q+XTXE3q7BI2k8xxUfMDHGcA
8hfXo1AsBU0OAelIPTMNKiWIIOQ2UqfrvW8CQmYrrAZm18WgBitkibZQjYFSwAg+KHj4MWnwn87B
EVzCxxxRHCT4+01TImrgam3ycDagyqilnWRkX9BRCwZ51fAbwMKMxqfOo6S5IWTb37o7JAGveQPB
blGQesju1Pz7pG0ujQNwpKBGsS0xfQt+JUWlItujo+it30Ke2omzIJ2b01TpboALjXFOdMC7+gyq
A01Q3PKA4XirjWYiClWOJpYCrUcCMORA9CAb/ZWDXeH2Oc47J8aQdvzKcUzhi0krTb8LEWhO/XpJ
cZczyVjrUcfbDHXSnNZZXrnujmRFCRmUdkhTd+eVy4CzlgbShL9JNcaXoQgA5VMEAWtDxkE2T/qH
j8b1YzhFkVXhpSjSijxwokAWCc7GGjyd9fIAyK9gCUG2/dUgS167CMoNo/eUOd7ygVviqdCa91fR
Al+NOz7epORW0wjFt0C0BuCYDPY9SADNjGVpI3CZwbVBHPHSi+WOjcfUpPEotPOEoeALHFw60WGx
PQimiiw4lEZxZx8NHujd5/Jfm5EkcUqQcLjeUYFQRhLgpJezJbpnJB9X++oaDrH6nxRjiJsSRddR
L3vk9xI+aJN5gEf8XT2Yg2dK/X+zkSaOeRDdlHfb9iIYbTU69PrXpt7d4XWT1vmjAQVTDaMUdTn7
k4c4xCYz1Ojvmi9w6kSlzf5CqLdZLh7eo3zbXKux6c37c1lsHS3olPV3a9yCnYAdyqkH5/q8Idwo
Xuvl0JEdNRWVFWJQk0iYUGfK+COorNEbm7Vf4spajxW2sENkx9b0LA7fBDhINvUGMvFMR/9jmD6u
gyX5jeEAEo6JDuhtCy4Kpr09K1IerCsp+V9Ti4jAqpODAxztfLr9UmzaxpDNctvsSGta5OqhF3u9
6nRXkabMCy5H5P4uRTdS4+NumL/DtTuUi1OBCTx/2EJYyhFMx2N4LZ1f58idODbUxsgJsgzv8h9f
lSMWld70mGQ+KsOBfmdau360KbnVb64Y2OYt5oekbM7Fq9m1+57FB8bLB71aJOGb9UsuNYAhjb2m
cEgZ6O8Zku5HMi6tpyy0ljfc6z50EST/IJGuX2WC/jJiz7o9X+pJ/+l3DpjNWk+zdqXPPHTNzvMz
yjxIQulC21gWWoZN69P3/RKNSL6EBPFK0z1jUHUPiwu4qCwHx+WfU7+ms25tIm7/oE/64jHpl4EC
eeZrdxk2/UJ5bZ/8H0ENL7S0QeC12ughpUJw4wgoncJ/22feR9bMGYjuwN5cyRzI8MlLsf62qN4k
6PHaKDD5o7dbDHhraUS5TPTQtDs/E0xJJpN4g0Yh/llR9Avd7z9cC86Gn7LveVZ5M8RNNe6A7lRH
Y9nCXri1f2c//K1JTcQKw+Jr5xfTbAbGpwGiJevyHa3nHQhtrq1YW8hsR8rHkZbh3XTRGb/O2sbG
OYtbbh5xwFi46P/7d5MFT3ks2FXGph0KFlUe0NUTaIJGvOeK51qOAuoBdHbCVBUpbZ35KV6w6r+Z
5YXgMqVpMM6MQmxa/6bEkXDUQ/IKy24EthT4fqYOTXDyZh4yjpgYnFnw6wc/klwOW3xi0M9TF8kp
e4EkTCENMYfPO08zB2NWER8yEc4HpRRE2svIyeEshTmVQtpVMZay05uYzE/tmZJT9pTWYgRDhP+2
R5rHXpjseT/f9/Jyv+7sRqIuBhPAdCY63vroNeYPBSfvvgMVNoi4S7GHDKra/Z+iK4zYJrIBFGFY
93Wtd5cDXG/KE++fDycnQwRjoLIy79erNmp5RvoLNf/QL8uCJAs994kHHHYHRVGSnQdV4OBnXM3X
P2sUtg6B+BPkpehTSP/mPw5xEQ4CuXaRmRz8x+TeTKyMM6e/xMAEJIkLxnl+sRAe27wndEXhVxMN
ZSI2N9/nBVrQQ3VuavHp1vdpR9DRsxWr4DxJp7vp2Po+6dnnYFsr/RyeplhR9mGMEeSVOAqFyNa1
bHPDhm+aaHBPUAAXVRtlLnpEydjhDmzYFZs1Ae3LymN9UfnOjZhDAV4eIjHxDlvgnjAFQpjVOkzS
ruUMAby2s2RtvPHYRRm8DyfxtgAlHo9mAOiqhH2/O2arTSwAFark9ZzV/3vbvDqweqLIcYYPXXIi
s/COMCbtPqC3N+I1KpV2PcakOT0lmPxfW868oMbLrNE8uue2vFFhlwQWvehri6RNTeCeGUDlFeIK
rMT5MkaSCfbKRiJIj8QxMKy6JSZxKJ0ICBU0TCUShggVd1kj9AQcydxHsdtR8bkImGBROBrnaKJH
0K9hTeooGnbL1OjTsPk5kRcZFYC3sXfITSrr+0Ph1pTLT2Nr8F22j8GxwRtBN4+Ryi7143Cod38k
kn/iZtIgx0UFa4B4ZN3/WeQBYy0uGU0BLxDN+cYrslens+gGNj6b9QEfzSRQ9Fv9JWJN96gGj6k2
ZcntSXLnT7VProM1nQew/c/hTVRVwZJV2wqJfY9++tYqqUIG8bz10pgbd5JJP8ZKLybDojx1cF8l
Lx30QlNi8eAzAa/weaihVUeKZemAamqZcA//UsKAzZXCINjmVbZsfbfSJlwReHzw/9kVmN7U9nZj
f4psKTmRZv+QDCqcBheD+Xrd+Ss2cLRNDNRZ1BLCY1Q4z9bkDzWlY5Z1D3IVNKyOA/DvatMZQVAc
GeLgAVKFtyUYxemxzonI8x5IcfwtAf32VxO8l/BfTxwFsqXIcSs8JMplnW4AI7kdJxIopqSWXmpK
pXtr4RgmjCeJUbQpzef7CIa0CZqbifIZ9QV6N1A0FpRIX+7V6JL8uuNF/9ixRjtCfspqL9VPoUtp
1+RpJQtF7B4U9/RO5xqFBdus/b70fJdYqwMX3EjR4qf1gIAKrF1PgE/IH3N1+n/KEbfZ1cm+xGCQ
3CPZv0gZG2ooRkjHlZq4RRxMinU+0MyENLtYFoknxrk0fcRfZaf/454mGp/rZTiTlzACqQT/eWqa
RcLEjjxAn6ozIXjG1c8bAgfUoHgKbk2R4oycTySO9SSclQT9LMy11484XtTFdj0GDzLs+1Rk0W2S
mRXCLinl+D1d9+H/JKW83xdjX0o77cDrv2n6igFtSIomWW0Qe4+qokL4newbGc1LuaZT2waKNrKf
A47whoB8g7FT8wKGTLFR+uyoZhH2l4OFPWGmdPErgB8fO+pe3A7tndTnYVI53vvM8WcBQX9UB3vg
Fe7p6VKtiCoKY+cHeobWTP7Gsmvu6xVupcPQ5RU0czEfjYSHh/WKzKTbs9g99peWtQpjbgfa1kb9
2vjeogF48yoHzCHPRgW39rFTjLEC7Egozn2+EHluTIJWkPq/217s8I0DOnrZwkR4Imf8pMDYNlg4
leJ0SR8YtLvX7CajTFXq3shIjzg2qsxGkRrIl8km7e2aWh1Ie1rZmQndLL2R0NcdLPI1ZcUJnWpR
IBsdFNnYZdzsFmjhdEXDhfo6Aerxze7Kaom/ixh++Th6NCQ9GtXaqJRD1vUsCEywsFJCznM/T3l4
Mvj2l9KaPJHu9zeIuamwp+DEu6pCQlq5EKGe2ohEhKUtYrFrRCO4wgbe4LttFEPF/x5gldSFhnWa
+QlIoUmLEymFzV5KCFXX5UZKdl1IasiItflRGpBLQLhc3qEauIQ11xT+NOZFDQCSTuzvC9FXt2zV
6GnVqlIFoDTYyDcBXjogJkwWINnoTV+tLKJi0Om+nU/aP2C6UCXQDR/cOhm1OEKVoWLtKvIyhz/g
6uBD0CNZ8X1nty6m46vCjFgMI60IS42LQXkN9AyqiHZ3Vw/rb+UYLw3tlut3dchdxFVwTZJc13mQ
tMFHgY0OJ+7XXHdXBflsONO71+KGY1WsmYM9cTtJRAmeuME2yFPoF0vsEQJp/CO/e7Mc435+oEU/
RirPPogiIfc+0uPsE81eiBLMEVwg0bNAwV2MA1mOlsG5hbCMJH9BG4pyEOlcwpwS/78Wt1a7zz8J
UMRd0aabG7TdPa8+ZHmheWbw62nWe5IxPYkkTNcqe2mobKCQUe38yTtyz0tOlK2zOMWBUEPs7tY9
aSYajOiVFdwv/JtZgcW39qbqRebZbFj1HB7XXoOnP5iZmlnkXJZJdS7Iemv3UF7G6l6ooNemGB5Z
2ouliBqSGd8wqPrr48GiLPHJ7MzWo2Ph5SW6rrjtYmRh0XF5r8iLerY7v+g9HhaNZhhtq92q7+9i
59pm6j0nODPywVThKHSzguZ4s+grOCYczodUIvgPyeDqidR7YpAY5XWqRpAP4jfe8jp+CxVQMM+6
KvH/X66pmVhtTcZ0DkuXp7bB+rSbEMtg+68k83UmLR8LG7tq6EHEsQIecUz7+cswcbZNkma3hXIq
WM1+GuPkGP48f6aReaNlgFv3GCsU+ZeBH/TI0ynNb5t9yUlWoVR+w1wwHAD8E5Ai0a1TUWMmaK31
D+aQV5il/pV4M+Bq6UNfI8ReCLzGfp8TOnKqQrNR+GkIn0z9fgAaDf8nOHYNqpSIvV2T+LyWLL1P
SBBFL2Wpktfw6EQvOOMtEutCRMQGxsCQfuSmqxtiqgMfhN7jGbHD+2p5zOfktWhcmJq4vBXHEzv9
W7/A1ja2xT37E+l6cr8/D0M5jS/n6Lo4PQbE9qMk9xT4bcNLVyxGjog6TEJf5ReQigas5LljMmw8
Sj0ARcQOz9L1us4HNol5ujhzboLgCr2Kia7Qp/dinpV+vBP0Q8FTbjuzvWX1chtn/mUZbXwBpLKS
VLdfoD3HDIgY5DNbqpiX5lRzQJK5OZDhlfdKJErOy2Tt7f2qIpoR96N3B39r7KiqzDvSkMJ9WKdk
IsC8uVnNoc7gJTs3a1XdrHXPpM+30MNT0inCYgkShH+FjuKO1zoR4BKt+9RYpbmqnO2/y47G43OR
EZAyQNGp9wKhpMvO0yNhLR5apCV35/XDv3UR3+gfe+uEGno9a1sdTVoN50+pP2CzFc75ajnhaYTz
lm5tNGaFyMPLJaJonh3j2NbwvRLb8i/IqSZ7E0qmnn7N1crhbN00VCpLru6vXb13jzYS/aQWvPWx
kW7K5dBZ2RAHBbnPi+TqOU2F/yv87bQMn/djndWyOt0lErkGKm6QJ58c7e6kIZwgkfz6BMQus94Z
UEAZxJ/3vHGGqhNayeyJcTlkKAE6HycoRyFPPzPdovheP1OTISml+q/VZVdD0ns65QQbeZz/cbZ0
qYPfrfPh2vzdiC8VPpY9AtjJoiuBQm0ecaz1ueY+UdrEYlkWo7Nmy9SrAKxXvtdRJNn8kh50/kMk
uDU5HmttGlyspXFI+MJI/jqHAh5dA7TiGfY/ALwWb9KWzvYsbeqHfpSeGKfveeuT0N3voNJVTeyL
EQbZcgqyoNJzTAVyiYVqQMnShlGLdDg73j91jbC3caOzvapsiFl0lINSg4GqaesZm7YXZq/lI/Uo
iExbdiaPP3eja4D3ow1jDUCvpjE0dManQLXRLS4YuIxI+JZeojEBajZvgzSnpDJdM5+br22Nvn5y
RbTF8lZCnJAhSDKpKe1GYCnkcXYTVLziMxa+JYBBHpMO+ib94BgMmlL+oH85HT4cdRynr52AVggP
8NOsxUrGT8IaU68D2cgkZIJtram0fC2tJPEVyi5KGxvkaDCu8SS+msGDh682XcOv36M0aBe3G6ha
F/MkQapbFLpAhSTscFkssW12mY5gu9amT9R/dUtb3hDUKrwf05EUoUUpC34Kkrf3XTIaKMRLs5ua
a19ZTv7fkuWgxmtWBGUbZpDCfSJiyFqdFkNTD5fkWHu++Bjoxi4YV/BqOsiQkUMJXdVqsSdVG30B
rN6wZfrGmACMiKdAtLru7jWPQnKjTsflqbQpKQ07gZBBl30f1qAUJYdud6hBjosaYbYUIC0vT8ps
bC9LlUdSX+6+hea576OOq0WB5JFFZYn928tIV94omMtORM5Eb6ch5GHp7BIaZgmuGJIlnzhzyjka
G7FyyKi9RvpXb7UvFwJFECDhnzhaGsn3DMkFEC0FbsfCDJpEYpC7ssGemsYhwiggfazCqiXGamtr
gmTMDHcrIHMu4g79qdhxC6tIh9br5qD+zND9cIjvj5UlDp9AOfp+WqTPZQnXEKfccYshQw4yoG3l
1vZRwYw4oyDib+S8eDxodcWBioNyUkUVbnNX3tFeal8FHjb0bXuJrlzjnpp4zflBuDqrfVsi8lcD
TXNYtxziPrHJyhsrpJARgVOd/ZZTox8CFF29/ki/y+1Iv874Kg7vHJAArqkv/AtEsJ2dqJZXYMEs
noy1zYW/Ufv6dMYabAdZST6mW1ZwnUiZeItWTqxcBovBsJOotXXZZdUqaur1yme3d9gj+q2XlV1o
nOgo8gDUFpklp1l7EWnirwbzkCTCa8zldZ0/pyhw+IDIXIzc3Irv/xBugw5ugGaE6EJuIzOGGW+o
CAA7w8/nig2FBU1gev4UauiqHzoH8c5t3/zz6sz/SqQjGvzA32oVQyleZi2tTRA0ioEDJsPKtaZz
HyZ/iUvkUG1eCkGCBe5j+wR8SwuuhjIzX814NZLwdnlAYlxvTeI2W9F6z8CXZ5h5FoKJ7+Dsp9Uy
oSTdSwI1Px97rWSgsonzyl6HH5rwBrMKB6N3DVRUFTpEM6DTfEhFBHObJn7DhY8+wzi8jHXTTFxe
mSe0mq7+e1RYclQvpOjG7R2ybqfJx3N5/iNFD5OGtbrd0r6xOlbwVbmtb1YaeLjO/EXmw96VK+yt
lXNOZOI9SM25kBBjF6uC6/L8SsKFGgROCISXAwWBC53wNNysdIiMVHMFIoy590DilIeZ1hPTneDK
N7JOtvNaZ2IYvmKypYStGknrPvL9jtKAYB1PGPYXYSe3q09NYlzZq7JIIA5lBDlpBn/QYTLdrmfP
6K5YCHJDyM2F1P7qUlIuVbtsKJ2aBabgmJ/VyIIYTJoQIBAeuXRvhRbiS8WHw1byPdv+8XidfNhj
x4PDi+Jj0xoAi1E4IFW2JHpBQNVY11JDrMeL7e846iCM+oXW5aNYAWcs4XaGXbNPg71aTxGGUmXE
XRH3z4kWLPaW5WDX+JgW4QfojDT6OMzZN3Tzpt6qwhkJuF3Ydh/XeZm3dvoWu1tgojwlAXHKQ/3N
HDCLp840tLlG/XU18qwOkWonc3TSid5TH4EsM9L9fjXSl8a1NykVFQdW2OQHCHzzz1cRSzbjvhUs
FJEqOuJwV5MelExNbv0xAZiI7Shk6Jo9zSaVB2T45E+w0FfWozrSadIq2/ECHia9hLrTDEGiM5Yg
RmfatB3XPfVmbIeRMiBrPpZFS37vYdAUqIiYEHc5gCnEwN//KZcFguwQybcwpWpz/RfWbxaaOiSf
2tllV80/vOm8qXLrpZ3iRSMEXCMZHxZ25qQMDpOsEyLisxClfIXBj2AGuw16YdU5w7Tm7Ad/XmPd
bjFWq71L1I5WFpVM5p4n/DR7EezY5FtG+WVC9bVW5MtN4g0NkLydyiYytX3ZEeXOiiOkzt1vLlR6
zy8D+eKK1VtTqkmlD/yR0LTTkFLrltsOnDNL9w4FtArcp1J6tvBaibe5dfZzWyQtmVmzjWUxf/HK
+bN77mwoTcvQ3IphILDrzYn91XpQe5PbHangBpd832IOaKfxZLB8WnTkTOnCLB+PY7lNikFZU75z
utVucpJIjCK8VOFMQDZkYSjNlConNQVQ+0WXvmGN9qQpJBXrIoE8lK2uLSjhCNK9tFF/IYLyZsW6
aLwkU5Lgd1XLRJ9c8xGa/nwD+gUve1jCnVBhWDjiznu6HGVzxG61n9g2B2fUimfevZafx2k+kG3p
GXG8/DEzer0PqPRrdao1ehV3AKesdCcfddnHq2T2Z3pL7XTt/8lLeqyt0yzwCvJVGQrQQxAbG8am
6xs+0XR2+LUDlE+pEGvryL28blY/dPMS71wllTENBxU90wmftkC//KFZXfFZvCq6XMm2PgIxeAic
UOTFtPGpx6hHfyojCEClbMJabfpR+BtjbzqFzjdbzKYxWnPrpt8qAFGIfK6blwGZLPHD+n5Xi2vh
BJAbh1itImYLpKRV+hxW7Bm+na617UBoP1tOI1+Cl3g7ePpYg28y7Rw8s6Uk7AVNgutbPJC4Xj91
n+XBixLhu0a2e7sSZgv9yYQYb7VrFILFY2WKRKMEkMX0xm9QMvFawQWyVNlOqiq4wZHiLEBDl+wY
1M59MYOhmn4QSDsv8V6eu8xSMtjK7GRNwUdCvm97J0T8dojR5swqlyCDyfA0IriVoL3Qj7sa3bZe
by1ibU9z1dETijpLjnxjds9SLxZphL3SRLFEht2g/xZafRwnO6l59LMf/cn7Y/Ptoqrs9M0LirBV
haVOS0k7wNO9YQKmK/AiH/K4aj+vVf4eR/hy9w7AA2zL6q5ee5Dw4xcYfC/IeN3q6o1ILJF4c6DM
Roj+2AFRfnFQtatz7ZnzaakRq7eGEBM4bszy2RMYqB/FuYnRVwY53y2ttN1XDBdHqoiR0y3c13oU
xBx4L/q51EwOMgXgBlwtiktVBZoXCqJC3ctPabcrtPASM2LCGmOXp082wSAnMQmPoW0+eW7Vg2eO
oDbuChDZF7EJLXMWKAkjBiCB12yL2abOVyDFvHWOxxlSIam5OLW6w0wTW//CmBV5t51UP6A7X/kl
WHK7rRqERm1thckPbkAEanJ0M515SvggESWnZB7f1smUOI+ddOhmYU1O1tCOz5ZFe3DPi5irC1U/
40OFoSlcmjIISNk4/LW06/pZgyPC/YeeY71f5egB4MHeX7Vw0QogMu2d3D1+qmQ58JBz9zvAxFmw
MLAbpetqd3ikTVPY9zaBdKiOg30gENSVxzuN2LcHitph0/mG3cDNjxIR49OWVALpWG3OaH33VCqB
ok8LtSIyipH3t2UwVVLbIoO5BIDEnR8gOkTfyRZmbTa9cCc7XJxxFySqRVngNKw9VVkT3i58xW0a
f2N4p2olB1OjEHcTHwkaCJAU4N7yNCd0Dkk3RCOJXJ3xNZ4hu0ZmIkw2QCpvnzn6uc8oXgSHXMxu
inXse3Xa31zQNVwylS/XRT2ZbdOnxfQlafrlFwldUvTLizZAVjr+88FS6C4QSenj3M6/NiqtU1qY
2Wa2ggi4QDf1RSauY9vQCbg0BY9vEU8VK7jyaTIXwvElfDtD7zNjKE0K+erEaEU0SQJe//b0rzwl
sgfx6iLmVOruXJv15tJJQtoK1+JPEdS7/12JHSmW+/c493jh/QLuBtzswhUP29q8ioR4Gwy5NEHe
oUkx3xV0Cz5mK0ABHrvu2vkWjPF9Sf9CFQcNqBabeUlaoMI+5AfTOQjM69/H6VStF5er9dhIQGgI
pPHtqC18KSHVnYAgGKPIyqNx5ZxAOFLUawFTAbCJkc+4Ww0jMhga0bnHoNpcB5HIyfuAsMWZ7/jC
OlgmZsFQXufHSTaW5CS9/S4xzEtE8S5LWFIzswHginm7BHOVZwD/Ztm/Bip6u7iwcsPsCqJWdg4x
gkj5XK2WdVDcQHjA/QaNOoSE6e1fC6rXinnMNgaCIwhzIHJcFhP5c6+a72Ivuot9J4WTIu49UmEY
MIcKcdbTKBx0EYhKxHGfa+E2K4jGXAVeo+bAKFdkqmk2gaRjAz4twlXCEK81urABUQ+oLO/20ppM
jxZnwScpEiki7vMNHLJOzH/77q2UJMBexXnj/KDfJvVey/FeioMBV4qdxvTFz0cwF10R0Nwe/7xB
JXD/h/kIr378BKApMr5V/Ur3CD1h2pMnyW3aKfJiDb+REFISyoCwxU/0RrUIAIZNf2onI+YJkINU
3pmKaC9qw8jC11WJHXq4lUDMFMdWad2OCEDQWD6U88rc1Q1WB73LsFjTTiRkGn02wFBN/IgVKIpW
+bIg8a7BytpPqE3OgqufLia1kc9ummcLhReIQG3us1ok6P/Y2dJ1PKhbtnii5sNfnyiqhu3Wv6Zv
YHDcsvZz5BE3D/yE8tCI64cIj1mQik+BXsUXSHO9/a6fXi/zlP6Krf8m420ktrkXXDVKWuPvN5Jw
gaQfvCYBivLOaWXfDDQ5ib2FDqVwLs/9w0TzunW5mnokzhHJe2Pr28gAwwRbDea7RMPFoy7i3aIe
bAT35whK+wijca9M6ctIw849FGRXstYmXLDvU7UbSBw5JTzg4L8c+guCYrEO8PTLW55FWFI5z2yo
bTw8WDmKYfW3uFZEMcAPVPrdiJslPE8Jw9CtPzYTgRYnn7on+E4kLJQ9A4EZvHBQS8GUvfp/3kc+
QnhhfGc5Lj067Yqk5Sc+9UczEZ+WUUAVabyI2NBoR4gm2n3g8PjAHwqBszwnYQXrR84Iq2IpnKuJ
LUNBp1GTT55bQOxwYv+VsD4U4noT7s9HL0COX4NZk+F0gFoTmltU4tbOSOC5EHPeMzSfKp+sVjEC
4V4BqNFUdvJ7/tIDdpZCZhaPNJfoopie+P9vIKq7ocs5QGQxANz1oc+h4cIvqDNTn3119EM00hgZ
zcGsiAaWkPXWwzwaSRDJgR70fFYHr6cLf9cxJQA6tZb7e4eLl+WvYwub/Re/p/sJn9cA5X9wjNhw
hz4BDXUDWOoeqTvUd5D4LSa0qi0I358gZj8UTSKWIW0183stbG6S4Od5uJMnpr01yP+XTeALV4R0
p1E9Bz3YLeGSjerFro12QFAHGef4hEtobYdFlQffJ0/Ml4sJ0f/PqNRGorWLsj3vk82NKdovJ7+B
h07nlxriQjwX98F68Pb5qqFmcEg1hDG2j149+eneoS0l37DcW/rr/5iZc68BKigtLM0OBfkmMZf/
QeDz/lkmZBH70v2NMefgd41e8Nv5Lbunz1PEzE/D9/ZW0yY/9vhdvDhutqxXNEJGSgv0H/+5amy2
caepBEZORHkL7UQRzfKTJ1FAdwItANTR2weaVH/JOio7LCwckm1UzDNZuDG/rORflGORLB0wQek8
Pwhp03li3IH39kDZtURvDARGUgqRdSRyr0rEg8x7M8XGg+7+AhNb2+k2rC4/WDb+ygTMIVuEDn3p
LSSuMcXDY0vzbDuZJlU7+b5kd5pgosjbkoFciM3IYUEQJem9pgCNMGGR3Ctu0TLtQNuePyuWBdQi
z89A2lW0MQw1sPEe+sHv/mNp6JKGHbLsriyymumXRdcT/VY5rc1pTHhTTIz9z6kiVmFDaPJCLQ1Y
LQ87auFI6440DCIlwILt9bqNM83MjkEcrcauFNeGmAR9duzoG6gYLYG3WzdBcN13oPSvoJ59UnNk
tIZu4elLzEfn0MSptJofZs7z3hcmPRlQ15onPZ7beP99D6aHjWrIsRSOLzqIrVKXv7egrrKmFxSU
fZXrYi72DiMO7NDC3Alrd+rdcSReVlkPDvwoQzJ8d0xGRajXxs+tWO0BUAidykrOLLuX3LK4vC3l
ayx+riu1sOyXGsNqzq6Lu/PI8CAXhiwOVK4mfNMlGPr3Si4/2W+kEQQ5jlGyAiZe8FIA1+PUswqD
If5R/4FXJbaSkoRKW3zUWzPNSrjnN7Wa9pm1xfHkc4tsvVz5m5ERqCTsKI8l3YG0kbpueyusJ2t8
wTvIL5s2vjvRE8hCCrk89a9jbwnzIukY/dUWuM8KEbmQsUhIO+AqbM+AYEAFFXE8RkB7fu7QVfj0
h2ft6e1WHHc8Hi63JPZH3n/YEiC4FE1EfF2/wVpoVloyYiFjXwb4ydCTjBUTIbW3ig2TDyJ9Hi/c
NIGAfZKBh9bKbIK8nS7nI4dvsUXM/fpJaif3EFMiYn9PQwlk5pIpQ9+AWLfvXmSX5vfgJI8Izs8i
+Jec1jGUW8fGk7W3Tgz6RXIM67RnCRmUPV+2DLwb3EEMmaNYT0ViLsCiVdUKKnUYDOa4beqAz7BP
HcyRg9ipih/Z0Rz5B8j1EE50M26Fpnz24LsdKH3Dy8aMvl0+ZwOp8NbOj7roWWjL4Ocj7cqIXIPT
VlOTfw1gRWCOJ/coBuue1aO3JLSFR9nbCvVpEHmfW9NFd3aknfsaJN4GVIUPgC52ZMwcKFy/i0rg
vlmRLLziptSnXhRiXu8qyVILVZYOhzsP/LI8TGRylbHJZaVemTpYQ4U2kzCOZ+haA983850KNNk+
rCjiaBU2eYQGBceZgme3VQ6jMjPKhtHxcNnECc/la07GJQ/N+pCmBScqINzDm0OYUwJgep4YbenZ
aHJlDocyIzWkLlqRv/oJLTQHFYq06vnV5Gmyhs7Dxi7UXGMvPoWSZKJUGiEgRVWvSEsa+R6OKvN1
FKivXCAXuDuAVbuQpSUysywqikBjglUVNASeVJWktwJ+LK4gBz8nMKCf26KjxqAfCbmmJpTHvcZz
6jg+i7ntlM8o5gl6EvtiKGt5Loxzv8ufJFWqdTEImMLBIh5SfLuY1VpN3DUtRxa/ezpqtsysS9NV
MKpaFHgHO/nIqGKyXf9YWdw3CaKoe4/4lZNnlT6C/KsHuyPHCQ3mpgklin1CaKXGo1SQI7w3fpKh
VJ6HtE0edYPIHiCthLTyzLxT27x4o3LCy85iEKpSKZQNsQTh6/+ARnuspPmg5jPsvJbPcctyjMh9
H/acgoNz5YYGeqXiql3aUG4Vst9h3aNtlEQK/66jtmFCHQCCb1FDlQkrFH2bnscZh6I2wntBzrOJ
soGXuYuvaDpVCVoX0XNXwpAfa/gxP34zAcNhG98kq3OuAGNWqER12k4ARDtqJ6/LAUpuVxk9oRw0
R9XNADk9flQYg3H01BkTRkpm2rMswTE+PmR1R7qQ+peI5b4WCr4EsMkgbhDH1yGAJw7mxKY1OYwE
QS1mn56Ba+2KAZQ4dONWeYC3sSwuMgq1ZVDfBY3uJ27DQDxEwaAriLbBV45MwBNXbSwN+v8Y8FcP
eYXsd/LL8qAtG7uXrO+fsoi0XHU9KeGy1wdeoJO3bj0oeUGxU00Tuu7sRWWaEHZBuXAUkiGCsKct
YapvA0g2Yz/JJkCJPFnxlfDiCQ2fhRaKM2fNsu6K1Pk71Neot8NyPpB5GIZnnkDcVzO2jCcv+1qC
AqU8/OtNxwj2GQfzH8ZexHpT37rAHZQrXnKAWE0EG5cCF+DXXa/4AadZ5COBf45uvDQvSU3lgMwb
T899JuI+9rr7Nf7q0+6ZXSmkdI7dhtJNY3OQxae96KtKY9Epn6jam6b3ymOc05AogWcTEieEeAnf
bfk0dD9VkD9GzLdn7tTfpWE5gLiIIt6SZBJFmzRuVKR+ugVXYQnrBGHkoMPc262p2viInki1Pf8d
zBTigSAfFLI6JI9HCZMnlms50GEOlubFqKczOpeEQivBjqkRUf4oXO9BFRfIzF2n2A0aDlTtkYkQ
zJa5sRSU4uPxebDAILa0RYRNWlxORjgeBQ9Fotc8SUrmWO/hBjHxa74Ntv2yzTQygzHLLOFUa4g8
ylolvwxmHY8hVSlN4cW3WKz/2GYJdpni76LbTgW0kzac7Mq+ucYtAWeBok7T4VP+8bPY9HFf1O/j
PRDmAOWV3SLAH1KnZseBrESYzAdK2TbTlxgopANCri1A8zFs+WBz0oiybQ5tvV1POhBhf5kNiEgB
j31UHwHsEpikz7rj84aveWvOKIdtmEm+/V6VNPgjr5OuD3ibm0lN99M8jXPNwO8GguieYydj/U4k
qZyQrtV+u/2C7qvhGcpDNSubXL93F1iseSqBc8F2mz7xZhaMWayOxTKsjbfHvYCK8cdn5gL199jO
hIqirkmKQRmTssog0qdXlMy1hNFP6kBvLcrtIYFfZdIRQBXmWfCUQJX8mHhFC9WnzqdveYwa3pVP
Vho8BKwNYzd8zQc0steTcBBb6qH7upZa5QWYiwHJK4wNJBXT+OX3vlnFLrIw0xmlNSBF0pJQessZ
jHYlw1la4eib3Ga36IXZOx2lI8DhWfojRLYj7kY4qcBPNHEl6EA2HSwV7AvW0DBmgBQdxW9nI0ya
RdgBMcXGqr/ECTnp4VnwQGCoQZVWxQnADZAoVwREXvBDguHeaXNutJl2lBxf644ejTA4oZISHvtg
NCgcVANrWVLDg4GhAGLE7ERYAO3uGug9SoSoZgALr09hPu4vyXu5JW1MjkNbFGsnAD0d0OYCSJkc
3er7ToAYAaI7hJ/dtGG+o5wUrm0roSyyj0SMxYlVkgi9bralpEy+r7aixCY/cI4G8IAyBo3UqZ08
iC1uj/YOINf1YRSMEZHnN8unM9M1BfSX/1uovwbRYk/FrvGrYKpypCCEEnVDvOXIEEg7AaZSEM5j
x0bUWo2xcujUOPUjh43z5hB4ROJ0MafXAxE3C1Zz8f7opk+KwXJU8ZM2ZplGpepfx9JtqOqpgmmd
JXxJKPDX7AIqfN5c+8wejxPWgIjWJdedls9iDAB3K1/qzy+EJmfOCRmIm6KMvmgbEIukYVJ1etyw
wH5xBRMoWpGXboMRR+RJzclcufWrSKLxR4C41cqVcxdhw1SeXRmogUmdVdecj1gYdaZTZRF3ALOO
g+PRKJ9+EWQXMS2/y6rp8Npv7iU89FPFWG7mIPGllV2Lwqkqnq1+edYFNoI3D/pjChY6RKCbPgHe
cnXugQCUzD1OKSmUyfaOTrph+MWd+065j/EPnyjbk7rqUr/emFWRzyWUUzbcQv8Idr0FdRu4qxZI
fX4dOdEi3Zb8oSZFpDieSgJmG2PWhhw5kdhOEd1SQf0pMaMLuZUg2CO15OS/gTHul+83q/BAH7Mc
b3X8bCrHpag7aHrZ2bhAJL+ZaK/aBUHOGQpCmQgHW196nf39k+jW0VrHPYmmyGbzsinaK2uzqdc7
JPeE6JRy8/oSqlFHSDPhOv1vt6JNSavAc8ChZnzs7f0XlODfSaaplBW34vclZQDECf+oFLDisq0c
Rqq+xVBXEa1rQb120OO/VaMNDCP/S4Xi1Kljbjz9zLR5rIoXgeLwEKdwqAU8NCSvl/qBgrxXpcY2
XJ954P8BkIKA1fNPHmyohxxeRpgOiykgga6tQCc6BnQADFOzrBUTrg0Pnr+jWUkuDd4t4xv/rs23
MKIPSyc68o/Devog7gbsqCVF9PR3oOftk+3cADcDdNKYOKfMokGmFiPOq7G9BoYLKYE0Jq4t9s7t
zGwwIa/C1L24eJ//VQNXgISXbaPz5ehocDqnoO7mCnGPH7QyZE36vBzNWYHQFZ5FUZjCvcgtlRXd
lO4rZqJmnDvO8Z1ITTp4domC6Wjy7Bww3mGNWH+KxtLe9Sd93uv2cLwPTin7ugkpKmnMxcuynQqy
uwuCK2WqN1qz6hLBXPjlpUSv/2uodfz0zFGlXyHftHyaa48IacNarhCVBjyAr8tT6NYD7T/IjIG5
jlJg88Lm/niXiiZBtq28a59T9JsdnvCXU1q5xGRxx8SGmcrYkU+/immu7aN9rjVXeLuTDrpvxzbN
EPgaTJJlGEieFfxtovVbq3iiMvI3eQCIrWSxdPK74TiL+oWL3MaW1VRlJfutb8t15XQpuz91Ml4h
TAIPq0yMzyGILk8ekeEUK2A1PUIktD60myvKZTRzvYXC0SkELalRI7TOwuPZvcEW44gGWpjwZZ5d
TzJcx383X25GaN1psRJhH53c7pmtadW4Max0SsO+3q06VJ1np9ikc8sGFAN4amqKv+tdzZXRgWap
x6xk2f4YN4Rzuq9LCPYQkGt+grGp419fDsNLl+016ulO9sOzqhJZTvTwpR16DPO5edkxlophieii
6JHB/rnFC3EJFDxKEwyUdZu9A5erNQKh3ABELipiYorCebmdTw2m3wJEDPTViGd1rR/X+j6M9gOS
hDZv92Oce8Sol7y9nNP+QBxRYlEBOWF4/LTpfDkiLgPalEAHcwsfdt8IOM/mi1DprlfmFtYsIg8i
WXNRgAtIPYo/gJLMB5V0uIEkVNtnn8m8CnmBSc941VnL+WvEaYgHvJQWcGFm9iuvS8DHn9wBqGgi
qHA7wyzStOELzfvA7U+qHFwoTnLmMi+1rc2JoG8xXOV9mfx77bEwgsz+X4E/itvgcb+/1oN3aYH1
vVk0M74/Gvd6RNXFo/BnxO7UxJMZotrRBoZmpynx+3Zc26jjD39XWD6UjBXzQaCuFZCmqNkYmV8O
PW2ySfwREL7zYiJYUMpP+2TpG98IWEhf/3s6zkk//lqJMyM+RjDdwlGFLaX+Uxy+zM/O9EIw5E2p
hnhrU3vmOp54fMPR+cQRYKEFlxdAIeinIdcAJDM5kdVST0mWnxIFtwE6b84kTwODWLiAHkheZUMc
2LPAZZvNVr++s2tNV2i95G7jG+a5HYIexdKd7T8OqT8mJ2+H8L5aORHo3kt4oULtX+bw7DC5y2O1
e6LIf00UaMevl5n9lOlSTBwtCHHE3F04PRY6v3SVOwVrGdTWwyV/0lfLiW7ra90zPikf4WW7/jUI
x4bW5HfLyPXaeP+sT/JB+TkXP07HPfdB9oBEMxEXwSKcYn13VSgdKMzKS6smSwIlmPFxVX4kcTzK
gGa/GfybZpQ+JlanEL6inL4/F22he1JnQeiS5AtX++qs/QWEy+kw1LIP2KtktEx7TcAry0X9QGQd
vRs9xzA+b2BFvchkxSvbWhMaU3KMnDh0t7vIhP/2o+Wp+KN6KzrxoNafVI/nNV7yIMOz+Zh2S53T
zcLI9XwiWg5D12iiV5D8Unq0+Q1OcR5N+3rE3aDO+IgSjvxKOdfUTUbIpPb5Pn30Oqd3Upgsj5fw
UuWfS1wkKC0xOs5JoBL39XWcESuZeCQxRjcSlt0uU5uMNOUgRjXXE+qO0xCopVWIIjil3gXO5bs5
YCyzFZQUuXG/4/yizg1L8i8Szhpr/QIvNoUOT0mkkYTUPeoDXfeq110Ur6dqCtccDXEF3yVYn8Q+
0zKtn9Oe47iG+XSFBDwv68oR6lR7KgA47vP8CZfhTbOmg9d9NRaz7MJ7Hg9Bgp/1RVwBaFRj7znm
kM3sCtmHYTmNkFk1K3sm8XXcE+x7b4MAXym/FNcHOczv89mPMD14aC/IZXVHOEGVOvd2JqGHxnuI
LkVJsCJ5eRgcRpIlHFgHniBnbvj1O64qUEIPVjEHB7sSNN2LKEGxSEGwSkW/AB3IV+bQbD9J5lh6
pBXDOLBV3gGTYUGr4OH+aOoMji3zq+pT3uFF/8hYyKgbxf1kctYjljOmL9ireaiaFoSm+ijqERzw
GgAeL4n0iy8lRF3y97E/qKy25qz1xcqf2yNHS/86f0jaQ++DKCEl9bvgS0dzeF/MiOpMAaR+NynG
pj/9ZE1bPRW+rsEJKm4LFlhSjEDG2c5l0Qp2iMK0NR8ouSvLS1thSMREClZ/oHv38q+i1ZNB+p0P
sQT+QmKqVodrcdqg/LjtEue4Qi3ughfNvj5g87HnSIY5OMveX4H778bU5rqYOOjcFSs9wjRW60kM
whAkUCOmK3schmGI966A4mBczz78MnQqs6KxL11XXWIokjQJTrTAz3uhyUK0TZpFfBEoLAo7m1MJ
/HobRHbJkTjfbYlYkv+ZWqjlBmoJxDi6ZJJUGNIkeA1lnbhnhpo5cIMwG9x6myXJ7P95iG9Y5JZn
m5aZVrUwe7R6xpLwglhTwqJVnlINrTUqq878tOEB7M5SiA01pMbHRKx2c2UUMDntFDDuvww2R2nj
ZOvF429COgybc0rKLtIi/ZxE2RqTVKEyze6JN7IzFJKM9zczsYrBT8veDP0Ka2k+040o7jmh+7Ho
h1sNeCE9wlrEDH06KdkR09obx/F7v7QCECOoXhhnNBy7IzwDGpqY2yM748nE93go+7Jyjie9e7Qx
DHVJlBl2p209yvyanZ/4IRhrDF+FEZen9oz0o8PkTrYEa5FqMjV0dvWN4VE2cf6EeUyou+Y23+LA
5DFgh9f7ubcx6wdI1ysYU3+E5sVz2y3A7jfNgY4QXii/6yOYHbcCoiXLyksnW+ZG0y7QfaW5OShI
UeAUko5zeCvFi2m0zlVAtqaRua721nlac9rLoP9VvXz0PmOQVE4ZlXQ2r2uCKQTkjw9ocmyt4QKg
1ndaTBNCScqnokvFqh4F4VZVeFZ7ObmoU4YxBViBzIPfuyUO+Wyy0H2MmX33unEfx+Vqjmr8Uvwk
RPE3q13+bzA/fgmbS6vDOTo5DH0EAy9Hz8cJYnfzNm6okqWnzHeuYd09J+35EyIvrk0xS7NQeZjq
VcY3joq5kGh0CRSgqK4Xxs9FhJ72Z9yVwBbh6rNkRodxzNTg4mTCNmXhQkdh9S6kO8c4UL3VMakE
cUYk7kQQdxA/adOwZCI3qd81vjy4ctJvJl41WOL0HFN+6VFxa/wrHXuCVDRuxIarQVm8HD3itD0a
P5s7Hq6AM0YHYK2SfqB7Jv9+bErLj2VBtXcgUF2f3xNHlpjX2s8/ILRghq0mPT3Q18aq5GmUqg5U
VPQSAJwBgqX7crgkbav5E6n70g/vXpt6WavGGZpjIH4oP1obLnZuV88XQ1eAyuQlkmoJeuaW3VDv
MEjx6KZg/weUczbOK8ZhS0CI/AbPQ8KyYktkNZBQZbJ1319jSZqMwUP3CFc2Pq5NPLjySISeGk1O
Ww388obC+uWA5m+BX6Esz75zfGULejYYMGQasVKHD83Lzof2axqSezGycJZGPXETH9OY601RX0Rv
jgEC6H0DrfARHYQgPFQY8udNPU5gR/TYyfJF+njXrL2qf8sQX1m2h3TRNCOVP9XI57ed2Lw9hUTJ
B2NLqK5MIZp/G53d7EF1dRl3KmpEp7kyph+rZ1m+5xnM96TXXN88SwV1EZPl/HWjXkkFtJjjruWM
DbjR+kPsRVexDTYtwJAveQdyUqEOhqzIuoSFL2sGNAJnSj9PZ8c+wmDP4ZkFMWAAJt0PjLpBjlc8
cpcpUEUps5zc6IhWKxbooiEsCJwVDmufWRhZ9VEwtR4VDd46rKj3/30tneAqKSBrfsty1RzdHWok
Flc5D1IPOXYbdAR9tp7Fk4pBcTvUL7frLPC0t9NCK/D3xCIwVBFmGm/hLXfikY0/6Dr6w42UkKhp
Y1J0zYbNJ9OgUb6+N6gU4+IxFSMVVttihDzfjIhE6HUSRe4/UYDefZ9UhoNg9jVfX3fY45NVLweZ
2FfbCagsqE7qR5FEq4kDr/Bv0/1Zd3B4//tjED2eg2L2S+e0fY4deVg0WfA56DZ3dH85w0OLY28t
4niqN2idRK4ZK35P1Yv/sbzFe39V3BcgtplJ4bVtDyfQaC5Rj2QUsaAjAYDxkcsA5NFHLjJyZWM0
DIMmxcJPPUIUzFB8Nha69XXTtch8jIUGP/9VMD0xWz2UgE4q17txmN35lGEKklZsbQ0rrAq9AUYD
GdUVvSWU7o6asHcDMjZxCWo+PFRtXJS4RhOraMJ4yqTJfAOwBBxJVD6jhdq1T13BXcT9F+7vvG2U
0sYKmf0/3NEMt+gQafP2E4IpDaNVgYCMn3cUA8VekpBPaRjGGS//3SSiYaUp/at2kfw92MT5kngW
J7F/pglTPeyccWQi39xlvMlgPwXn0F6dpZWYno58mA1RhKKiZbIOtCzPFYC62Lt7gbJMQKkrlRRI
XTSATXxinhwUpGBGVbGe4kOABv+ZGmzUnbWx3AMmBSmyOYC/CPDglT75h7bs+ohx8qL70QZ1ICZ2
EGRbX+c08cUE+zrqhvuVR8M6nAGhmrZP4PKQwoL0CxTZllxp7jtCO8huRFaIzqJ+U4J4wlOaerRn
7zFrsYRzvxu+Zkm8f3xP/EqMMtNN+xfJ0SeRIo71MgMWIzTlndr5wCflZGboR7EJpwSUUSvfg/7N
xpmGS+aiDiOHUttyjAoyKB+5y83OUNiJIKHZ4Vb1Abek3DyFC4H0Mg4BzTjmc8yO89dOLJDcA5y/
s//6gWDSkP15eiTi50XRlqj0QpgVbyDOhdDsFowCbDXYmHH6MffRNTRERGUXdSG8qvYPRdr9Ph4O
C+Av9GhAixOcQbpNqV8/X2pJn3L51Kug+xII6EEYC15j3j78cCXN38cJmpQ/K4WZQ8yovFKKMaaz
MzjH46vS8hEhm63w6wC6kSkLcxAH7C3YQOa6VacqkWDRWzJOsU5tQMRow/YF4cqAowP5GQb7aZg8
rCupTrTfUcBj6MwyNPcAPhJNrkorwcZ8CkjY1wFtFTJz3qjT+FnSxIha5kQyUggcsDxdpkp5MSkx
/ygkwyGxuPcHwoCzILzI1CC93sxQvTdOniROax8bbxuJeSqrygRxEsjURzRN46GCR/+5NJsHRDlt
sFZOu6q7RYihPeiSkKO4KLY0DE0Rwa5r4lRKhgsRniDsTYQPPhQcxpNBhHXZVGwgtwBnKHxVW2O/
f2z7Q7P3kSA5ECmnogAFiyuxERoB7laQz++082ul3JHHYXeedJflUtyKSUY87QA5DIi3Lj3mh/Tl
/XwKkZdYsI8xICMR9HqHu8PAyOwPZnhC34q6l1MT2N5MTdhtWwFNkKi7f1mOLYaN25XE3e57gKr6
ves5jXKevOIUng2uENCU+koeD/d/afr2ll0MyYud6ArUG4Ytl3qE6W6odmn1Ep2+65VSZUenwn3S
wUkWjvpQzPHxdRTuwB9AjG95b4094XSgMSnGuGMsGPz+MK6n60E4bCsqs4Oc3+z0TSsfQTGkFaB6
4Ae4isF/zN70oMebrooH5MXMo9e/ijzIunRR9oVJ2qD68woFT9DNHMgAEjECyIuDUZdd62ALgTRv
T+pztf7zbDR/ODdEseGugIbV2xbLV89RPdmykWIkT9FOZnFd97r1m530motqSwcx41GTMGuiopNn
J9LenIQZ9D1dpP2divbpStBS+T/fipKO9NbZ4IAqURJr/dNBxv7NdSFNKAEUMSfyH/NgSS6NWx8+
daZgrQ8NdtA2aSWLKxjHVIJoEPrQyEy4GkFhAe3LzjCIfFdpQlUlNAcLRF82sz1BC7uiDz3f1a+R
jgvcIpr5mgaLgENpYA7TnfLZhwAZDMckcZkEHGMD98CQtuRzkbA+EOnqzu5TO/thwtp1tyBNDIlF
4hTAN7HN+M7XZ1iyNiVj2FurINSm2D+mCwAUSXKO1v26yDr3hCQQ7K4OG/V8a/RGM58hygQHxDKL
8Sneh/roNKv1bI5YtvUVGL8C2WHiSkSZVe9bq1XQXpBGthWlCPlBoqvvlET40mskbZl7aspCNRTE
+3nANzLoHAkEqDtNqnBtc4iXN36GYsNZUoerXLQsAH7L+AjOM9x8kvN7rqhMiE6+yuJi5VMf/2G/
p+Ne0sTqtOeekRFPSa9Q2mZNS3Z9MAMgIqh9B6JTcyn/n3G4xoPJD5hbaXkKuLU3vwYVdtuESH9R
NEwEaH5LoNlG1dgwQ8FpDB2u6pOIlSEsGKES3ToUbaWcAFPDrm6N1yQnvYGqz+zBQnCrTOk7ocht
fwjmQ2OtHvg+gAz+CyWUpUqo3NWEox410N2j0Ye8jW5rf84A+4cT++n+8QW5k0lZp9A4G3q7SS14
TT23P6f83kWE+OF4FvGJBon9Jv70Maz9CH/BWxl0LfvnImiYXYWwiTDwki1wI+8WcgMeKk70vGIM
0n1zaWO/hZHG4iNrnzgrQ7u/mUeq4tZ7L7s/NoRh5+qFnnCWDrCmZJIjKIJ89QUdG4rBPgHXwrfQ
F6snUQQ8uTdYI88mJ2WDdkJ33RDeuSPkUk0zZ6PbFXXz2GMVnhBgS2KruJaMlfaKOnuW78ZA4L6Y
pe/bgdADX0wLLVWxIRE6DTDm9dTFgKxAJTzM6IZ32IfeIFaH3RME22hgqmbke/e8/LocN2Gpf7d4
ZvRVwOawFp3xwXAQontsp/MWPi/1rb/Y/nz0WkAj+YnlqVg46cu65RIrqJ70Jn3vNgN79ZzvjHJh
7mbQWXV+O1oj7ZcttI+G/zPPVqHhBr6vLCKwP2Gb4qHTZeLryFAacxzkZwotJ8oMVIEF51lMdToB
JnmsmhP6C+SvrI1O5Ga6dcIk3D+pxnTnKS7K7G6/YdvUVOLCX8sf+LDZ5838WwWonD2sCVuX/HYA
Vvg06/RGGva+XYcgRQogQo31OY3YmojOf1lJ4ROaRxwtzYomOAA4GoeSgMeQY/oFE9tHLZ3PPlVj
Z9YV92/0sz+ikR2b1qIzHVSXrErwL0bfCNP8/IPhe6p6ODhPdVXG22YBgcuurS6fXVY6btyudEuK
4/hO/osK3FXa/zkeHus1OPtKPJN7BC1ijql+ZASHho4BD7BUI2kut+CyVkYp7kRmbN1RDQDKDgkX
XWnwXvGMeRVbj0WvkMaA05s0embvMaJSvjme1GRsU5KzDASrwzydNiqgeISz23uLubD0Z3kdPKxe
ISb81xGB7N2KegEPw7Ovp6LsWbL9sYdp86F+MnJsT5K331M0OI5unObKMjqeh/9j07GFfjTpe80B
CXMqxnuaQU07LfLeYhdfwtXsbjaTQaT+aVXiyA1lp1sWSmH3j3hepcaqbQBUn44iq+Jrjilab8N1
WuUrSTudU5NQ+RXIiS2sJ1YSAzBChN5qCtxshyANvETe1c3NkgLZfrg/24uTl3EiILHFYrXhpF1C
qIGO6X7sMAaPcWRNmRAdDgQ2Tb27a2DcKhvy2NN+KldTdkBDRPITeP7zPg7sxHsEPLxcY4tHjGJ4
F4SS2/CHATWhbH4AFKXpTyBSXPHLQ+y4/pWhj0JnK/wybl5vlFej9e99VvoLRLR96K8FIQR70YaZ
HCTU0oQj+fgLYolvtyQK8CYL6CphMSMuVGLet8fA0lbSAL29+WBeeUFFCNOiAQoEVg6WfuQN2/aM
RdnTinm5gudrKSReuQVYGCJBMSlKrcCRX0NpOz4/zGYKtK3e/dmOolbQOfkgqM8zdiJn+q6XpOT2
Xr8dWylinDux28ZzArrQLP5uPiKUgK9XxVYWtTposCMo9wWICchZRQXYFpPR668K3v+x994qHt9U
v46P/h+jspdf5zppNz0Q+CdgtbdgtrlFl+djMiZGcfY/OsCmpBYMrBHVqnrxXc6b6Se1FemTYuxa
PGEh7HTULX20ktADux0os+gvr9A3+iRzdo1byDWIyv2fHjcntN0C+RlRXsmELTyXdhZRYtut83QE
hykWiEydqSP+qLkVpjIJv+TeZ6746tq3eF8lBWsfkDpUAxNy1foPzrnRRieY7Eo4MsbHAv4rrm6M
hkTgNel8J2vtGNvQEUP1s0jw1t4hlbT+3mZQTEQoebK8EBr/zpEnfPBpiijAyNhyfBaIL4iPhW2b
2rVpvay1+fCCY0/WxrCsMyiQUPFK8QFEljT6C/4dQlzu8hLoanAmaUExOQnD2uS4wtvpdTkf8+G+
zW6lPgfiHlPKB0tRKlPXefAQQ2PiAff7cy960pQ80x5L2lhemdTy7Z8vbbHBOYET6QaOwS4io8we
eyRjSYPX6z7EmzGs+obwZQHNR8wtNMeEdoivK+qdwsvObDmPy4fxMEwdZP2D9nbvu3nPKDBJS2b7
YGdTj91TNI+RYJhM32tlUGbk/y3GIP6yK+mBNpZZHIod93G4CnFwxs7F1bmv1Xsw0+0gXKV37cOZ
9q68YiZsI65QYZbtT/VyK2YZpxgLXdjDOeV3ZTAR7cyb9X9lW3P6J11IIp81sQe0ig8UKIfEIJeu
bWB7o4scniMGD0/BwAjOOuCrvbarA3jdT2TJ+88fFIz6O9YHlyhKnSt+q9A4A9GLchuCyCFKZhgB
55y0Zg6X+1MQGmzxe51F6JrevyqGjUir2015pdTbDQ6tRYzhVZb1aaDaEN3AICmMJUhU/FqV3/qb
zPtzhpy1tJbcHqHfeZ7qXugkKN6qQrgkMkTJd0CPuDXmKMGYb5SulJHm7B97ogOpFcrvLS9zEeSD
w4CtEzcpO9zs8t3kYuT3gAyO1r8AU2qAbmOWWFLdzJEcb5TBywjIc0SvuuOlVSNc7F4ymjCZUEYy
0hktWIOVT5IZS8B6yjw4hdGxpKIm76oj9BnolnYYh2ZYu5pqwX+nJAq2Jc5VYG+agX3Vf3hHeGMt
jBuZV28//7ZjWAgfLr2/qTjgbRLCCDo3slplN3J7oHSHqnXjPVfLYU8IzeYGSthE61b+obNTqyxM
OxvYxSH/BlnwBortj+y5jKjbodndoDrSLNny1oUThR1XZM6UVGdEv5CJlD1rAUhLvmpd5r/G1Lzr
RnWwTl0KXBzZQ0mrhiFwpTeM4Wle8mWS+3wFLQrFsa7ntvlGAaTJaZB2D34VzyN+HRZJY2MzhTL2
tFObj2xqcRXeRtJnLMVdYkt0uEIF1cB2cq8NhxO4km2v7yIkRu3zrXQ3nAaF0G8nyY6xQ2rgymEw
KZ3Ezxq41hYitjF66VAvwLSSZqqJ0xc0ORwoZV4m4vCBW4OwHZfgeN08M5oxDNK2h1PTZ8Tf65zU
ueKcMJVlQkLewoL66yWip0PbEF6lE0nJXbrc30jXRAtoBFTECCn3C761Lfxjpu1DUDVUyLLVGqBF
TXx9tYJbEbifpOkSutoplQSSF1kQqygwu2s11w/3/GLRUNpKwDoIwgLbWRx+9jLoKbSGcU1eyTDV
QEL6ynNa2UOYUrxvvcojO4dwXe38CI09IjHQCdWtPdMqp+xgi1TtVpBBpWrTjC/KZFrsR3P12W8T
rLQGlvPO+7kWm+AQD2/BDozYqu5sH6M3oDJ3aWeSSvttDBfXBMqZMwDfvGpjw7qM5Kp1QR/cf9Sj
8+e/HmFIxNX8mQnM6Q6+DWCcZQrI4Osec6LUJ8HWz3m0wfQ37ckvX+reCx+GRwhXHmcdDW/FsOck
rr9rO+53kbmjp7BzygYEKT2zj7dtIkCS4/Zazj/BvkVu1/FpmJJ4ICxY0+WIZa3xoLe7xIMh8lBb
i7GdZDdYvJ063XyJzr+FmrGnEUtNuQ/SLuS0dd6dMv8+2sq6fCKL/QwMS8Ap53PGBMn6nbSLGv9y
UGqfUIduUUCbxTupe404pg/3OxFeCipvU83EWpfJ+y0mzX2VnzEsDL5Q16XT3HIcnjIhwmEROC0h
98+Bw+mkfYmn0dm+KEBeeXCDbg8zXBV88T8WlmWovRxbfeEVN8VJ9mPZbavHJWQkYVXsrXdGQeg8
SHUarvXz+UECEhhNbHzyRwbYemKJJirmT8FsJGECyJZUYmYEZFKod8vFSH+CHuV52P59921+rb/z
GRtqwNm3L1jMMZ/xuKkJ2VogMBScmpiWgyBfOgldVE0qTdJozHx2SRH1GtJBO3yfZJIARO70Tf0U
MpmeuvAZkNy5zabHAFa6ObPjaRNc6edLYtn3oEWBIR56xx3L6IAt8QAswo0eVUaR25xVwE/gy+xX
OZSKwcfZrZSr2/7fGc9s0ENRzVzomzD11utL0LaGaVKVYe5M1890AS94FDS7Pwn3FY397JQzbyYy
9ZJ6+OXN49CA7ZtTy5NrmTGTQKxED4JcXJTRjk8pYZGzbr8oASjLrm6zIbibedVhh2WvwY++VHdc
qG66VjoMo6uUqDu5SZtQHIBjPhY7QXoWCBXUWvrPjn5Eb/i0eihTzWZG/wYLbryW08kJ5GcEIFGt
8cm+SX3yCc7P4jvwF7OTOcYqAgBkjjv3PnryWchSF3YHmiCVToOjGGJkY9HCmZYaQ4yDiZPxM3Qq
Ue900eYR6aOXmzV0T4O4MJ0pk1lr+SaGa887EyXUW/ICZ/c4dma1T4CkrayRd/CH2xznq3S8o9gp
estvKTrMYzX2vHN+/AylxOg/sgIIAtBHzHNfgpqaJ7lEbwp64AKQloa0tpR3DrC8ibO9v4Ixzp3U
wCXXHYYG5B3wO1A8ol6tvQjY9KL9dJR5VRurlbxurfiknhv082OXQp3oS8R5DlEDP7Cc03uOvdPp
hmos5EMKsAgX2OK5OmjF+xiPQ960b+4fzDiM7juOcmf6G1U58EkDef7zoB4yVcAi8cUHoGKEhHBm
qMhxGh6tv9JU8JYw8BHPGykvo4ZsAuHgTwJeIvZM1SPYX6hHqWvNQ1sqXrC1s3YJAKgSxiTby5jc
e4N/A5CDMfNyXrsU3VWz4mPeH1fNHQRxJ3RHtUZ5H7MMcKAKVE1JfqhTXQTyOPqCQuqLBd23RCGY
tmtMhYaLBLC6ovZNaWAGKRkQQbcFk/Ds5iIKx1NB/9/I22GPr0qL/IB3RVdoDRfBKaT6mYFRgQ2U
Cug+bMj9Fl4dDaPBzCITkw6GJdyVihWA4QYXIWwTBEIJ1+CSr6Y/haoHnrNFopYmO/czOqU2W5H/
HrTMVpiB6euVAE9yumAguMR2B4csqEtIm3eokS8M719jGrDHCQJ+evMMEj9x15rgyICwbaB1XfXZ
3NVpAsxwL0vTsksHMaG3Flfh2vF53C4IfuBIE98s0FLeKdNgbGb/GIRmiuLz8ZXSogEd0s8hNOqk
W2yQ50FuE++RPo63gUTdKft+TPt7qs33IJQUvFPrsfD0fpFBuxuDQ1dnhNo63r5sO/EIxjqGCByo
ZGp2iNsOZnF90hA87zEA5IT8lt7F+b5yAtlTOJov8X/qjXHoYC8JgrsWM+zKRtgDEzD7iT6Z6/Wb
fVjpYMqwfT2ZVK2ZCTbz9+Pjd/0bliSZt/4kXkiXE9lRPAqA1BiqXiAkGqtxNgFPqAKyT6ruGkZw
DCOK+WgieXhw2JmIi8n1g4T9TqkMFcvchyK/I3NI5Inu13Ypv5T8ly+ie+KuZzqy+8sREIU9Kyoa
0XwHluGq9aGVMrggs86iRR+JgWE6KXa3u7YZ9W8H2IwoKf9AEaS6NC6nF+L33fo/YNnCTHdx37gm
8Ljfk78qqo77qCneaq7M7EBTI8QOMGaxVScHZeD66O/s9Mfu5RJjzOjI3R2x4x7fPrXbB7YgiMm8
/0Tadf+GmgapetndKNGF6nA3DSgZIasQ6FuYfcLS29uR7LTMcYwS6cFkSx/p2Qwexg9/yCEywEXB
QqwzhBI1CZNMMApNBo2juIS07GojhBnS0qcy9tMZ+c3wWQ/lBfsrVxxK0HNHmI3qYd9/nmlxrOPF
AnhbCROQZbvZGkNU5/hIXPIhD4SeZYdGI04vcw07dnY+Z1vhR6z3PQfhnDwykJw+5c5B4kh8IEHZ
FKAis6k9GqDLQa4aVJTEKlc6RSctdg1LpHEauYY9n3WI4RpJTyUtutABuGQ8UQPdpMf9EeXY/0/0
HE29iNNf6Jo86ZayHAzjT2Sa4b0mFsrLfNVTVcddq448cjy8RoFbv3daZ865BK4JurF8XJyUippo
wf+Nh/8tg17MzAffXkwzDTj7dIE3/SjXSnlMru/uS5vhGGgT+0OXRNrXCK/TNyDcsvrYaZ+odSfs
UHmTUogw3A+L278TTZNa+eRhoWAJR2wlec6CH41dJl/07O+HyzptOPXLkrBiohdN278nuzWihQaf
zcw4M2XxOu9CUtmvyNQG/oFA7TMti4UDFnD8X6NAniKav0HOPpnIboV+1yWuZX4h85lgBOupAH4d
nURYJuJmsAfA0GneBlBWFRo6t1MN0vbJtHm0YsftQP4EmZNZ/P11Nt1SG8QP2byOVC472tiQqqDZ
25eI4UZtk8ESfAzQNnWEUIr4sckUsPD7emMTtxkR/XVg+pkcytv/1Lxwp1XYN/V3LGPqFnmntLey
spFmOAjjoXlNsm/6GW6jzcB+Iv96Ezg04bSG0zBuZ6TV3GD3QQUoCDTX8nQXOiyPoEwtpwXeE7K2
iMBpydMoCx9QxmM1uDLOtlS3v9+zCYV2mxabSqURqiVrrB5D53qMIe0auT97UtFsnC7oNmpPC4K6
SR8TNTaIjnon85NYDpJ/gqnrJdYkmaBmRW/PiDcAVBhC6HGBCqyx1IAd+qxL1EdSFwHvHhzTowYr
dxayl0uC0xcVdl2O9BxCrrFLgCrD/ljZha+CPvtqz5Tq5nJfs/hINGfAc5sVFDc7wLyLrjfvh/Pl
4mZ3VNF60yHCksx0hz5PpGNYuBC7ouCATqRK6GxbY8klNcMovIBdXErzsSIJhANiEW0w0nHS2ULw
PWroPIY5zRRme5yHE7tPHfOXlRPFrP+Y7rOvkY+ZAZBEm5l3li3+3gTNioiB76jdQbFntQ+0ghmE
9xylaTw86R1xlwDAV1fk9BnwCq0FbgF5fYVr84HgLz6BIaK4Hz80q46QrnEUD/qSmoxYc9C+muaW
m85en3dhwXVWTG+UAsrbPm6UhMj+JFqd0WQlwEo560Vhh8VN4lGCLlslPiZgcnjNBOLG9W+HoWGD
FNlsdTAlkBTQoDK0QwqRrrFASnQU/wdOGzBJ6d7Ln5wqaxANWMMkYAFiCi0dUXW77c+KGD7Jjc6Y
HzVLY5WGPJBQi+RS2WLGR7ziDZD30It7ARIjo4aQRuuJtOUKo00n9u1skmmAz/laEoicB/MWgu4M
kjvydTecH43UPcCIvk9DNMs60rTo77hA619+DdP6+ZFUQ+G0bX0l1w1LvETTIR3myCYa6gryxlw6
GawtHSMWFLwcOQZhkcVUWf47gQUBQA9LIS0U1vjON+nb/L8y11E0RPHGq/AV8ljE5bn2Od4OcmXO
MdbDQ1LwAXLNAcfDmOrE0HtolJvG6FZJ05ig95nx7fYu2aQ80CmcVBf+N1nAw0KRsYvHLn73RxoT
YXBVEmP1KtfU41QhFFGHNHmg/Ky9YIoxkpZtlD3RD7LHCQAJAY4DjnqhgbgMlbv8Qrs//WZ1Rg4K
euAosNLsLffUaQtgPxtqoYgzzohr+5NaHWbsRkeDVNeoC4u2dMC5WGE5JIeATBXxBLYoc/1Kzzbb
GdwdzBVFqvjHIlHhGsWtawa68exaJPpiqnO6EEGgIkjCiKAeqhPjfMEmMz15y85k2WEbOLazOCEl
JqHy+EaStH/dJEs5w8uaBK/jYyelMKX3aUVaQYGBhAJcqR4+JPtNB81crhPxqG5k4dxoOIp72czh
T8YOFQC8yPbHIvydV6GmSPFgGCuIuCdyGDQa47GhfpSzBrZKesrNHvlrQ59SZZZu5+L70YKri748
PXsuQlsxBPsrkAsoY3pw2SgdJnxJiWYzxjfLJETWViiC3CM0oz8m319XExvl/AY98NYqnIrv8n5I
bwMU/SNQVcLQg/BJj4Ux4AEsb0+b/cw9J2eI0y0hT2kDm3LXu/H3RW6CU7WitYYMGkKSNocQaNtB
MQBrL/1EcZTVz4JEJXlCiTaIIerKpfAVCBlWoAN7+KzJz/vqnC7WfeVxfIjz5R/vIWr84k7mHpu8
dFUyHb/fJ7xrBP7gKArDSLZ4F/CPc7XYOS6WKSns8R6ySxgWoAkcMEY5eepxc+bE0MPoWQA1x+SH
/z3bhbXMMYbzpI2Nvnlw2y7VQSBEEq/DtVJYHBPtbkeESu1QUgV/4K0QpSjoo9BTCVrjjfQ5BzJL
haiqporVaZrRtyckwud4SIWo5noV0Zynhi5imnk9oi6Qc6wu5hj7FOZo7OOrX2HV4SmTlGt0XcYI
PA+JnKU7bkg+0k67RjZPtpCDHzGMwni25/1QYr/biaD8xYJLixYTGXI1P9oCgoVwGpFAh5OzjrJw
P48/v4UOmTFU8PewAoi+Ud5TnhUGxOS6xrChlQmST31mwustu3At5szviX6Mza8dIqicJuc/BnuC
T/vda9pRFK098k8J8oUpeO2DBDorw9ot51eHm+8uRv+nINCRRbzZJ3U4k1+KTZjEYVlezUygySD+
FD01ZaEX9tlJn+uRa5Cccsj7jfQQmyKochD606OC/+QZ3waUisaTUx0HqlI/J+t1cjqtPieYScO3
B4LmC9k+V2iYeKs/gAxdS48wLfstYBEq3w6rAVPIy5CJillzv8zAGFjGVT/Z5aP4yvjILThh1TJ7
oMek6Sgh/aJG94sc+f7iQjP1fspkp6NYywn01aDmu7VTmGPbZ2luu0i8+qpzxLHT/4YpuqFYPKxe
4VB/6aMjrwfJWki9zBRNPhGBJ3x+Y0xLkfFOjfuuRkaJgyMSF6IAmCXNKz4S8xHFiaAl8OEqZILv
4WnKN2Jq2QlToJjZLY0yh8wruklmfwqz1JevuCCcE3XlVSiJnYVbevmo/EsLY1qvAtPLL0DARd1+
eeCxYbTApgTxnia//1bag3OzNYgrffplaFylTaLLk2rTy5fzhLUvBYon9KR9+z8RPY1kREJiOgpj
hxqmnfnnLF28hZXwCQpwNn6pTxoA4UVoReY4T32MBklIC7vl8z7Kr7+ALQgEORpgSnqL6gDngIFJ
4M7C2vXTm0arugCvkg5p3B5Va3GsXPq4SkDvbAllkcfAc6QCP/ymzceG7+rwIa/eA1dHJN79wL0R
S52beKfPB8UnHP43Dw4fF4/Zbea07uDjV+D84kHWvPDUKXVi9GmO+lWNgr5bepPVHBFdHHIaKFXK
v6dvuAc/zE6J9lf7bXjztQvxjrxAwlejnO6a3saYAF5yTERtVp3EAJhtJP5+xlJF4hxPGpY7cfc4
KSTO+sk9Z1u9cm1dUI+0jhH2d5boBKQy3d8hD4+dgcHa1HKUrbelYjPmiHYWCm78+RJT1LxngDLi
m1RS9jUs7tLieDSaAubdQXGvdK5VoajDqtlJvQ8oPwpD7Vn5LjObuZAZ7viEOhY76y+GP04Sa7TA
8STCq86meWWrH5nULqvh4U874mU28CYtRcvICwhnxnogfDKlIZyNn26X4OJ4Cdxx9Ipu98PLlvCs
MvC6negtO6XW2Ig6Q/GrEGXumBZCgMuhesxRRpV+7hV1/cRzIhrZ1dfyKY+RGIL2Ba4uTEPcxK/v
L5E3w9ej6sOBTmDSvinkxuZUQh+hQXOjbJDNXy2cYqxFooegu8lijJFC0nkcH01SHzU3BtdRakjO
cYF4Dzsjp9kXcu+Y6ADDqO+m1ssqbdqOQAIEugMUYo5HVRKupKNoF63cahV397amT6cdPSlYkahm
JOi7yLr25N/G12dUAei+PmhEuYlbph1qWJ7g4l0QoVGycKM80uKauqml7iuXDV4uEGnT64asFzH/
NdLaFU5olw8psoRTX+cb8nPbiSeSUj9K+VMyajrQ8z4cWpyRrA1LbF8ulyQZqwmF00KJ6FftV3qT
OoOPK2fukyl6uEWFvfvB+1FTvhL5V03pRY7p1jKQdFQkbUSETwJoE7BNYnXzO1n/9gkfelvYWx94
L9VnMw+fcOi7XKg4vPgj/K8ATYue3ULQgRLavnfW6rqIP08FBy5Y5hXJEZd7iBVXRt7ERw8KJyPq
ugHgQNFvatKDG0dP3behSZSy8iK1FELcAvynni91XQBXHOYIsTG8RId/eBsRAATBAN2REcBQGPbE
zEKr12k4kLCP44IyIspzUS7pziI19eilnbo4cBzWOkmWRvQ4UkFiF9ySLW9MudujMwOB8FWf36cj
8zhh9XQimWwxOdPQzTqgi5aT97xesVILDJ6+/piQT42vZlSTMyfstnOZww9n3KyNDDku3c1XWUFl
NIeA8TAuh7kR4S6GQI7KC2zUXs81KcDMU6TmQj3nui/5PzFz+k7cd+UMIqPsUUv0lSZMFjvyoTal
sxQlN6cBc2Y3uVo8xmwWM3099ii3/DVKhUweXfsgo0u1QRZRoaB09vKO6BgdxEBgJInkcJAmZ9zO
fbpZLE54GiHtPN338R9J7pwSodY4xLMDNCQbWGCiCZwN6c0FFfLiexBp/BTEYcg2yZzb8nkQL0Nl
OqnYD79NUTFH0GFw66WTbZcwv5Bcwx+Rj4EGQggQ1VKNNInKmsWX3oWTolFZ15pQLOIh1jsISf+E
xwvK0am4mOqxZE5FIz5Dr5QE/QvnWCXTszQ7mvRPRJp3nFq72ByVgd4/1cZ15z6S7Y955njQijWW
dVHs5dQpqjGz8L4u+DRZyimGvRpfnCz+iswhjbUl1LRgoM+rjFtKBk8bEnanipXg9uvAHOz9Ac55
FHchrmEacwwI+VKTutzhE5/7ONkm+bi+OKObfxAlTq6AGM3iLIx4kigWyAJ8Nn+bzGU5o0LM6Bl+
E+gy1g1TgnfmkWFJKtFJ5GdMHe7OMHt1cigTYYK8KNKuEByz1mGlM12HQOysDHONW0QRmqcJReqU
BFGixAKfVRfCGFcaWYQpyhkjOCcoOvcxAmuw09Or73oFJ9108zjiQstyCJjY00qQYYtFyBK7BgMp
TC435CjkU50GqWFgnitJ5Uanvhn9OVScofb6Eq/M/+O6VQl675EU/uzSI8gY2Uut1qVw1N8FPSNg
0oqdFmeKY11wh6vZqWBzDfvT8GJiaTrUL3z2hsbb+36bmaGkeAyPZHlCeKNfx0kbCxp6T3dBoByx
EbBtadnrSshmoMrShmnCuNuRDbEFRrDcJKguRf4oN8xVJFpYLz49etaWC0KzSR45tKO7EeTASpU5
4myoX7uhgWeCw0VANSS2X9pndcskI8IjaJqvGz3n0nQXzp+9BAL131QjcrMjBqQUNxzzR339EI0K
W6ZQgXcLfcmtOLYMocNAJTwTCH0SyUpVX9uGtrVPaRidyG5MJCRXqlGTVgTdhG1zXxOj/JioVH+V
uvRtyUcqJsoqbW3xZqK3onUtz3EdVxqINaSWwmLT46/1mlYsXPYCRRdZKwEpkzH684lLOcKKnPPK
JXitWCkiaQy9zEnYlKBncJI4nsAUslNgNklOieLbjubJx/RWTTQnjom7pQaxJbj7auVPZdhmoTYH
xHJadL5gsyLlEZ6BcPXeDWy1GsWHRXA7XsyWR6l+duZZhoXtK+GUXC0ku1KeghYZR9UXKsFbHh3n
97n9FgveUwatn34bgtkes1m5Iz6fvZoJ7zyVxBUVXFLLpvRmAR0tEKIohW1tCVoM21/SLXSsAPyQ
dhwMBSqdBSsXuUA1tXjBZxs85w4omZpZKJP94fWXTarEvPwLPhgTvx0iJk8KFSVlbaOY0CQ3ZY2D
J4+jAjSb1vBdyIYFylbMVSGAjWYSeUWDg1aDCq1Dv+ufwx3KhPNIC2g1KyYqHSLMaMeV7Ccs9NY5
5ra1L4NyR/DHtcWliCJpI47g/JRH2hRlZVTUXLOfpZdgA8s4JpJlrZg6uoMofpyXyClqWHbPKhVz
NQ+0jXTHin5hx9an9m3hb1Cz5GKe7bDaS4pz+tOk3v1Tj72r11v9iIOwAaiIPMQngR3f4ZQJxW5k
/0aB163MYwLrsoKcUfYlaXly4gu0+3nyhsg4HI7h0tN0aMERG6josHILDXeiAz+7/ni7ZiYxMrLt
/I3UmT+KRXX1csJVOeNalvCSFEKirzk83HNHj4cOnNrZGI9Mdi+ER5xua1yMgOeXi7Jd9+zP4F7l
2FviLTsv31TsH9RyazmmBTqZzDGySRpMOOf0hsQ0Fk5tir32UEXbMLwjf20C1Q5AYdfs1Eeg6Rqo
FW0RzcnzH/ADeZctkS643fyeJdxa+/kU68FwQV2cK4vVtzGaC+T5rc7xj7u9OifIzorX2RTsy9Jw
acBZJEXEJSrXDBqVyJK9BjGOoZzwMQ/aSzmt3zez38h3hBXXj8dXSWWOotM4xOp8XYwr/CT0yOki
2kODZuzzoJ8/BJBsC4JBNwWSu3k0bmcdfJ0UFbVsmj8DrxlCogL8tpuzrjJ4MLbwOBWMxTW+Febk
wn+Tx37LQkwxT0vzfijkF4KDh7RiZ8PnCJR/38aI5pNFNN57K6z3ZrKk+8CeeOHcFc1XsK4A/BK0
NtmdvJddDFLvTC5pE3XNhAP+cExDlFvM6F/Juyf/yxpxuY4MIyx9qZ4ifq8aZn24lQqVnNQEtngz
igSbjZxSP+tInY0SnWnFwcoMnR7w91DAugJHL4873OB4cxnlfHQFb2dW6prFarvc1Gnb7A1rRSp5
BttcbWjWwim3wXd82ynWWa6nDEAP9ta3q2P/X2wfGMTCCkMdH6DM32CUMKo3xrn2CXT5OSTY/pJ/
YQ77sKlGGeczmuKMFvgey96xkW0y9RPvi953wcliaA4Hz0rs0kP3Hhb6b28IxlnFym9ER5hF9+tZ
0sHgxPQ8GFQxaqmJsc6krl7smmuGwkYmShIFc4np695TiVebiiyBU6y4RrzvrDDEtN0lgZuQUzlj
qvPjtlsjTEYPL6I0qPOn43d4uwCY0RNYx0mz88f0c6TCD9t+pjgFjTSJFcnIA4N+xZYm3SgT2qN3
cJaTjU3qKred2X9X3rb3tw8y3FPCs1KzJ6acMmvz+wS4TSeZP1AcJPnylvbaLMy6NJ1lrVKc6JZB
Nav4vJTHQa7iOaBvVTZoDAd3isYGVZ4QPMpXzY1wgaKDIabdq7jdaH6MYDxTo2thR6vE5O3zlRas
/VNek+wf68L3pZ2XU1L384BD7Fndub1SZ33/fMVaoSaxhvMeTcneWRV/opRsUzJ1xYVmniIGj3Yp
8TTZDZV+bsCx4bzlkHbpWMprhrIneUU7IpWkeFO7QIiIgxAAMVyxH/oSnXPfdh12uRRXe2i6pXS8
QWuYl5Qg2KZl72sBbsK7Dv629adQrRVFeXIh+FGIzGDC3SnfmeGFwfzudMHv0CD4kR2C/cHk8HRW
p0kwgWwUIBHwONb56Zvzxnx3/7peOS5uuCXWpHKWC4c4IRpNez0B7d6p/Qw+5rqn3JDc45B1HVuv
VmkXgod0gt48wp/TjpAnM4S8SrGO+ewV4/NuCjyRrJgZ6eccL0LGTrVuSakDKOEH+sdNDpisM9nG
ffCKLTnrnb455umXg89ntXbit+j/Yf/HPV4Pi//ujbwoxlztz3kHv3QbXGvlhl2nDr1nb5385oId
A+ws+8B5ovfNdH+xKOend+WpBGPSglpYuq8zonijj9wVLVYlyivear+CneaNBIu6yea6dyssP9kg
DkjqGW0Bb36VqYTHE0UWUbXXKYlK4Rs1rl6QmToQBgxv+/Pv8/WZohbAq1rKAdPAuQ3cgN25E2Fz
6oTJCaU1wrLLz9m0zcsthDZxAPabi/GVonLx2IOhSmyXEHScEEqO6QlbIzr+Y25Mpmwe8aYvJdoc
PJ1/xyZQJPlbPoduxYq9Iq7ZWrynk5OMx93OCvzFFs67qaAP4/cEVCQTZXKAoX3HvKH9K5As8jB8
Ky1c2gNetUHcyYsPZAPzGhIBJD8NdXMsjg1eEB69o2iM6HuilAL/G18dsDVGC1Mcx4BjQeIXF4ju
/A39qtzzAnHwsGTmlm5BilcUqJttgsoxnFq/fv4oWaV+pz0gGQith7EG6WwCSJZRzEqE8XI0WP5m
OUCYGi2HNhQMTINtFjzCxVmdxDyZG47nJsplpIAUzvlOp6w5aV2TysXcG4e6caqMht58/WqGeFht
p7WDvXlLjQ/Xj+srgIQBe6k2ZoC85eNRjsYkFrEXdsK33vJbOD3A3QxBUUpsDCNYLQr0X/MkUPkQ
t+Gzo98Z5Us9muilkC0tvE91s5vVql6QqiWoV9qES+4x2C6yGFK/nOq860IZNVax8FBOdmUGVCoM
HHxVinD73Erry8uOzWDUSNSUI+PJv8VALhZYrTvLmP9rxqiDOEFURHG/8wrCwxB5ve82t7tcQPQn
LaRdwVQ1BDiX+cQfgBEX53lOVA8aFE1y7xDz8G774r/A0g6iEl+Sd0nZWxa8ezJHe6RxVPda9sQ9
SAivn8fehk/EcDLMpUQVev2wCiLyweAQlewGaYN5YCiSk+0WEJoEQiaf3f2pjURT2BM2vHVY1xda
osLap/+tDOY2r8pkUr3v1Ybd0NUayHJ8XoXQoEG9G4pQEyf5XMqa3gtMBbgBe80IEm8y6Ubqwqhm
RFU1VluVbqTfiKUXQ+24DToGoJ8FxwQWR9tfUwTz+iV4nBrJraAbs/Ue5DjfXX9BldKqlXx8Z22k
k3YIomAeVxkVCftmBx+r7R/BpUHpPsTfSr6B6lBX8JZEoC24R81WwWjdxBZ5KNJV1tt7qPz23xOv
47Tz2a1spexZsSjAJRm3V+T8V0qiQkT8DDEGC0Pp8x+PoRJZ/AvTpIQ0j6dU8V2G7JUcLV6Mv1xp
gdoZMrom6sJT0anCCsSusk0wVyV7EW4nT8qLmyu7qkImQYcF4M/6CddoJXAeM4BHiyzqHc4uJeC/
3zd3UOFPyE2/jzXSqufwexzsYyVm4buoNd7tRUvfFlTlERxgDYZiEaaNjyZa49BKqeRn7u5peYpZ
OwTy3ihIj0wOdTCHhHVJmTEK1UrwJXKRf9yuqbv2MMUYoaltljbplvKD7MtBv/1o0fnbgW8AVCsJ
Jis7cY8bWIRxQjdegrrbkjWJZ7QadfpLEEe0fMdsWvMaeRk6rjdv7IsekE78S3siB6OTVS8cAUQg
FtZncpW3msSg7lwruBd9HwOU18xw5Mk/Tmo9919/hNtFT7AP6BNAOuSfwWU5IP7huVEAIC4Wj1Of
BYHZg/9G0FBfXQ6lqWp1+KrHr+F5dl31Ba+SvVcsYF3jhWUDJzIuwt7nkt4WiPEYoGu+EOHt4pVs
6DX5of9GtDq2hpNEC7LZDn70Ph9xsuH9JZ68tr8VvdudWN8M/vbjeRAHOifs7kAZI4snmd6aFwtU
VWE0+OVFg4bGuxIUBNXqei1gu/cR8Owxh6wMeXeUOzNv7fTRSYusGfYVdYWkIN5vo/dQYjUP221s
qpY4bEWI1F8sjvgvABmFtHQbCDvW58zdOcUCggHezGhtMB6YIGN98kgK7nSAzH1EphDs0HHyR0fA
KaM8sEvoTJQbJmCNIOUIpjEFMBbJEAp4lygvxVHxDlK/sRWcmpzg9crYLwjNVNG3dag7Wa446t0g
nLqfvrWW1O4llpn7FI1EzQh2oQDR3IgEHc9C8KCWPXBSvUvC4cKlQSETvdZbR3roONzEQDj692jw
4GZlUN21mgz+oMI1DYAIsWb1MhtbBBCL9/fRum+++qVLIrsTqfIHoYlOVXamutZXnl2a0jZQgTQx
GguLwKqRRtoaCzdEJTHgvN2i2S8/1kpuu5ZIhBQnSczfQB4LZ6BSD8AXQLE7iRZbDYqoSL2HSrCE
FElk2AECW6BpJklZydYwfkilFGI22+j3rRnaSPT+nbrmVlLNOTfrc4qGIA0AAUVflfBAdXljkXli
HRCaHJMwJLn7NjTdeLha3HeOfD5dZyV1iqmToiXlJyMK8hEbk9xN3cLKBv9zl6eFtw2cK2gcyuaW
nwegzY4Zosr7J6LXG2H5dA1+lgKQKn7IahYfCSPfamH3fvzAhNwoWjbKclxMBcbUs1bo7XWmz5r4
mxnBbNwZ0rpTapWWPxaN6HQRPwaXzWLs48OxUzOoGTuqliVMr//2msuczihd0Q4aCOXLMlNSyE8r
pAT/mVBs24ZP37CDEEd9c+nh9yXl03ujJM836okYp9nDm2fgEw+NbG08YjRmyebihjSE2l7wcvAK
K5gxMzG99IrPy/IuAJy7H3ffmHs+JoM35EVwboZYeTYbXTCnHWVMCZIr90hj+NVbPpxU7mmDez2h
TQL1Gt62Nux4TyPokDx4jYe3VjID1bKh8pn/71FoRD7fSnbKcqB1USiAZfFwpy1+QURMr4LjbmY8
AP15OOdVVdwWkM6gtTP6QmayIEP/5HlDvwq5AANcnqJ6T2e7acDi6cOvTejEHOwPFCI2gl7/qfiM
4T4sCB5PwtOKH/rtFpBziTycK6NeRnVQV/cTiZqmyr+ikm68RQRKKKSb78UjDbH9wcpvtIqtLe2d
38hq02tBpjhbgJTd1aY7PpSRq5nGexNYk1p/xuF1ha8zP7lcgkoSyPHtjMxJbtF/NiebLxMnNuxg
FRRHNddzcrbyVodTZjIK/TD0z26DaciaBeqBI5YLkca6GPLiZn69gLEoqr/Fw1If1lRpqIoiiLEu
sr2iTH544yqyws3P81HSnaVWI1CNC/BmPJGTIVvOoIwY1xHfYF4oY965BtETYKO+fK/JrRlUBeOS
GIr43GiwjabLWRfo1T1lnVrm25FPqhI3RZlEyt2FNOsMhUqk+5LAQ0/aw4hvUibm/60qZfceTbaM
05r2pfLrnzmkywhIuJmfS8+nIr1zmNgnkHtc3fE0NYt0YxZI34b7P79tdr6EjLKQwwBhR1t66DVI
pGiI6Xcs63k8UBLRgF0jIQctEYT30IulCud8a/x0/OYYso/ldjSBskD9dgZYUGB8xWa8tbdwdZRG
xuee7lU3RVBhf8DOx7XkwD0amI5hi5R3Ribwg5B9lWy8ntC3hIxC72vpbJmWvEQelMb9Gkr5Omoo
F7FRkrw0lr4OcxGZQ79r8Wsbx9BKgFuciQK9HsiPGka/3uDdlzuRXy9uYhb3ivYXloDQzgxLG99Z
cGNdqOQfO5GeDNX2hqacas3WDC1R8QJCVvhrJ9FEEULsaaI1TaqbJjJtDzpTz2jrlcqk97ZiHj/9
2oqx0jD29ajuR/rATHFgNNayqHPurhZPrABuLK/HpGkf8haMGBA1lru2DHR/EdFLvXhFZbCr8f9K
Pw7cvdwWiZJbN5g2ibxWtvcgOfC7vgkvZFu+UfKE+MRZvthEiVsTUO2kLBhiaWzGMNIbcavtZNPT
7itBYnc7hq2KtqR84l/qMN2LpyiA+Q+saU9iYRPmICOt+S9ZR9RJ58hip0pS8aqmq4eyOm+qxqTI
FIwVgbE/uquBJ65bC3GWCpT0D61umYJp+dqIfl6FGgpcXjSwGmQgagJlszTYWthVTd9D6a4jHARP
bKV6F+DkeVc1sqQg2SfLUIswEbM+LyW9sfEIjb835f+USWr1IoSYqpNlxc0BbFHrfoTraMq316C4
XcgQ9+7A7tdWc7viwon+Bb4eyP/h1UAohXZPrR3jo3t2/L01KfsUA9dMuYLUfL6wmNAvkFf14tev
Di3Wzk95veSn/HGcKVFt7kAqdwKjO25Id2rhiVf6kXBsS0sxeNSXudadEO/0B1ks+lISTZicO+CR
Mx3XhGzl7vzQFtWkSwjriGO3YpBulF3w9Pujt/Psir2isgzH0pVRGpdNXSSCPWbM2UdXhho7K0Lp
ftQ6OeEaoPkm2BiO4GXTeKKxkBYAtuFZAKh/1ySTSDy51wwBSt6Eq/+Xn+7PU/FVzoCB1pLWTZKP
TbGdMgjUCRUJqc4FpUY2t4Z6MRaFLCgIuF4pd0CwwY0sRb6w5URNw9EEmScFowpJYSRyzbSQ8UcX
w8Nkv25aRM7OzBPfwWLZz/E60Q+nAsZ5oiTryzazSZa0ykHH6dR55x7V57zqddjxUt64ByvelFc1
lrd8Qgz4lPL9q+Ku3+0F0i6alEkTok8aFavjKafEjjXZxff/oipQ362FL415DrLAWrYPgUGS0Mva
HenFUeJUVkwW+iJb9ehag/JYyNj8m3Tif2w6cOJK0MjX6BbfDplKwGfl9e50Sr6vFHLlT+t5j4DX
Aqh53AzUjLC4NvJYs/gy2Q/yrjEaiEG/5HAh7IaJ9qEf4tsX7wbk6qQnMxNAGpJwTO5AVKcgEBQb
8Me30wel9+Us84x0TShtVCoKoA135BY6JXvD+wsTE9eZufCew8bSagQL0r24NlAb355GW/BFhdeR
oGZrWWZTEhg3PzDsFRREOJX5R1GsRb4vXTeyjk7f717cmEeuINVTKGmQo1ZDlapp7Ym4xh12qNIB
vwVd+01B/VojRVlvusecO1BeFjwgLpjG/6ipNvydS8YI6nTJKXQOFnQ6gGwnppwstkBa+xpQyat4
W6i1P/rs7AUFxEKD/tBxgIEE/d67m92SxxJReMA5taeTKWH+7jhCq4sUbJZ+ArMOEmsPsCZWkn2X
RfC5t2w1GJpIpG42WxjWzFKEtmzTa7Cd+VjUWmDZcB59UMwh1qFPHdJw7Get9yAuQ6meyc1rplPu
kl5Es7wnsg6YbHzVVAPLsUdKwi7HwT/hU5ZFHmG/hGserPTJJOszJ0AnoRF6ges8u9jte07b//Vl
IvXVYqsB9czKTTVTz6q/ayaVVPwBElfklLqsIAwG06ocL6wMS+ex38Py+V6TXEoxR8xMCCWPAcYz
ynm5eu8tyy0bprdXQopXL+4Hlqdsi49U4zlrJ2YVpEqJoRZgyKuuOpxdeNGBxI1JSCBCR7Wn7F1f
qhrNCcaf9N86XzdVs3jL7V2BLsGbM35BWiyQo9Dwm9omlQ0ytpodc3kv41X9reMuTLKDqiU+zRIa
8C2UdCzjMJySLy7Buc7mD4+oBb2xVRo702g/C/m5WtE03+L1PZowKGi3brscvDjsZpZbWBQ6u8c7
Fkl8OKMBBDBK5CO8/VFG0/jdpKdQf6zw4CFRqxEVIqYfwy9zy04fbtm1stmzpduZJtHCITbfTw2R
GNvXaacKWhgHjy/07Tk2YAbM9Q3d3FFjmN1iPtrcgpsCq3Ziy8Ke8fKohzQJgsJOAVTT0p7EssfH
l73ae2BN6g8+GGI76GfAY8LAwkljwzVBOv/5TdP9Az8dp3VboeP2tMXdlubqBzWftwy4JJoAHxP8
byb1vlay+WTgNGroZ13qrm4LE90vgzlouVtMbicFOLktHE/gsbJBMGapzREuq5t6/n+o9GVaXwo7
BSTO/29CoMqPou5JW2j8Y0cBL8unTojC6db7SbdjxYuXv3lCCO37FSSrf+a+WA2UXVKzllMcXxod
YLC9nbkt0R7ud2XoWdH1Dyg+uy7ACi++RtJLAy4+LtSuJgRQfln+iuLzqBWNLg9SStju8lbVJvHn
G9dVWjjexD498DDY+WdtS3S4XvLsA1b97FHQVFYHfdwZgvQT28vZ29oXC08Honp1eDfkTtWl9/lJ
yGBqgpsLiTySWceMzxYkgyTZ0ZFjGbVnbw12TtohYpSw3JqqS0c9FanV8Urbcx3tr2knAWUQmPFk
YbbYINaaX8VT3Ll0FC6iBJcTSRMUwmniy3T2+0hW0ckExMb8yPyel78eN2ywfmw1yG05rRYQ1Es5
mxboHeZu6aHb/oj7MlM3hL091v46hNfq//D2RX+TtjwvxjFZw6Sow3CUIExNh5BlcmIFy5wzrhEh
HQbH/lzCEnCED28pIHQ1uAnmDqXaSwOCrvvkrYAMZT9O0oXQxCLRFezqB765zZbWyI/EknPkNRif
KTJ1T+ZjRwwUsXIYM+3wlV6AKsfZdogU76LwKYr8VI+8ZoPyA7dsx9SI+3H2rDrNra0a9aOwCoc8
+TwLrcK0df4dHYNLZM/iZE70FbvIXxTAy6bI/3KsOgjaBhwY15ocPas5tbKhEW4vm2IiGnF10mAi
/9vlJlzVcF5oJvYko+E/rgsz0YHEBOsw5VYqVDdZJDfljSZ9heX2ygZuSdhJQyDe9jBqOi54n2Qg
dWgRXcIzxMqLHVuYWTsHpyqC2+/NCHv5QCkUT8iHGM7LypyDcfW2vcHUzxO989lnrg0GMPxGuC3r
Z3Wim/5LLUp9zv/0PTgo1QRUwkt4jwl+ApRbRN+UGXfbz9xu0bxXX3lIGKS1Mthd9jj/0QdhLHXz
Mrc4AoHfiWS1bFOCccgTvA3J2LIAGNzx3FfSIGny+3QBgg2KTsfRlT8D3F1P38KJLbIuctPK3YSg
yMMeaZOpc8ufn3JwEhLe4qEYg7HcecC2szyi4GnA65ZHBkWiHQE4lnvaw/D4uaKHEcmaJU/42oDw
TXgWhVkZ0NYbfv5+K0+CmxzJhLP63r5WrK4DWYDvjuMKJ2P7wJvQxn2c6Pv9b8dKteSydSnGNu9+
lqil+2MRnpEmJy+5By6fqWkQOQ4/0kYEK+tKn3UsSqR+H0D+Lnd2H22QJVJ/F5hir0kWInjQTelg
iBpiNRlKlAA67o6wGGaYqiggb9VLANcsqi7q/nHhSbu4mSMpm7AI67qjbCEz2lsvWPNmhNCbTsGz
TT3vXfeKtw38Ugt1Kbv4rLsWxY3H82826YumOoMB+8BbRV9R6ZKZsf8nkDbgInQsKOTSTLgjuiFP
OaUC65K6Spokl/CzB7CNZsj6V/dXHMjkEIYALtZ86SFSMyUajuqLC684s2UX153dUq+mSIv/hLYT
VH8yaTgBgH5nUaxTJ3WHcvEghvWoa2MBiyn4hNZTvWDtkSPJxsclaMHzVrI+1rUKg+szObzjQ77w
wPWTbztOBVis30CBsq6z8LilLnX0ajgxq4UBiL/HIkkHoL+WIkf1Z65d6XDitro+TWstMY9S5RtJ
MEqXzICcdlusMy6jJ9u5M7IZpxyBpB6Q2RTq7T1Nl23TezqYOOwdF9P5QkOxkxvDQ3i1DtpkfIrH
9qa1S1qISJpLfxKLi8F0OoB9CsVTVvCQJBT8cMtKEYHs8UBew55moaCX/8XWejm1R5wg/7uu5D1E
2nKlazwGqzrVSwcP64XOHVUadnSUFpRhaNWfaJ2xSWZ/Ckz6tX8jpPkKovC0kUXs/lnlrWKOsVSP
Lg+osNWTl+lNvQBlTvYXHjkc6jMc4A/X6fP6dlMVbtXjS0pZxpfC39dTbwBegIYNYCLTY5ETl4qf
IMsYAkbNBtRFDtmsq7I3zmUAZSy8aVyLHT5mugSdbE84edk4nWxEcR5BzyfzMwaqVLBDIVVutarg
5lyVGpw0Ykg7DLFnGX+f2/Buu/AyY63psWsC3KqBU5uvHHpiam2BcOs5o4xhfiorKhZ6c3GAiSVL
cTS+1IkBvDLZHzIMv1BGH3CUDHb0O78/iYaRwCvm+pP7K/Y6QalXGfPkqwH1aUo4KDLeYxSVE2ds
K0tuNwzL6JaGAfRZWTv7ZIBf9GH145mzWfkR/03RxIahIL/LN65Tss88RFeMULWObQYpKIokLn9u
PR4g81mT/ERYizSGsfmlhzqIJU1qAlGzO3/A2mZF1an6uEw5Bprs/7BBXi2dw1iuGxIBY17PJkMT
kLBydCaY5dh8EQOWQRgTmPzu83+jWX+JKbwRbvsTbC9o7KkJ87b/kQh7DGXRFT7HtGyeTL3tLW3V
nN1NzWesRfQHzJV9aozspL1Sg7smdQ1KsKZSoGzAHD9/EnWn/HOatp7CZZju0cUuliSEcFCPqLj8
0r8GfLMMTxpu/33K4R8GuoBIYJqzQV1dJtPCWBNfhUKJEyyJ3CtsDIYmJD8aqTtycyB/XkKwhWcv
UJ8kB9P1n3F3UIRI0TF7IYrWnLklGKJlGxz8Xq6g9WBO9ZlfeVXVGdbqhRxtdhXwK2vGocCJURIQ
kM1KTolhcnKwFMEWOFlRnJ+UDkzusG0n1FnIewJohbcaB7vsOZAWeKeT4DF/8AThWSncqwm1uaM9
U3JbaAyKHC/ABTV9oMSTS2NqfVezL4zNmNjoLYkhUF804cOt1VW2lTp8AdT8y8OSHyq1+YSEIsWG
zOcLq+qPyVO8LORtgKvm575AgSEx7YjmofVxYNaNOlkAhlJFomUowSIh7K21hbTj6KpIgHytKiRd
AGNSVQzs/lqQOkpjCDiAwRcpYPwdgWdP0WjoQ2XzL4gv9I0JgnCj2J/8VnqY1jqeGLxeu0hNbRDf
+jtNNo1jKmYncKrmei2KeDiOqcmdThwgykUeviHiQe0hP0YHXjL2IIbLsTXkkm9QAJp8SNG4eGkj
OSNBw4FTmmcNr+shOJ0xxgFkZFv0TYj59hPuY1/AAGGLyI/Hq/0cgc5NRQEztxgQTK5YAl+zcrHq
8EFZD0GyhMD6fygGmSjxOrgG89lCP2CsVhZ4NT8twEzUB+dA0yPlDJssj3VZmxzHVCU0OXGG/Egc
uu+WEtG1gIL6BmRnUBva23COw0UPIFyYApdOicFBP4dpLL8nmGE9yA9AJqvUapqQK9wQR6pX37sS
YPIZdGRU2sVGSXii7I9a0mSC6u7gW2c41RcG07z7PfbAciAw1pO8/6i/MEF0TZL0Spc4v5NrNV/Z
BH4JtaZH+OENxGskuNaeENjkV8lJxvQIyGJPZuUSLVDLwvnt0mOYLctte8+XjCkqVdYqQInBybq7
UaYIzMjoaC5XyLL7z+rk7ssrEzuEC5W3OhItLOJFCGyhWgSXXc5HItM+ePvLF2zeAo7z3cx2Aylr
/QLkEKZSDduv5zbQvp07S56Q3R2Jo2cRhvZBwEqOyshZVVIfgXQN8mpTVDZDvNMIdBqDfis6uBvZ
YA4x7l1Z3P7pm6mlmdUY2DbMOuiH8liH9Jo13yy9F6jFSnP4xuy5OPCgMHWQlPuQMx1B3rEHULud
ld1UxOQ/QaMp4VT2x02TVsyjNIAuUDzQCBBDlJmmhsFRwKT7TR0o1tg/dIhnMy+MmgZd63QKD4NS
jxZUl1vyRl1wHlh5uDIoTZZkot9EYbWWNQSxyZXwvWSpYuKNDM7LuPecmXqvpduw55IGMB3EUAT2
RpRGwmgw85IlPyuZVUkbqb7iHZ8E9FLud+3zjJB0QtLH+VgoSXLN27x/ElvFRvj3hjejrg1pXxGz
mVFhbhpZ64qoUu3OvsT2qH8oy1XIC2kd4n71hDXovsno3gvPfJLMZGa5Rk/3BKldas1LCuafLCPT
0lQgaWtmw2US2ov5O6fZonRdEk3dlFZX4Y9TNk1rT5BE1Ti/Z1tvDD9q3f6ojV8xk7y1Hs7ddC96
mPJX3IHMsV6Xm1FlJ/qzcIh33o8cLiL7ztPwydO+cNuncorKMZkPjsT7T4iWQembMH/Gf1hTKgyr
KCrhAlusxFN861/xK66E13JbGMjalrPExH/ipOXDCp5MaWgsHq8kVYPQ+2uzZ+1GfKoR+Axj4S0F
QSr7rCaJEEdXmTKo+uGxMNcyJRh6t5td8yyW9+YAJ411NtsrHomF0tRQsUa7fnOaXZry0vLMeTny
+m2UXposn5PTycDWDjdTy/cTfUpojUip4vZ/6CiLFYhiF49qub9kocBj6IN72GxQHeWRCyeCcXTr
qZwj9jNZph3LibvFGjDddKc29bEbfY73LIn2nGB0mb8yy6WG35OAK47ZYctT111UGdY7+pnZ2JGZ
1LZgAFAueNZepyVBRxGpSTua2+Ai2AglpeL79BDPEc79LmsxJQraRJKUirHsE01dHDCvH/tXACQK
6ZcaOIcdhg395UuN4NFNTOXa3bDUl4Lx3ZwxU1GwhuJ2p5zmYp2Qfkx1ZgNkBXms4lQ7IuxYCb0K
E0QwULubwuTMQbqM6sPOMwq3zCnTVgLb16xWMl2v6KrfGzLSiS2W8BKxA1W8ya77zcfN527fiTTb
N8lIAGwFaAbocgh49+kO/izkemOOhks7GkyqpRYHRKZFuObZeMFxB0bkEkW+E0Vl4g01jajVpjlc
D0FMsn7Uano8kQW+pqMeZ7w7CO8rkjzjg33JSTMnKtPZ+USd1obBE9mJYSINh7EJjGHGug/TkS6c
2XsI5RmqffA/+P2beYvNdAI+bjDwq2aFs7BGlg8smsnockCmvDsCLFiunVjgXn8iWgV5O7uI6fSc
/OyYqiaA/q5L24TZGMk0gCfVvvzw02Zo0idvXNZSdxvci2M8d+cHmmH/J+o+gY9azgJsXUqhsYu0
sExFAEnAS9/Pl/3xVYN+GF0VxZQRzgqsX9PMx/fh6LAQX1sQCeEp5Ygi+kTG4Rb2QX66GKtCDz1L
fDKZ0PeaZo9oQSZvjYp4pIfY+soOxn7YxtrGF51YSwk4xvc4ddn75tf1bla2d2Zeq+GDwCLcKiUt
FtAfe9tgxLjxgwp9mNqIGK5JQ5FAnnWg/Pd/yDX4AfxZqvtJmLkgvISUov3s2H7c7CH9HKBETc6q
bTntt5CucJJ7O/fhvwWH1+tWa7cIT6WsibQ6H0jOFGvgoEYgodHayk7HLbGU4jzM4kZ9IooOJTjx
H0zRDvu+4cjPQws7a9B2axBXS0sYboAT37WUOqJslYMafmIOnB0WCrzllGONYUP3dsLWHarom0zW
JJW80+d5KhysHBJfYoHuPeIx41X5IkJ8I2adbhlQYkP8qxMi4LSGCAGjNcazzwgD+IQHoFfBtEQW
2y5OGjpnsOnnWTWoBqesqvJ3IXIQe1uAh6oGzg5qVU+AqXN/vtH9GaL6tOaMEf/PJLqCfQva8IF8
VvLrCPiq8EbaLABgoQ3emeOsTHiNkVB3ugOwKJQimeQwxrQge3Gu1+I+4j6DKsc3ITz3uRNdwO5k
cnoL6Ika1ywMgxJRqvGGTpXQKRT8HNXxF47AI03c+jWM0bgKs+hlvQiUY+EhVmkVCjRT5durV7pB
GnB+HVev0N9sIP0aG1F6uf5nyoJ2VpJ6w5R1uUYeHqerd4B0ifWHsNzODAk7xp7BI/cd/y2p5M+x
dgKSWZnPOLvyHb+i9sgBQ6xBLZfnVefPuP6fUTgMP6eS3EPSIqJjuA2l5O38EIzGI36o3iSMBM44
k44CuAsEGJPuJS382Rdt93mF1yHIcxAXwHHYhnl7Cp34fySwN4ZI2O8VJ/le+JcsHVwb8bcKtQuf
cbSGeRDhqx8IsF5g2qmpnsU5NShAnNyH4ucqlkQr3t0UUg9Q82/fhGwb9Ex6q6DAQbu/1g3tFXec
PGRBxCgaHOANH/SfLmwyx67v/KvJcRxs9JUsDoN9PgWHo6t9YaI6hGIprvPC/NS/imDWopYzG1zO
J45ClKqr/xeQjD6PJrtbb0rwcw2vorrWga+2kYm6BZ8uiNbWm70CHtLawu7sJP4XT9JnXgrfCCBz
q96qrrvySMMXCaQGC/ed4nG/aqKWHPamC1T0nTtsEANIt3zyEHMu9gV60kq+8qa25EBuEtd5AXFN
0D2B6K/muE71Rf7M8b4IkT+hg0Zjm3lDDzdSb7aziXyC2ixGk8b6JBTpkH/8awqIfm1aU9ZlihNj
APCabtu6B4BmaPmdBHNoQJglmf8jqb1fv5mm+yiVbDCEwL02Jk07PXCqpo6y63bJe7L9uNCHWZqP
R4XW+s8ra57tA3QygzbPuDC6K3XTIIcvURI/begi1OAIPXeRRT9rOoj8rfP1dESlElrbIfAWbnUp
TgAciSr2dCoO+Ndw4wuOP/YghrJ7GZBKjiqIR6hNHhYQGF7cHyOdXB0bk6K9I98xoE5k/Nyblk9E
ikIfAXSZacadtPHTclFZs1/oTZyIyRuJbbNP6V9vbouROvTIom6gCpE2R+VaSHZ7BrTLOB0Q0VCF
mr6ShQ4QDjmQ7EOTdETPb6D4NFajE5nUwpvs5HVxWkZOnibPoc+sNLVfm+6Maqn98QU59bD075zA
x49XsU/Rg5Wsl7sEmqMEPSUUDi/YW0/MOfuyFV+2gOu0FIxf7V/DCMZFogWoO/RxelHwDvUqsz7q
j42mSntiyG88YynsTAoU/PWvHn0C8RpKSyp9mJacFfF7x+PU9eITVJqWy1k5KFcuwvcFxGD4yNnV
275qcTDdOo6jcoOgpG6BT2wVVyfuPIF2h0L3PhIrl6wLQPNn7Nu7EUqzVAWxry4RL/NHenN2+3Ms
9ipz7SHWmNCqdD886c9yF1xAg0w7I+/JbeHT2ebVqK4QDjLZPVI8yUAagNu+ENU4lKjw59Mb0OYH
9mzpzOgADp0RKKItjgpBQi/iij4AodjlRRVhoPaoRWKmT/T/2I3h19uG5VUj+0sk5rK7dj+HNKVp
6K7xiqSrqFSoX5ODm4LMvhw85E655S0nLhMxz6z2sV+Bs8A5uAflxLadgONCvjclZINJ6hQuDP0E
TTcB2U3DFspZIA8JA24XoTZco4P2lqaVPWvGkEj3nzniGCOn3+zxYiGE+Jyi9MvbVNLC0Jh28dIV
TPzMYGV28+l3maQN1a0xa8HRnrZc+IHrmTtk8Rs8TPQFq4jW5CJWhiibmVqFGsVx+MomuaHvYMxG
CoqjCSWLZkUOmnml9NfWOnNfglMvC1YxBE+OkxObQqR1WQJFeu5ozVvP4oi4saUvoaG07RzZboy4
+p23tz0NU/IV31YEqWvdk5kCXpc1EM42UpfHiu5pfmOb6/YJHdeDVpeQ9EXipiNZx1GPWA/L3RiM
5gIYVwPehBRSlKwjI+3K7BbSemACOJUpG7x26Iod692k9Ntfs94BlWNJQVwBl6CphMIF08lFn76r
v9ESwNgSELtnEgMZiIp06S2SDmIGTFggXX6mDYIb4Wtncv457PvBLxm1DBZadQKEqzd3PYUNl+bc
77vsenZ6aW5Rvb4GV2/qPgU2Ls6c5VZWAG+nu3aVndSVNKPDXB1413+QjNeHGNexAr9cLVleP2Hn
snlTUTVoBWAUXIJ9MHcysPe/xDNigHTQsMyXlDiwcStJNIVuqjGYcVJlKS2689p0upBywpatPwH1
kCEm5WsbOZogCDo1MsemF9FsFzxx7KJ4ih2XfUAnpkt9zWr2WUsfhDu4lFETq/janfXov59J4MC4
htrvYar/dhdrUFxTmEBuvt8NQ2WjZJeHw8HdBphaQnm3BBkOBdBsRiREkMhrD7BIB3LcTIhIH6Hf
MKmEdLQ8kNjcGeBS/fZ/YyHQIeDuV9Egfy7p/tcftGSIhc9kHYdf0XfQX6qGZ/GFVyM3rjHpLlJq
1Hz4gZwOsJQB1yskYnZ0NNrT2SicbfH30Sb5E3whKUtNS5R/nFdGhg6f/Ok9r3pZfh8QyntVyGTI
7wywOLtmyWTxEi1Jh4nCsTn2ahhaTzQlklKuztAjCMbhImgDZsRlR4Yg8ULYPJgH5oRKWoel6oc3
KpIpg8kDXSs2KwxiVGA52sM7ITUQ8Yj9e1H4SfRW5/uj75FBQr0Wr9FezLoHQOIbZwJl7VhpgkW4
eT+6Co0bTJKc37RSv8Xgei7LCgrNbhy6O9peV2NGhDkpeF3VK40Hnl5u3BN8lUq3dqQw19mQaws9
7kU5SESrCu5r6GTChiHShBiQNiSvXeoQSFe/2shvNfdFn8o+ofNEkSyZldG90ykWT2f1FRhd5As7
b7gPMx4jlcgPZp7cQeotp+kRQQtRD1oO/UWDYJUh8w5Wv2LBI1HhaG22CjEnflaRZCba+MtS783v
cpoqv17zfD29coe2u6hDhMyjpdvt1Csk0OhzpEtMAipH45nIBGrNClIfvfP5vEFxjcbIMV3ajXbz
f6OSpBKH3ydRCClllm2sk8cvn6uVe/mKMcp9dbzdB/tfpE0fR/BAJpBrYfJ4SjkrzCHLQ9FlLxXs
kc1VPMICbrIQUO7q4u80HSGTsHvUc+dIOZlJ+MF+uPURA372IIG44hLR1FF4QqFBXz2NptiPuUtf
vOYT1VfqXy5RskwsZcd9SDnKgY/hYKzE2nZWLXwMFBtTwYxBtZx1+8vQulUpDMyVEEBCq3YaBbUO
tBd7oxxxSieGxWp8Fux1IBcsOFnYb7SarPw+YxqQsODh1UmqzFbpKfxpXapHkta0zNfN7pueCwzu
87k0Fl6Y9SN8MVw0sWQ2qmzXaS+4WYUyYPwk/ptz/FwvWj/QSGXfKD1KhuWGsgwTfVVLO4sWx25o
m8t74hoW3nEwQWvz1//XvbJLFzOBR69gwh/jrrfiLfogVpW9oCXgTdRDikbGerjO1KTgP2nDWxUp
xshEUCDo3xEdyeLZ8nX7W6Py9KEv0d7POLvYedIfO41ht7VgjPuL3NG7v7pJNzDmQdhqH+Fw5+Vs
B0MSj6gq3B2ydPoXJJ+K1jEtOwKq6/SfG+xsqsFSyJ6eYWMBefSzN0RTLdvfJYmCyMjoTxPhKao0
dGJrqS8iFj+PbhwP9GK20jeN8FdGCbAHFfRPACQ4gpz4pZP5+vK1bMcyqXvGMeT82IAFdlnyCdVT
+ZkQdfTPvw2gOBqC3gmNXNTWZ1Oro5Y9WIb6cjGL/7S+yVQRSlEU+iGq1qb6Z6r7BluGmh1p9j4k
6DYx7wwGnPgVPQTcHO3aUy0awWv/7zGRx1tpegMPat3Jkojgqx/3vpsJmBoVu7IO267owCIDh59B
YLwB72VNC0flg1FJMmcM9fC+VE9S7EixpcsFtv4Ee5wtTL9ixLhS7ienHZX5OVSnIh4P1maFEBlC
gM7BMZ0FdTYaSYA0/aitdBKTShNMFr9rn4bZCbiSylYffHUF6TLslubOQHURYaVnkfdejrrJraQJ
FRLDZ91r3FjVu4CF1YRbp1oKfK4urY0+Z3+yGsntfMct/an360nVeEtV+gnHZJuuosrerYLM7DXq
FzxhWxr+vEKvd36/XrjOgvwIa2gjsUM6909XliO1q5j6VvvvfV5b9ZutV8rQ3RlKxKZ+9HZfEQfl
uK//ivq0sFfYJ8uloB0Yk2L2A2X0WYrPUpwkEbXe8zk17jBlq/Z1c5h8z2bPTc2+bgXLHgWiOXLl
YSbuAc1D9jAJ77mAW1Eh+BXZJoQl0ngyW8D+RA612A/ibXMZWktggn1Leb1fQwpkDMIviHWt5hw6
BVWZpet0+iYxrcOJYRTflbVbaxDEhKCTf2qHMdRCXL7w4MmLnveeANoqmi5NG2VwQoxTeDxJN+vy
2R1mjtQ4bFj74mHBdjSM3w45JIypUGFzw3cI+CMewiB7OYhWTnb2tYVizuT72QnkOmIk/7dOJxHT
M3gAlh12KV3YRFz5HSNEdGiipF7vtJVrRmDs+4R5t3ngUSFldow9jq/yV2YKD2SEQVcr1YVYR52F
HOC4oayKaRSePze2J/sGIzHxlxNNjZhmR+4Truf32EmH4OhGI2Kyysnd24wh6QvCvzQzw/BIJH24
r12Watlb7WOXaOXIzQx76d6Kst+aFu9M40B/fpKXnM2NmbUqZky1A/lvJXmEK6Pie+k20KasXjqx
xQjPzpDtp1INQtrja5gZgW3td+kvL68vT6gk8uZ2R2aQSQXXgOFQ8PSspaBNM9uEzAovlNAIejNT
SUczjqmH4M587IiRJVDJs8yrrP6YTKewMnSfa+ng6TNUKViKgQ2UAQKwV86DackGJYvourmnCAlQ
KQFQ3cUayBPhTL4qA2rWPTAHfyRzKEdLwsev3NiFfC/i6e+9e35q2N8RjlcpNp318Cdqgg76caIf
FJJWC0V9A8hijYch0URow9RY7Xwg8AS7TZbj0RWXVRnKownydNMoi17cAjR27Oxs7Ng5Ei099hvm
R3eH42h0paMCwRox573JCMdmQQf6rQWD0zaFG4Gm1MLCjveH7t/2X0S00LCbcaUlr/LdYlmwgPag
PcnOeGdRc4J04Dmzv2yylvKCuIGRML6D8EXC31ms6INqgT1Hdpy5F8a04zF/Al55J4sKJ4U68P0B
mMGe1K/Aw8N9vUJH7aUjN14HpcrFo9ffoBDCtXOEhW4OYqm/ePqHe4er9bpvqaxOM6EqsocscoZj
sOxLU07QXvp2ouQuPxlDSETCt5Qf6O20z+/saA+FYZ84mKLoCEeGXuXA9bJJmmBMRilAUBeEwA7C
47lKYHnKHvglUlgdKrLDWlocAcNOJFe3Y6QLVveyTm9JhjjXUfBnlymEdtB857EDu5xx4uKe7wE5
2USwNvlSYPD6FWW5NMVfhGz4hharGL/ftdeXub2xOTBNoFacOZ2aWiT6xD8NSJ1sFaVlg/TzwjAV
IGG404jvIoZNLS5m+I94CgLU9gC67HV5l4SFvge/ntywcPsHQIVbtmdVnr3en3J+U8NRxJSmC0nz
+N8NvneP6WSduwY+gsSNfy1E6AM/ByjyVt4XQ7xpmdvu1DYueo18cDWtgBh3rupPyLa2CM5KaSoE
YsURQMs3Mud2duIBw++oEm1yBZ+S47QUsGpA93TjdBzQzCc40u56FJStBuAIpepHXZQN0/vhXH9Z
d1g7UJLZXj96ufLpCHlX7Do97VIP2j+677MOXBwOxZxSN79Or6NGT3XJGPgsvBYGrIx8tMxx8mbI
bPi7IWXfPro3fj4YkhPmvsV2XrPoLnDMs02slQSWeBjLr086X4QbLN3TfQmDrangxjLl0Ve8TkCB
6SDlUMuvRpCcAtM0wiCQLfEypZ3UzB1lapJhaEWTyR2I48j+whlq+omLHqsM7f3mRD3w3haKd4de
ESxayw4bHqMXiJOU523cvb1p0TUz2radN+HOkhkGubnP1VxG8IYoWUNSwTDwfULgM4wXJvJFLocx
1Wqzrld5VUh2rwOXYO8PsA5UIrITYUDFFConcS3N5xdXqlcqCKcj5kDSTjfNFIIcgXdRWnOlJ5FO
b3Xc6UBeItKSkrHb8INDt8inXIAAK/GOgU+v4FtHqrXx1B+JLGwd8nf4PksSB//GbMe2RDjFLW9C
K6bdu5UWZZUFKgCopbzvmB+wiWXFtNB/LPJt4jS4QY+zGUPEf+RYXxGAp5d2byreaZp/bCE4fEqB
goCKIAUpLmmlhwEfuwqJQBc2qegGxUNPa5I4XO64itP2Hg08eaTqIC69ECUhRqji1IWrXcPVxU0o
d4I9B9UC9phgEZUt05L+HLUKv1YyAXxMknUyni1y/CQQtFn8D44RIaAm7HjJQmzb1KDWJcw7Ukan
OaOAYS9FmQ2eVeH+fYdoQppWLt4ezhS6esPS6xgq7w4hN925XEbuaH86ZYVXJB0IBd3mQ/J8X5nJ
9hvjQTaitKUwFgb1HOuETJM4EE4+2N17fP968Ni2RENl+4oId95cwLKJ1MKh5Po4r7/EJeZlWi+K
tfokQgPif1SswWB+o/m+dX98S1Q9SQe+wYLLP4NAx8wlR6j3Jv3pn3TPYJKu5mB6TYpen2a+dWvp
qiTILQFYf65xof+eff+zPAI8hDfQq1GlsXoINsAGzE7kzZZ2MHB8tnyjuBUAN+wUdbkwI5rdjAAi
U+R+opFxYr9uWN5oYX3KYf5xG41RK8h5kmmtPr5K49ynUcYV25B8vJw4/4pVWHIORAZOCaWvW9yY
f+w4w/arWZ8mCqT3TrUG51inq5x8vDutBR1qv2brB2x3jVWqY/ZotnnZk7wyEeeN3difNSh0W3e6
iG8pt13WMB5K4kVmRZT80ka+25u6fNl8oMushyLg7fQ3LSZ35Vy98XFSs+dNDly2kyUAg6Id70sc
19QZBle5X358se5ULfF/OnNRL7pCX4rq9wwU57xB3kAPrx6Dp7H36WT+CDkMMxl0D+e5bbSdwJl/
KtdecTeV9T3MyBT7FgckIFGd44uUBhm+4sztel/OuHZdx0QRIGr+aYXKbWKR2qsEfEmq6W89POY9
M7BYkkhJjB8TLeSOwCkAQtyJGcFKqKoE20kqgrjUmZiOheptL8T9eMnhBnAA7qwLhF5LE39VPvC9
W9yS0DG5okeKiagOlkl3kctpV2VjboNg9TCKc5IcDkh9q7RkqFdKsPgB6q42Vwg356cAM1VwWUHc
qqVHd1jRXEnxZivkaNDbbG7iJovvnOlwi8jdlv+VTbRPFTkrhOuKumdbouhN6kwiC9ruZbAcDDG8
FTI7Tug7REW5cO0y8H5a9bXNwn2+q76tcQ6ik/hzJ5YMf3Lys3p1Ylj7sGAJQQKULsxHsvQDRA96
6J8Zo7QArWC/Y5QeBCfp9kcewgOwA66i5yrdpmlGln6t8jKwF1VN5OyeQl54rXXcntohyV2bmCwC
XLXLL2G3SPAo2d5bidNB8DN5lCISlng/PSiofuZCTIRT2rDv/A6Fwb5S+EjlWaOl/2+QRc49H+Ro
IR+A7CRoormxKQi37ID359Q/fRwm/cAscE/Cx/ECZTpEaKUkadM/UEtW6ysRM4h7niu4W6J6Z6wB
DhH+vCYjsaLN5hTV5VYlw4Xrc4ND6pNPBfnrax8ryx+9ohePPMIMjqRAXK2sBZ3JCkjdzwgPEst9
odB6t+8LBjJWuiefcSF1c//0XvDdeFsXnEU9pAt8qhvSzgN1CMjDKTzPLxZAqjDGhI5H9MI7TZas
I5ZLhdRZdk1nDCUBr8d4XqRqHkVqmIayPUL2pgWm3lLjYFWtRbD1ITmNXS4NTlYrH+DREdohZGip
x4mMEpK9NAXztBWnliAUiw7PtI3TxMCKlnGXlAqO104xtqzLXjic9+A0dRyXmxrHkMNBS4qZYya0
bIBhs+c/jNmepEBNcpb9SGBHw0rceKLkpfWA28IjLlNVyuN47qlPBdKvoIuRbxaa0DGGOyS3+dIV
l+/tsK3k55yUy3O0p/n44VA4RLW8EHX1DXFZXWa+o55GqpgmDOTzg4q8wk50NQg1C5HiQZZ2KHrH
wL/C9GdmPGUqMT/WibJtEG3ItiXHHXP3VNA6O/whBMUHVldIi2uHTLi2dlhysL1P81UQt0wITjiN
EkA+wogaBJreAA85nzL/oHNRIK9xN8DH84f86CGsI6krbnt9mw71zskKYthO6Izrq6MdRp83G7nT
7gF3AvpV+y+Vp7Au5aFNC1f5JjACIYIbSOHKHJfezGqTMBWj5RqJMZhBVb4105dTxrx1eya2Eg0x
o23fowjpeKIaqSF+sP/D8iygU4bwOAVsjAKM/wyrWLwwm2yqUFXDlOkUzMOhV2ffjaKQ3qO3kOPj
3NpRdQnWdR2UgOkcXyizoN7rrsbrMdMxMzDd+2dopN20+JTwqctmsrWxbb22PsXQ4MUuCS4Vbm/2
P9zZcTNsFB1XuC9TO5wwLFgnt9fSKVBufgeiiHSimO47UOpVhEqktuGIrYzv6u1f4tidoCZKUAaH
IIPZJYdnnJuEuDPrB5uAxX/AjGB1ane6CG25iaJjtxA2xH/RlBq3sDFKYInvYCTUVmJ9/UQbFAg9
nGOxZ2bgWBRxcmTxfZtE8XeVhdxqY5Wa5iSXIem4MqPhECwbI0ra+vqhtXkTCsDvhNgWKQlwrtfF
ClsacE3Fdo0TZ/XpuuD8FccSrAPR3Ab/HYzBvs5Fh4k3DdMCG4c9HV0JqvfqPduUkavB5+19pRE7
l8vzjTUNqjJT8cYNSDgLMSLbzDaNOb7g1MabdLpew92j5eher7L5lnJaeDqpRRJGHWCrbBL4TLLN
qtXnIm4N3W6kFpPQVANwF0p+oZ/7Kyjga6BmMzYyKgSy9W06geuEeb/dp1Vcb0Lg9JTcVMYsDcDV
78YIMGWqmndCTEdUKTQ/BZfOB1qqg7Pg2aRT4cJMguG764HeiNWJm6aTw6KJ2dqE4Q/xrAKnzJMQ
jLQhXSvOW8I5BjdDNdQmnuV0GGkx/urk72EZvsVVYN39WeqYLLs5jhOVymkVz2QsghmXcCuPVEaC
Avral2VRgN6YZWiJ02c5Pt34KQRcC3AFuuFBE5eZe/gfDT99k9bg/+1Sb1SqXpqOnVzfyt5aa3Ka
kcO0caRWjug4zqUrWtgLb34Ty3Us9/KgVgUAlsOFfH0qEHopth3WqF8w4yUt2SDbB//p1U1X/wNB
mHNDQCf8KbhWNzpzekp0na+XgIUSi/xYAad49N7afdPSwgEBasjkJWcU0xM4+UthwrLHuunMGF9p
OsggfsD45bcR+cOQZPFQGCQ8SiZpC30fg3nkFTyZhN2xcQehGT1XtyMI52G1dBF7C5O2HUjac7UH
snDjlUP/PZt0ghpiVep6xPuqmbij8PLPKD9xPoNpQz/IQVXJDlcLOxHSi/RXdvXxy9IgdA2bcN/Y
T8tIssHTRTp/DmV/Ri1Zy5fIYSiXs/qoI98yTsYQObMZwnxKJfwaUgUn6H+OhCXRHszYPfxtO4jh
EEvVOOUf47v2GKIVqE76Gs+1fzjdYAaMCThuLlqYzDRwBEQszP6Dt92+udr1oLX0YrwTgJZ+S2d4
h2Rw6ZdVxJPe0XIwy4dBRfxJmEJRNiYwIZ5ABVNwiusciCgxnm74LGl7z7oi8lq0w0ktPDKjpSAn
Zbb2YVRfbXTT/rTtRFwI7IF/chCxaLiBs3CTtQBZDsT2vLOdmTzWc/9Mlj+JKzJMACyj1CthDeHw
ZNWHV1n27W7GE8nvS/QyH6xB59NwAOKqyXGZhhQEHDljk3CMVqJEkt4WsMHZugXy79cRrVJZXmgc
NlbkMkS6o/+0omUBYNbZFBT3OJmJoGoCn1EPoMqxf28BCM8YqYGITqOPMEy+8A4eAczCuNUO4QzP
Cb8B5oSx/qwFbLVzDtiEQsJzoZS0MWapPC1ek+8NPqU9q0zXmzo/ddXRSF42g/ni+lHtNSrbAEjF
O/5S1AK7b6w6xoZRkvrrk82hnN3xUQ4PH13rT8ZaLo8sXQoeM57D3vR1c9Kz2+K1JB+EQZ6zUJbd
7VF7iajJGSYsTHP97XMmxcQeX1n6PxfsY7UX5Ty1ZKCOsl5XYMCDlZCNIimNPCTYVOYAD34G3AoA
sAR4+6InHTP3XWnNMoQbYO+1oiO2NZoJr1m7IXIDMalw3N5dGHfMNA4ZXbkgXPqPK0m8Z3wij7ub
Va2W9Sz/rlaltsyMm1SfHrRoLhHdICMubIZl16UM7IuWR16Kz7S8lMIHCoJ1SlSe8z6gaP+g6nTD
5Ign4ZdoNesxDRtywDZNEPYorFp70BXj9mDFfg6ssZAd4FjO3E0b7ZtKh6NPw3Ec2eexUsYNEG5j
JRuoyIS1vdIndsPNLnDarBo48FXZtKpOy5sXoGIQAtP4279lupLCucgD+YG33WtSebMIKqc9L3Y/
2wXLhk9psFx+4G9pki4bryu3iWD4XCEXu5HKox655Bsvk41LYOXy/y+b8X8wN5RdaK7MUSPAgaGL
UC0q+mPrMGgy4QFApGdU57Ck8Mqg49GKhrwKeUp190elFigzzz+rEtsNfXnMT8q5J4dKpLAznyvJ
/ITxZBDasdLCEhEzkSoo/itrIYNWKCxjdZSheswSsfFk2+Jbvthu4QzxkCFsv4IUlmFbI6K6x9w9
uDyS6bWqFA+3Yc1/vmBDUnm5miQRo8m/bqtCFvKTElFm5/HGR1jMVuL42n7GJxN8Gotm/5wochfh
pdzQapwv5qt5Wdha+HkUaYbSD1tdFK96lzs3cM13JQF0Zv0k3xEYDUEu/dPkc6ewMGEmI2PzkG5f
X84sERCZZb587ON2DJFuRU1j8MOHmVzA4OcDSrilKeses2LnSFXoFHB3DRwikW7V6d16U+7+ujJR
4RKLqbppJXeZqkw4lUYKDFSS2nPkts/jzLvMz7wJtinzIVUemKKvlUAqtfp7omcKFk7zycZtjjKd
cHsf8BQI9hldkkqerdYqHFqVa8QgsXP007bhveS0PQhCHVd1bCCYh1Bo5QjjtXmIs3TACjAEaduk
8b5mwXeFGFtt9mK92B1ST3fO26GN2Up07iiiHLfm51mfd0my8OiqZ4B1mn0ncKCEpAotEm8sfmo5
XJ4YZgKY0TQF5jldPAH4DWftmX7BRa2paSi+tYV03afh8pOVvFiJIo48HFE1atgdJiv50l5CR+x7
svy5v29GlmCaOvyu3wfRziYZCp+nxDC13rxtpwjojt8+I35JvQTs5Orv36OLefZ/jL/qymheUy5I
nbyl985JydNiUEY7mE3R/NcOWszoG51Adyah4xmutoCboVeO1gcZnbBRKQfauGP5RafaUNdgew+B
cv4p67H2oC0+G2v/j021TPPvAXg3RQmTu5W0fOIRGlLiuKjd7+GqIEQ2uShtv74EEZAOwMVc50L+
T04B5dg5W6TEFxhmP/Tguu14vz/lu3UQ42+MjT5YKh/1itaO5eQFiPdGannfTGcQqPTFqSmhO25I
ZNa0dhtqSuKBN0YYPm4X1UDefw8OtdxIcaqxpFpGMnRuLenGtwPmuBDdvkBvYbhLUqksZ9TtBcxZ
iWtmN05iQxUDWzuDbGKt3ic1dAFfXqwQheCUUyjmD5BrDWStrW2FuFsXv9DDELW9AP8zWle6p0Cs
F0e5Zhtbj2ZCVyg42sv6OlaaLt0KsI37nJOafl9QY48Ak/Gws/3wfdKGcFwO7wGsE0sOBmfHRxNd
rJ01+XzlvEwzwA1G7G41OHbKAL9sthm6JWfflH5FR22YGAhVHd0nBgpsN6z2cC/DB3X6bHPq1Yc2
lJIykWUjkMBIIEuSGi9VZZYKrrwB9hm/jY6xHoTFJK7eBbWRdFvcSwNSfEDI9LE0AHu+mTsSRFiZ
WAp33fLPt6OP/iS4WhYqAvFRZqc7hsi9+jg+mnxrRpMuphG8hXz2Oet0IXoDMamHUmZ8yqIQLSUf
dUZo4B4LVhyM9bsLdTX93nk7A/fvXv1YesNIJ4bQuPvBJs022OdwcIlkd04b+WYN8AnP0wcFJ+be
YRzXQ5rmVWe9HZoAOelsvQESrBVjAdOjKYTZM8a26Mtl/f7HK5aKh1Tx/8kK0Lm6hlOgL9fvpgH1
lQvg33ibmimiay39gfEfF3kjt2LaQHUhVQ/s6shKO8HC3RpwC8b35IRAQVqAA8qdei84vKF5aPl1
xm3pnKlhPi8XeXsZYptrI4KWXNMiESPVArt74kE8zZuctDRHnU+dGt/SWaexDh/VTHqmWqJGlhnq
E5JwsWkJIdEnx2FzrxAHEnk1NPNihZxjxNxSgYszVW/1529rpeRRGRZRkN45gLc2lVT+rM1Ynedn
yrzJH2v37xQskTexuC4/rwQU6DEKeIe3UZiwT3tJAE/G0DnO4k8+O4iIRtV6SYg2+u/r9LapoxmA
nRO1S9+MKFgBMLeLNRujHYtFio1xjyNr5AZc7MjHIY3xpLiYvfvXFbI8dl812LSnAnLvVYumEaWg
w6WEps0TFBnov/OfFWQ1NBRThSGngL5jPsSfzFLESBeo2RFmFXqG0R2S9Ul2au310rfGbh6vJiJp
n53jBcQ9j3pXgOv3HFyMJtJmwI4XQeMrW19Klst9jVgnzsy+7BoXwKPy5PnzaBPtB7QCueW4UPXX
DMVRghTrnUqNR6gK3YOqQnOw6DKZwgSkU/xZbJpQkS9osSe+3sOZnBr52kP7cUXVoJ16TZlsw/0x
Jk7xwD5soTcvNPgw8Ttbi32CBAQv2LtXR/gQqPv4Ksx6WMjFaZ83SAfuOm3TDZBDJIPJRJyAuy40
g8enEnCQrcFWNGavbgfyjZ4XRHxgGP0yR06rVLpUYtKMGfGEM0XBCYxRKeM5+K51IRwGmEyzybC+
cfohXkYcsloIYzP7pv5Z8RNnEqvhEuUdMBCmmvywwRnYL46Tkzvxat9yWSREvDjIPoKXegFoQFPP
uRYb+aCk/KYwFENPhBi7yTipqSsmpJOqGTrxaV3rN7qABUs46soV5B1KBuke6CPad58V1BRDUUhh
K0/mqPT4ceneOypNXCWUq/b6lLrAxZNy0S3qBNu+h/GEJppGEC4Kc7MyqZzriSLbMmjX4Dbw6CTV
a8hwkbtKZcWFsYqJQfbam8x+5d4Or8VZLc+dnlBpfWSGjsDBgwVuwWIug7S6ZE6ITmhvJAbgUSV8
qxX21ke7Rk0avoLDDPzSW/eUuqRS/LBfp31r31bbM66KTk9Y3loo3dL7CWw13JIpcBqVBVih5xcL
taDHhFBBGINgdMb6UKIJVmy6D+bsFMooarSn6SGyRbsSYAR9QbSd39sjHPA4G/oRYK1lXmHBpoVV
owkBfipmqpPisVNo9+HhuWZ/VaOHIQsVCzvEFxnlsgVIXqSqtVbxXiApY+3djr4eUZ1JMcSBFgE3
pnYUC+Qux2bOAnfPqnF0KRBn/BnPHZt7efqi0uUowAwyTiQOgUUe+bubF6WL081Sz4DZ6TdYdvrB
IenM5CeNcflx/cJ9mBURvrOkuBrkhu1p2naV9y1PhfhqVJydS4UexH25YU54U1+fM/0TfcTVOc4S
ruz3VO2VMzJTkzb/N8s8xhlMmW/P7sa83XrDc0ZXmztz7jkvBlzTqtQwFZab/Vf6RooNqf93FmCd
3zbNsylmOuHeIrB7fCzz+UhJ2POyNTPkKcCKymzVDu7iIgZoR9s96Eij80N2U605+bSjEHSPYrXv
hjg2E3asE9uq/zYhTThkPghWnnH482tRBNVxuN67NkIbxNrlFnxZfSwY749leY6mb0D0lKPosFDt
Zl307Sfv804rTKIJksGV6v/JNdATP0GiNmcHAnI9n0nAvmKwhDmiW0ePK8qsxWjf1I4tLZR+Yotz
3zqtW+TYURelpLKMEUMrmK7uFkLQWCvql+TAzqnVpmlia0W0t+h5V/fzmGDuloqONj0ovenoeyzZ
iaYYkJfT32VAFM9sCTQGgGJmayzexV4MODQqwNWkmtIO6xajkp6alF+rRM9EzpnqEbd/E9hijKvz
1xv0b7fRnWJkGOkJfvX7Lw0cXpgTdTyNQFggh2RRufpuwdJS6cOmQbWQIXAz6e33O1qKMq5hoTlv
7CVtQn6yd8tq38D4T8SN/8paPeTgMYYlAMAI6knyyBVPpErd/EnpT89rlNbE1RnQve+cFlH9A5gY
kNcKxKF9eWxKQvTqMkYcAjuxLMl6qweVeG29Pdv0fyDHxeDtVsCxHaiAtTLKQdARsEF4iNFNTEY5
NhdacmTM4KY/T08/pqX7qtw6Yy2O0AP5mveCbY68GRHOY9+loBgzlJgauaFuRGpqy+Uss2yXOYTC
64D06uhRUkSarlNM3S7QVT55QGUQ2mNpVJ83QGM1rHybLKGBDiAkKUY2zB1G9vddXW+qpQNzINBs
ZvOWxozNZfp4BficKt3N1qlwvphkpx4tFYdkoBMGMRVmrnFeJK/uz73uYnqiifN34xc8hU7dd34l
3M2YwLYqL37LAi87GwQ22t/CWM64D9+d3g0OqiR1RtQNy4JXKn0caGVQxShI4yxthV3RDjtZ2mag
aEE05qe2y2w6UwwNWvxS63R+BAmtPRj7IRZ2SKiK7Vq29sWfPQYVQtUuBbGd7wdY2gtt4yh06Ky4
r2PuMxQlGvLwGPCHDBnLIcURWwUOdWsHO3CA0Zcj/2pPnl7poqvU0DjndQEZR4c5Fg/LxTbzqlfS
r4bezoyECJxANdzBl679HLX8MvCZTXDWtfAtreT/FF2vEaN3dEvrDc1+OW8J22+Y/fVJCSJ/ao9F
71BbgdqslbpUpHhCgFSkGTWjKFAbu2EDmUTuY76z2juyWKoucTbRYFIltxjRyjbaGO021leoQqO1
3taCihxHmjIQFN+Jm8r3fEWLiiJPIflkmdGo1Cc+kJsXdo+l8n35SUujUnHkkBSmvwMjmSyjhJvQ
IbLkt2hfkB29nN/SalTDQFmW8yhgKaAh7IuMBa+pbmaeryrTRQKMQrOvwiqDGNAUyKGTCiWv1AGK
aY5YZnHv/weIBFz7FFb0QHuT5JXuhO/1Au9o36eLeIew+ga2OJgmLOBlwEnwSq+TsKE3toQtRULy
Ku3e4U1TKOpIL+B2BJ6KLPZGaREEItlqfLl4LJhOQztOS/EwGeV2OehnPa6Tbf/rByIBwILetGow
m7ZoWCoL0jgz5DWz390u1wqbZ8vbpeFoBCsrYdti8wHNEmlwZqWZeQK0WUDvLq4NTauxW7U80HEA
d9dbiKC7PdXEv2UVZqKnNJILHuTGJx++B2YknPmQieTxKe1dLKjgrD9zLY5+C3ZsIaJdNrablztm
ZCm3GE1AMaqzHtUXAylawIVmixK6vHd4ziPhzsxon1XZOxlWKOh4hOHqyFkmfC3dv2Allqnsrmk8
tx7lFVQflsG7BrG+3A8KqfjBr6R7zT3zVJmkoRrlPpcES1CrWRKlHePQRzOnaz81x25GsI6L2IT/
ZURDD/su/uOlO4eawRJqGBUv89IlErbJ0fXUioDgkMsV+Z1UtSUJxmy8kLm7yWoidDqhMJ5+CRtt
RvM4ovE+SpJ7PO+zNDOfWEFks+rIAYxEi7a1ZEjWzxI7bTz9fc3k726BVVdJ/DAEUii4mViM596D
51Gonm2uD86jqQFQko6Dni3pLETL5t87lTQ6qXCcpR2VTvvjQ7CCTg+qQm0GR4W6PNcdNNtExk/H
CJO1DyPk0wGj6d4gSympKNRmdfR999INzGQ1ciZIOanMR1AFYKdNKOc8nOf6v5zr3ZBPAxhbn3Pb
IT4wKLF/wGUpW8sZBYOnWmGCTPfyAN9tQA0BFXrwam3TZKiULV/UCIQzilWc6G/DWGtBvjJkCf+O
e8aa9guPwenfXvzTdrUsE+g9FCJfXLnr28qXGNeCoog9EkYW5W5Nd8+1EmkQxkzrE+mY1+t+6W+5
4wvswFCj4notnDzzvkQCZsqiIv4Uv3Una0brOnqZEDjb5uOtgOPveb/WlaMi2lCIBuG5B4egsyaU
Ly8vFYovqw8tyjZOSXOxAudr8mGPPI71JrWKPVuFMNKBwcJly4W3Eo6KQffdcEMxfjwXKDNTJbSW
GQXmu+XYFeoxZFvcw+BJCgwssUkYroqbh0MhPKP4Qao+sbqU3myVuyytIT3sI5EA3kOy5k3JkWdD
Q9BLT4k7ta/wnw/Z00y+kJMbpEwiGIDUsK++a3GMC6V8Pm8wTY5VJqBZ2M7/9AcEFXns3Bgz4HeK
iCOME1Rn4+3pQHtnPUFJlOHR9t20Byeu7sZ5UyqpDSv82UtwCoKDAgGBPDTEwxRCSORZcTM7VtNE
pkJP4tAd5inuobuVKfjcqZrepESe5s5w5Ho9DMqLeTaAOr4gVELjpUc24NorpqN/mQNc6h7LxI9H
R3OhrMOjt7gUufW8wrkqIWiperEuMmDaJG5BUA0uMd5vHqhjypqoAbVj4VKiYLs/F4SL8Yym3Rwd
k6c/Js+2ePCZk/WcbZs3GwDqq52+H31Oe/z4tem3rd1Q0UWwJJ4Hlgz2GZPipiQ7n1MhD+96GrY+
AE4fVQG8AbY8Mw0Op9xBwP8UQ1E9I+ToT+wIx9QYjXeEOwkFMa+HZxPp9cme37h0Yl5jZhWeY+ns
/sMvBJS2Q6iz5VJVK/CDhO14GztrJ4guyz6KZmNOMU8XQ9mZiTCgKBWEQV2SXF9MlWfvbf+gw5JG
7RRC5Vk9Uo0d13rU51Lfx3J6WbWLdFGnhy7RLgnNexK9UGhqIdlxP3yq/KobdMVCmvUvvp27SpW9
ptZUAks6IId34RoyoKZBYq3rgdTgkmT9a5E8QioyAwDBR9tKLk6ujPHU0tNj7/Fs2zjc9nHttoZ2
SKB1WwzmP0ubNEW20KzmrpXT5x7oi3WM8ynBJcOvE3VB+c+QpDi0S9RBjE8kzvv4XVOQuAMr/iqh
AY/pc3ZIn8Zd2OYRReAMslBTYphKhCo1lffPyIM8fnaBTEZphts+KtH4AM4iIbp+el1Y4MrnN2tp
3bSjBpEQXqDUwzI4O4/3UIdbbpvOuVyxN4tbFK9Mjuh+dyIkmJbll6zVqA4oAXKQuwPobJqKD9Z/
GlLB+5iv8GSYJYV/qcVKy1TZghP/1W5c01XFvXJ97A/Loah9xtPckBs0aehxajwOPMltZNwlgQFG
evVfOHppele+o1vfS15J3SRuWb5Q0IUNu8DZibRDGE56BXpxReOcNJ2R1CYl77uX0/EHsPsmDclm
RIFFknhjDy9UXv0tN5ZNxqxBNyvV9RpnCBtBir9nkgPmC2CzeQFjfEbDvJo6Jc5pU9p4UCLiPhyp
6lb/+YHzUJNohW0jP+aM2lnuAynzTCBFO9mykuZiLk/kYP3xYnwQL9AzNR+Pn+h593eTPmefvVYU
jniG2UNtbBtIsaOzDd+G/QpnQr13EG5oTjASI5c5EJ1uwpJh5ET9qOJCU++jr3qVbKGmaFN7ayhx
T0gmnTiTvfaYilJP/UMmHON97HjdIaydUWBYDnqdS8B5Ga9yZVwrrLdezvBsKw6xQYc6MWMFI35w
pJ7wLzNRLy+SJ/ura0DjzzO2rkSGPNRw0OPTgKfhxXlPV4GEhKjIomNWBIDlMzQUsbtoBEIfcpJe
bt+A1oK6W+5JasW7cznW7Q/8dbfnZ/lTHkhIILHNwOdbP0LqB4TOAAd0fXsVf6FK+lW0jks4JstF
pu9+635odsfTRgnQK+dAsA5CMyYQNvflXPCAWeMg+fr0NkM9X4KISVhXjVMn4YeCN6GNZSbtxqFs
W3apFb29FScSHFugGBo9zDYmJl6K+S9lhjyppOovGvxAdLOvqGhNSufvqKnP1zJTlGF1DBNQEveE
g3HgMfQ718guMYy9I6JzByubHGM3soQ7qkmz4Tbmjs0VmWTpp9Z5OBevnoAlMwIOCVNpNnHSd79D
43mBwXTu6l2VQvtq+Dz+uM0NMHk9D1HbrCiSCnhOupOpvNhd5WjGfyyouZbNDRO9EHToT/v2e8Go
DecuCKKXquucEKRG4nAy1dEMLE87c5QkK8i36PFslsQyhLmrmxyWQssSfI4OoWZwNa9mw3J/rBGP
q0EaiKAi/9OFR+3y7a6nMi64D9cmrcmep9nyLioVpg4wHVujUGTfUvlGnAlTBoEX2Wm7+5B5jLO5
mLnnXU4OwQee8PZxA7K/WT5IS4q6V21/l8NfqkodnfN6e9p2ZKjuqZa8SOHXbk/1NG/2QjZ8+o45
qjKlvNRjs0Nk7mUndJRxkMfgJ1Q9VC+GOju8DJVOSbZq2i4Nj4kAwHlL55FKPp+F4OBbDl8ghB9O
UXGD9PHjjyEi48fMFqLSb7KcEy8wxJw7riCCRvuOmDrpNtUd791L01srVzyiPGpPDWctHsYOC88R
RgtL00VVPqJqWDbltZJvZytC5fbKFfXfNr8Bsw5F7sfMkyPPR6wgOd7YVTu5NvugNUMDla41F4+h
cjVZU9qU4qSSGfGSU+N6o/zbGfx+FGM0/XEPuClatcs8hdjjz2K1gpymkETO3u0C6kTuftR5DN63
mpK2HHy8/GUBNsAySTA8/2KAX564rq9sGmjGwUcwBGvuyJbV+EYnhsxajWGu2U0lkLeh7Pg/LMOa
kNpbM4huzzK2obEus0PDEg0Q6PUPClm9fgrfI9qO9+C9U8TIZ9F5L40XSliqr21Vz0O6ZKE3NISJ
c8iw3vVGm4MoYmHQ4br1DBnlXQ8a+zo25VX+Q3L1DjvQkmTzWvp4kZjsgH7K0bAyJ6sgrm/gnsnf
tRvZoJSxgaIx7dYhPHacGsyYdJqIeZ8ZImLH8IyYO2TM8APFOnw3XxKYPOgTTPaCe3rNghcIRxze
fw0OOMduBWAZ6H6AdXWjHl+kZKGzkG/R4DKex88TTqBCcsh36q8/dA4sjn7o6BqIG3t54goMKJnR
0hb/nmB/Rn7f9Lh1GogZ545EsF9Uk9Tf8IoPbSicAhrxrn58GUoFSuGovZrl5xoYYd3vLjD92xwk
aRYqQAByjbtO7L6m1Cfauz0G3EG6izXsjiDyzLbxcYzBe5AMMMUezCMnNw9VQOt6xnpnf1IFmT1w
V0ESA1TmvpMBlZycPaOqFSiPTF6FdDVXrriGtSIeJDLknc9bhgwGZXYvx/TT3E1T+q26wpKGv6mu
g3F7x/c4jwvPc8YVFLAVxZC8hNKmOfbxs3kE6Qg4a0sLbVKPuJPfzjMaLH+t7E+Dx0YRs9+PIVXJ
M+JtXOo5HrrflGc0wjbtGlVwlA7Bj2+NCAZrY+JcVQp9rp0o4yAoIBHJ+sten4KyL8vszUtQLv6p
IV87861wY3li4NxUKa6FI1nO6ME9flbRFBdg1Xwvz39HwYuyqeeeeLhzGQOFKQAbhbFeP6zbqOSu
9R4aK9mAxpvV8nWja231Gf5UENzvHAC/+5S9bwRqIk2tJgmTEWqjFX2RFJoGJ4sszlitDj1wHiFW
5I92eHx5n+6TglxASsMUo5e07A9Uvk+4u/Pv/a41A7dBDoSv8OYmxgy2eSysvTPOkt/ZH/8MnSDg
5qfoQ1XC+ZDP9+KF0Aw1bSkQr815QzqJzmguc9500kMowKdzwZIl2yMy0GSNaEh6fTbF/vot9ofw
naY0MnqVdTZYW5TJz2O9/J/+8LUb8X97BiLTbMKk5WA5AFSqPQbAbtbRfDftVWgc6ro6Lm4izsen
w1KLgf6rYukSqgAw2QkZrxLELOyAd3v1dVCzoNCJoqLUJ578hxqOnrV7FGU2l0QjjrSorZpvWmvi
oZKAp/9gMkFlTpnnkd8vY7wV8T2CKhWLkjiI4pxelEhGH3T837YD/0/HcQl+T3da7Cyf+/3VNqsl
gy+QhwsdKGqEkDRNW7eDz1+cL9K24ljkW9Qb7dTrbkdIUJI265pyD1KuqwJoU+xoUfUKBl61fsOR
l1PyIF/duT0bc9Pf/PvLydcZd+9Crl4lsZMfdmKdSPzLqXEdlfqY2qiruY1F7XW45ZpUIo+50waJ
YQYaBAF8D+xj6xcqpWdZAFVpyRjoKyWdlczAjVCQCAZ2UffWZ7W9ouKO0YtpTDKAJuVbNhqZk30g
3l89b8dgnNxo7TSAf8pVSamqKurXnydg8aVbExGxvXnkF87FHBo5Q7MS+kCprq0cpGbrcbkjsGTt
3VgXImljYyW4hmVKlK5OR5LzD+0QhXEL/XQ/+37Bc2fSEOirvGM7qmjDcskxwNsxxIRHIPM8QfBa
5HTLKrLBJyud1e8eCnjxwEtHCcgjeXvu+Fadbd+kbytfO6YIIWuNfYzencdy+lc0l9WJrs8kCIJg
yb9S/oG0VYeVS149l67AUX4rEgTV2SdnkD/K8IZ+5yFdEbtdHMEzCND7ix/RPsc0+kZmAzN2WzZf
8Z2OgNvIrurPp/fA1ydHYnnCON5+8dA0ZTf3S3frvMrxRIkLF5qbvikod1J4rHoliFXifr54Lk1o
AYfK/uDRbn9n568jCKoQip8qEcZNpfR/npYxc4gtTqaH6WwjYclQxOpBXaSyW4ua6oQMmO3o6eQe
dfhmZka6gKEHobpgM0aCf/iu8mNaHQrHPmuXhCUYpIHSNmxgXiyiEoVC8Ua5nd/947Wiy4PeWo+W
nBxHTOPS0oDWJaqgqgv1z+x0lY9r0T2VKVpKNeoa5hM/6B+JtKwanPehr+w80btxkpn1MiYy4vZ3
FeagSHmqMMWdCLXAfFxOAadGpU0NPB7IZe1uKoVjJ5mnY9z82RnkTJCQWvu09gqa3I6uczF4yp3e
eKlIP9BhwZ9oQeld6zx1Nw7HnaA1CHlSK4hEsiUUiEn8zqyrwUKsokL3J8OqRmQStF2+BmyJ+Rfx
gjA3B9MK5TkTsE9RXvaSV7IFUWez/oaubsgiTUv5hB865oefNYwk5puw/jmwWsGfAg08h+8rSQNR
INp2XcUz86WHRCfW/Ps0GNGHxuo7vyjoLKOUfa/OS4dHzlRnwBEse3WqMK3eIrW66Z5PzD7mT+kO
gTf7URM4WNSjnGpdNvtUuKOuOl2eJOD9i9b4vhuEfVmt9pi5QUqPH/aQmUkYikdlb9zrstFouooL
YfVMqnLqYfz3AT/nZQoilKyYhOUofgkVO4DNuTB/PglvLUThTcxXWjeTXXmcQak1G5tSBZRnjSvV
TzC1eeAJk/coPP2M1ecwvpmXoR78LrCEsV5+XfDM5KYyDMOSqocHMFgNsiPfFWgsvmABbu8w5omH
UgHO7StOS6IXndwO4swuGjaDZOKMScaTCHrmgQPgXcEsc9DupxPmfC8XD5E7FyBBVqokIFjZq+pG
DbSym4Dza4zOpqMZnZ6m9Jw1T4WBE+6uMswwHjtaQmXTiSGFfAhnaRaMeWI/dbRehj2iDJembjj3
wJ6eyYmqXAH2HT7XEbAM1lEoZGpT/SQsmCvyPrFqdPX3qG75UD9YyzwS4cWXfIeWTEtbemItanjI
3QgKX3AyEZBZRMMQSTe1YR2dXT1vWqSgkWbfA5Q/qyYCIizKTu8LiDlH8rfmoYxJ8U7DcJQ+F3UM
qFjZh28YbrK5zVAvVjrl/Rk71L3uL7kKQ5xDn/0GFXSWruuRN/8LKc18A9fPV4bglktfRxXUSUpa
dWzM3zqYebE1FN1esgeSdWrDPUv7uk34q6Osd7AC6k31NNjho+3qbmkeQJydaMAOjBk2wR7HiALF
wDoStTkA+zVA3tOBw78uXHZADrVaWDmEBKFAKatlrSH0FmGlrweeZC7k5N8DQ4rMrhSHfeRO2q18
wi/KH+frFT+DYDKo28JqUyY91QpO1MdNaarfShMKn+VZ8c6ywHy/uiIG14HD1MszPVbBqs5RiSJ1
ieix+gG4HabfXHe4j0yhd86JGVz9lJ63LeQGYH7QxHhfgFZlDjiE3MmLBipuyh9B3ziAJ1IT5kMV
XJk5UM6bmNuojbK3Pcpif1a06msaWmdV+TfVi6XpQgsYtayq1ABd4MlLSmx8asyw6eYaQE3PKCNs
neV4u208YMbLBn6oCIW7jmdXtOrzIfHczYWhYejbSQHhOc7BScJkr6jJtbUnHZWHvtAMqeU2Kdvy
dh4tRMPaPXBzckKgraOUCHDff9NHwFqaoQbrYIJ38e8otX/h+WD0hLdgnzkUn6YlP3Nq0waH4Zo7
Y3yYzlZ7SwHyIKwH3Pr1GXkwHsklyT33YxfJ6BoQpaAbNUJXSS50V+t9NS9NUTuPR7JCAtc+TIis
cgCJmprbABvUeWCS6xNsT8q4bCtIGcHVw7gICwfze711xsodrmdD4b/kMTbSwks+K3yG64f/Q24k
NTMmxova8Ekhmx4rwkr4mGfqBONlWMFOafDd9TPYOgT5TAzA3rM5ZzTxyAKhyjD2xelXxoFQR2it
nxmG1E1xEXYo4wOq85uvOF/D6+hmZ/juLhREB+ySPUg2eMU+2Wq3EDjJ4d0sWpie1f8pwqUCjwZB
gFIU6gHBleFWg7ifR6st9/TD9U7tGFLbFHEIYfmW8I6i1LUY9n7nnDMrQfTlcVyj3003SZHrYDmY
b2Q2Xtmi6IkQgJSrBRLzgxjgRAIH9/VjgEW5cJW/uzPvezd6jA+d5+1jjIHiy9olWaZQvfidY3SR
5ItvVD/8wXNryXcPqsqW7IgHIYgmgBmgJllolPu6q2W6QL9vnp292DSF9mzZbPiVXC6PqazR4gY+
smhPgmoB+KnUcvlU3HXoralBtCn3pUKhtK5qGkjFS8wgUBnyH+FVPz6ohuzQYm5RErCRmwtrZIRS
sBALA058R5RPKfoM29FVQDrOYCNiRJCUrgT2/0dzui2xSB7cgOKEm9zgBntY29+mkOyumMwTgSyz
r0thhoUW+F50pLqv76PKgLBzcEDAdD9+5t3JeCYf2dsljdFPHm4BAHhO5oKOkPe0rh7G7UCOoUSw
4tHM7h4BL9tiR8W6h9kpyUE4J7BCOb8Z+pegHPVLNnobBrfExI3ytuQDC55lNgiJ1ZL7EuAHM0kG
tK9OA3cCcI/DqSlZSg1q2McTAx9appLKwZqtFTqMgzTp61A4K7wNYs/QZUxCTOfsYJ5905z+l2pA
SuxdhpEQRUOnZSMSmzRSDyGPao8gILp9pLt9yqrNmZYEdTWxL5AEjr2VHiRfqrl4wISQIKHSi1Mk
Krt1ruBrzmX5MLBn8KFPwcmyqImFDQLrItsBX9/LTbgmMV0eu+6j6hDytwkITnANLLZdTPYLL9uz
e+ZdOyw8Szkv9+6Pst5NlJQUoEXNI0UPQWwUpBHdjwTTK4eLqaHcITXLLYgR3a4noFmkmIa/SShb
IWX5ED5Y2ZawR1FZgQQ1l6fv+uHfc2Wh9twKzln82Gqd2PlWk/XcYbvQd3ugPsjJ+ehB6jvFghP+
NqdKyV5kzcPq828y6MjZyw5k7w3g+au/8/LLHO+v5RknVmsJETieR54an8hMw0BLyDt11Db5nDm6
OBwT5v29i4Cf+xu9Uk205lHej3rVYLUPqt0pjx+s2+XmAccI/vvttur5kOF78m15JX4bu9PzQ/SB
acOzfheqDgIGQJ37VqgcKj1s9b5WS1dFkva0SHsQ3VmaJzOZKyF4dBd4i/ZTx5b7u2X3zsN1UNt/
52dClHLnJSAoRc8MTLEqaazD+wK9Q70VMhCwUfsf5VG3/UxrNmAG3ItFEzQf3e3SE9aodKnT74mH
nFQHEOVA8ftopGEp94ugTAR/kxFEdu1xxrlJEWcTKddw+f3AHNCq8tVI9k9vEWmPkRcgqJfcxM3w
3tYjQqRLRvNV9DpCgDy34gcCVC7dZjl6IJdZuZnYxiyMaIw+w5lPTpP996kwy66Q8Kew1qTdJPxh
4yydsgIcYG51v7FtmQcHGa8WDWpCSVcNvmLPn50JciLA/EWq2TsMX2XElhO6Ee2xp5XBr+bWV24D
6m/idAH7r36HAI65MZU25ZIlmuaFXHxsFfxTux6q8GdCjja0dlsZV7j2WoU/FAgNtXRO7LenxDUa
n925rtubCI+Mtp6xemSEonugn5YCEDJIVJxNyjqo48QqqxqEKIaFMCb5Q5uhNU4vu0WNtiEuEIny
cg20CecsIJVKzhO8MrFMsH9yBKw/XO9GAxlBWaXEmV9z5TEcShKOhGEk8dnlL9gpNPvgCIny73Yn
GPKm5BYTA2IZUCPbJ5VU98JSxhozZGyWToVdOXBQrSZNsjkGGIpG5Nh+M2NM5Upk55/pHHlPvZwa
XbsGBW/17dXmJA55p754M0cP/tRrWGOC4HuwhdT0picegYhkL7coVgGlMpaHzC51H2nflpKwogAg
XN7Z5B2O8ZtbPv1QLKjY90dY16AucpOmgjo7wLgjdPZFqzQKBgJ/wJWEYz1DiRWWXb9akYiq/xDf
szwwrAsIqSHTLN/ykNI/nw3tgBXybmWZyFYMWuI4F42pQ3Ooxp72ZTBLgxI/ex5mxrzQF/q4mrGz
77BfiZ2XiLQLnSOo0hRJG9IFNwvc5W01OhEYEB+FX+c1fRpS1NIgJMqZ9JPJqYoqYa5wc4gz5HnV
li0eDcFQEAKbc2KfOZduvVUuUs+yUFT96yN0OOE0uJFjJ1NpVTIG8y0o1fEcq5XTE8eHPd6hLYGR
oFkQD7TG3yMIFAc5YYME7UZvOQCMKiMEnoCFaKpttXHQE+glamL7qh6s8ZEyY26Tau081tBByWo6
HYiPGaQIgqTfzohB4E9UhUGF5UjV57Hf/ACMza0LHWWvhY37DmeSOOid3Pv0AJYnGTWcE8YYRSk3
aDfdrYxbUchZslH8B/uaE+EC/FJUq+mB4MKxCFuUYBuJtqS/vN3NqssxSlpI3M0VwT4EqadK97u+
yOIl9CQGA8AhB+NH6rgJpGWRVC5aaA98w0fyhjnQkkAPsGfR4jWDkW+3UIzrvGCzDWXusgReFASZ
Ib1xo5ZRALXz6Gsn1kt37Cr+GeBdQNooCjAG6TwcI+BDyQ36kOk20DczMT5TzD6pdaSNTs7WoXOD
xMsX/foOLWwf8fZFzCzfNTTL5zAJXhiYnVAZO7/EslYBbFdQZ3SillhKsZBPxzql14fm56cJjTsw
js6fSv9W/AjT9UlDekSNcYj0hp1VU/hlet0VGqxa3WKlTpDJF/BICbz0T3ZeNHu3LkTqRoju4mi9
DVjat4aKL6kv7q71m7dGAsag//KH3l4Fd5ANUR0xOdKbqGfHgNtbzfAjzmM3Vu+jPC3CRGzMaf54
RT+iAShUqI2vTu7AUKxzHskx9dEL5F+BoDyHopQCIgvTYfk3wUAtkoWZogQRz89gqZjj2pLP7Wpo
lmjGImN+mQR59dDJ3ojaO4uWpcxSL8OTEL0kF45UI/By74t8LCWhvlSSRLm39jSGuqjkTMLH5Neb
nIUCpBJG0iR4ku0a4vNtH0odQJPR+YjEAR4fXPsRqBbuUU4R4EgEtVtdFqK2qn23jQFjBxxePNG2
LUlZ2XUKtc2hbthaMI1SwHSHVb7rFG0ZJkmFjxuCSKR+aq844czRl6FnXBTL/UFaga8TxJNE/KrL
Z7q52d/++9osYwPrkjez2r6iOQVA0wppELURQoywxhqjwsEtnZxGhMAw7TawEtDMbYts2JbN+4xe
53d92bZ/9h1Azg2vYmC9Ot1d/t5jwJZFR28tBD9I4SW/apskVFayoQVxNr1A89prqkL6f7Hh32SX
paXrtiBnVAeks0LWmDWDZjXsb3P2O+6Cxc7EGffavLoAyZVTviDJVRDz3z88NKmfBP9USM4cJHP/
TKzAkwTTB7nND3cZWamiCKn/Q98HEhW2kY28B4lQebSKTLPSmtxMkqCtXSKIBWKMRO7I1umaycon
KjfdHhJ5EXBl5VbGH/FJa9J29NyVJy0MFQhJ75r6m+IWYesXnyvgAl33Xdx+yCO/o00ysBbospSw
Yu9owL2He8ZZvz0R9gqtAQP0dpA54u4Gp2c3gVp2bg344/qQv3xCn460oxj66pmeucitvAKs3xcH
IXjRtDunJz4opZiwHueX1MRusnpf62iIeGQt+RNinqP9G3kegaMrOiV3x33+YguB0eAk3JvBwbw9
0RbDGZBQ0wpi3h3MFYCi5Gkobfx8j/xHdt0ZdLIMw22jfAeZ59W4JtKPGDL8MFmYplwjupXD8PNj
hOdDibla+zoDbDboORqNA+7aWJldp7HCQuLdNm/zxrLAEB2NYxEi+sbRot9iUjbIxPMihYl+nUY+
9eDG4IhADaLQDRgEE2oDfQf12xFguRCso1q4tX+VpdKYF5KGFOTz4MBMqaJWu4TzRAgsnl28+jrC
Z3haVR8vDHpoE4yhmjgXl0L699c0dMrvexcr8XvVYq5+Kpqafhc9LDETY/hRyn/jRJI8zXqfg2Ju
mrbgUod1SevaLX0+QQOirjj3OvlWmRoawtzlJvuIY8aGpEUIllprGKdoTJpQnCMOfre/axkE4HK+
weDFOSEmhSvLr8hfwdHs++cWZhRJNZquXkcUQ07a1jnChuUX8Ne/2DTymjv4AQvNyuiDYZDCRDOF
Her9iGL6A3QX0W2oB0jynqLQ2K4bI3HX+CVJ0CiKHkcrqveiDG27WWlyHb5sWW/3zfEXJqior2VW
5JS7XS/3AwKA5CloWJPxKDq6U3IBQ9QeBaPQGvi3HWNHKrKga9qXOWXW8XpnjdEfwMpuLxXCDalH
EqQbEswrp2KCUuZhpbsXZqs0r1RKqpXBiJVXwONiA31LPjocEqVuNs3szO2MyQPhEyhBU9PpP6y4
HRsg6km2WzikRp6wWHYFW51OuDn2ZCBwKhZKM8sDt+ApYYMNpNTe3q/UtHckoWEuBRAW+gupddpN
Ui6EfgCwmbAvMBw2KocYOguDR6H70vKN8HZN2r01mbtqqHr13TzdoeN5duoaMEmjPPJl9tO6HCY+
qMMcreuZF50Gzkp0Q94zjKZ3ZSp0wdJDGQzaJY77fUwQtXmCeVAz32eoyY+an2geetqpLoS3+r3O
9uK/GLzwogeq1FDIovEHBfvK7siVkPv6JURPJ4VgoaOPjRguZV1CHFiW+Nix+sBQZiIBtLxfq+Qf
IfZQYtv3znAc/y3oBHSrAt6VbPYqvNO7vjQWNWjNlC40UOR2bwcU6hXRbE4aQ6A+MqEi2Jru1Fyj
sXzTt7wEHMADSiL5v68a9oqZNF8vAcptmYYApDEctrxAzFvdfI9xwbrsKrwoQojcIWCVD6b5LLfd
6qTmGnT1rUVyfQgdVW+n40u7gX4Fwzpk51meONlPk5K7MbPpKpB/cciy+5QRvMx5M/jCxrPnIjOO
4OYytnrhZOVi12O8V8t9ybJY0Hoy7Iq9iYrUDEjSGjk56Cvdf1G4kjoVNTsTqKnETV9uKnhqOIvq
Tsp/cMmmvMO68CfknmqpLeyWbZUBLvFc5G9St/y+9g0Eh8w4A5GrS6gEdqEq1KVaH1iJNV1GQyUw
PseX6lUr3N9LHu5T0brirg3FFA3DF4kmraamPbXQVGZ26sGQcjfUqcx3PJhfXe0ygNUXsWrQ0ZTC
iDnTZqnnjgWXHmDlxymezOOoWSisK3oGQKg0fDTUss+SM9F0yB9bNB+WmsCgshXDO9tNR5tRtGJd
0Oc7NZRholZl5GA1PUz3HL1/MjTVCDZMQizcsAAf4rnfpAkmsSibeNcfzbzcboXot9ZnimDjHEAG
jJQ/bY+spJyLXc4ZqIslS67Rjyl8HETdQ1B0jfi8K7Da+oVnyg4yUD0lg5S7lkv0R+DVji8eC9lT
YGWaRfNUpbTp3wibFM1YSjZEuMPqHCh8sysOJH5cCpT8ctc1UHDR0ree0CPvO675DfCX38oH3Cum
z4c4E35EkGpW7dtnrKhgW96mwJexmcxVZ1W/xVtVKMUiSmfm1vX/LdRJ6cR2jXq6Ww8+2JECXz0L
xgpHxo3Lfv/l60pgCqE1E7AIgVRzQJXRiCtKCt7vUeyD2+qyRQKwGsPTC8taN/iyz5UqZ4iqN2C5
r7GCAQ2DZyHdeRDeStK+GBn3kVUzRBzUpmID7iue2YfwAMaXfqbbra0Uy2u3Fkg4bRJmLDRm9uh6
G+DFdkcYVnNynVzM/uhVJtInoVWpO/Ds7vH1cIOvZEb6fVdCWHyIboQnpTLjOLHJGznoKNlrsagr
IxMlA4SbkJ8AuwpIFzzp+TeAHfdzOybBlynwFx0wxfUh4mJqABSKt7m9H6JfMeIbzied2PJ2lq1y
9l6HRZ8gSwxnIzUmNXhzd7duMKUa1ds1xO2mt9hkzpCsWju9rNdmytXEoDIVhzA03ilHNoPF9FBt
SIRCU7yxlv2Njjrx6l9mVS+o9zZ8ErLnisiwwX8lGifiP6xagjPTNV1LxKIp2ry9Y3XSOuoi8rmD
VCVX4xsutC4qohhzaStnr43WrN2VObwBowzBwo4MWXTnalEIdI14nsd+2+c8/uAmEpZ9jp2S4Dwi
wPYrKG+0ZTv/ZMEhAcAYnw2+ut9UoKTxLxCkoK3AkHsdlE5HECm06R284hFOowXP8gBfaifPhdOs
ai27JsodxFGuAmRRFGHcZwePVcqzsCe/mhHwP0b2YhGOU7x4x5rMa8oZiPo8KKh8rdiIIagEjxDm
51qtRBv8NTQ0jIs4rGe3hCs6R5hWEnDrOyTGkd7P+ZJuleRMG128wHzUzPJ8eb5AMhZxa4CyIsvF
0eYfwPhPha1VBB1WoRgJUp6P8D/g3QqpWf6sp3XIeA1RKCj3FDKGHAarkx6uNdiihzQioFUN6oxR
sLBzGX5ScnzL/y7LvNbb8slp2PCxBHK2txHjVj8VjdZR+nuVTRO3y102GPfFeZOEpugMEzTHunlr
5b8YlswVH2GP0cJc+GxE5NL/x4qYUilABC+ChlJ5tRj3Swsxdo4QwRfRVrqIlf6SrlrKbT18y1CX
5XXQP0uZp/V5e+3evYHOkc4E/RX6TQ7Pb3Z8KzC7CYHSj/a7pW519XaZY83Prmxor9IUnxtNdX/C
0k1CmZ5O7HRBygxEE+Ygyc1LzPh4ZYwZfK7AC/UdNY7PvTr64Hf2vNgSpa6/ZtdTxVqtsNw5g85B
SGEQRv1qBJsY9MTKh6rCpRDWUtRMJUoE3K94oUJ8euFMWHAPeGi844SFSAKy0fJYmeqsRhNEtu5w
3e50eQ9ESEjxnxRKV9C5AKVThiWqnN0XPsEby7A8qS64OIyvoMZ+5zTfU6FMy9D/FMolCp5LnK//
EbJKQ45oBoKKSwHaVKXGGl27hJQMSEo5C65uMZVOUcQIxsKOkGtblDVZeFdGXY7jT9+sUAlMnYBa
BNEz1P1YxmkUZ//TxYooTPvvbBkCxzoGVwbe1+u/n/LOPOPWuRjci7Jysxfe7stC3Lk3f7LoqCDX
p0lHhDMlEYrDUp2k7FTqinLvX+UlS6gWZuiOIkZp1CfWhOgQ5Wi29dGfpA2KzHHW88k0ci8onq1P
TzDweAnzPFRdEPCy+eqokceznlPk1AlfkpdzSKRLmrQmUGhYtQvlQ900gX5SDxuTIJO5+xQE38J5
VN9qHrRnqEnW5uwSMNX/bRq0z4Dp9rCtVcdzx9RzpXop1r24Xl84yn0ncmFu/6J0e2MN+yfmWLJo
33TEp/v7AykUNh1989wIWohZTF4+/SF0Yez6VCXovC7siF2vXpKT8jmWsCGzVKgxtxBMtyRT/Suq
UWO5rXlakYarqYgZ8H/68Ed8sKBQh0v+5FQgUOMy23QibyfT2rGpdXWlc52AdR/tpVelmFL29yat
qA/lZuH3jJFUoULKIfhZ0bIB/jgXCFUDPKJK2YdflM32fR5fOIFfOdaZWvb2ziI/oHMSN3wngBHU
zSOIK9j98NJg1T1Fn9ewtd0E9Oy0W4wFNgtSakKfZyX1njKlgDJBT4tF4zFchTYSOeWcaCCmbbzi
2PmW1AuCA7xGE/VGEx8YhyVSZRY3ztPCieiQIKNXzaFwYwNqOow6UUw9RfOaKTKINdtOF/Y6GLIx
C79TZS8L7tptfou/Yut03lLVNrCdgPbojieWfqCVDh9l78rAJ8if7vO83z0TwIa8jP6Sl7/hG/u/
uI/PUx25cFlcBXAPQftoC58op0/GOATMsyr4JvY1LeIFCeTnHxdMbgAw+/i/sJ1p3H1/tJt5Woh7
A/owLPsks/kKmQhBw137Wpv98qFzLD/8o6bdBw8kkQWFBzN9APBnaa/7WluU2jabJNHfJiBDSGX6
CEW0vSc/y1El3je16xbTA7DwDENjdglsOkPB41Wgg/Xr85deahQrcTMPS3NTWBnr8JH5fRYR8uas
M4TXMujHHjtHbKTzJvTMjxU64lg3UJJco2fgOR8W/Ntrvqx/vSx3uuB3VqKT3y/1ItXQvUH/eBwz
cIy8cJCPw2hspdW/KUNmFNI57vkYcAhmDwhQEJg0OeNR/FZ/PeltcMN8Z9DQiWS/IMF+d1cqyis6
CzVxhuPIkfcUsZK+j7vNaid+ZmkMtKk69Fjx4iZrd9fMbvLDZjsT9TwFcw7p9itlRg2oBd4BOYit
stOH8l32m6Jh4yNToPdBGbZOZZkbYtesoReO8gHPb1e+MkyE5Ulr9Ofp7gMtq7uKxfhltXlZxVTl
jo6U1fw3WTcAgmz/OXPcbL7O4PPqH2zxqPpFbfHHDc29GhpXfHHYnGWSceA0lJTVtTG4J1h1aPOc
UmIa12yA2PBS4WJG2EKnN6p+tudgMBxd6ewjkdk5OMXXpKToG92ArgAFat4loeX35xGPaSLjZJaj
MjLvznptSs1vF0+t9vvqNZIo20d9UCZpcDodIcd/4BQKpwoZ0nc7LboDk1R4SDV9ZxibaRbZ+dvV
a1OxtzRMDIkhdNv+MJqudWSDxAV+ufNl1YVJXrTDGg03Umhze7SeN/A1LpbaIP0zQn3s6/uajknH
BpnIZujLWpmNxOXbVG+mUDXlSEMiPUbG83ATvXh3hzvjWFu7ZVTOB4DOpU2m/XUiB5jDXJf+a0uJ
dM4ErGCLxJ0OH6OPCMzBwhrLPsrQ58Mx7tjbs2nCnDQP6TknQ/BU0FpvpzOfG42BvCJ3vJX6AsW6
I/2Hx5+39l6uaHMPY2ArjkN+08RwHlb613PLqBkHamimT+6oyfDqDtIXggAeE1MRf79cBCd0FnTB
dPblrmXhJApwj7TyvStJbYyULw23e/Vh/Rxh6dR/sr20nf2C/R/XMGHdqKVBJ8fLHq+Qkfotm7B+
9GX5smF3TrFpSH5VA98ok7aart78WTt2s5+Vf9RJBMWNfkf/TCB8gXFc53bDz4GEgKWFmFO46x4e
KEY722/a0rYRQsiG5mxsgDyrLQWR3dv9uF0Gd9VuO2wmmAl9c0U9GIHob6RG+sdecF7QNz/BNDq5
yY17FNniAKkYBACALGQEPLu1IghmZC4BkS0motpOgudhrIharl8x9fUkpGOJ61zlJ4rubW7LHnuW
8TR7UYpEZiO6l6wr8zMGjHN+/+mH2JV5vfn55mslvrPduOJHSJNuWKH6v6lJ6hGf7yKOH/yma2ju
uskdVWlLTM1jA3693EHr5MRzh4hMeljJSg+V8yV5CtZIYQCYnFi9OaO+fMgKqNrbRgoO9Sq2u1mp
rVDl/eJK5wSpJhjdeOHXxnrSDNyVzKGYcVI+c05/Fs+43a+7nb6666HIxl+Y38xh5JbEfygHQ9/M
VTUkOT6ScXty/naFoaZ6qlxTPbkeEdZTvdE8lR/6T/iWKQEq1ofsZijVKD+7mA6HMBmfVkDaaECt
ijKfYCUmvDmfF1zEe1AAVglVm4uifhum6gS+E71Mp0zlMceXnn7TikOKvmcrdLrbnxYt7wNRddF1
gqtiSFC0hQw60aPoLGJtIBIyaUWAUNs9YVHb+Dbu315U0KNjGIcexplMbnOMKYqomQ1FgQLHFDEL
SWTWrPKkZe1SArnnyBZM19I467hdQh2nrHKloYAmq084o26qoYdTz+7rXNI+FqReuwTV66/Z+Mq5
4bmevoer8hYJYCoGDV8neUdOITd2zKL9E2JrX1NPHBAaaiMwYcRQ0gDRY7bbS97T2m1SMpG/mF//
5xmgZxTQhYIAibALdAOb41GfWIzYRW+fY/mdrQAQxXr9RjVxQbHWdyjGxNnbp1Z45T2WHK1O3RlM
i/3JQ+eeMSTK8FyVwLH88HmyDSiUt2tDzeW4OXIyv2u+vjGNHbfw2OmriqKMUxi81zdNxG5di2dZ
d4di0+ZFNsgrqdVqHas2aa9UPh4uDV/OSbsusG9NoOyy3zjNZyzBrwPshu19EaISu9mNJ4tVIJgg
xuC+2ULfC/gmrfKYOxSGKH5KuB2SqanvrdlYFwMr7vzDlZJD4vbxUIQJRbRpgL0+mMnrQw0Ji78b
Hfu7/T/+AJdzNQtZo3iVcNsE6ftZFm+rOEkSGlgfey2P/csHJPg0zju7ghpvOZUL1ogPG6tqZpo2
b3vn4vmmCqORSjXsyrez5yGCkVcunCE7WN00PiWsBZooMYG9MM2LgKZin4TlWDcdDBOyzdwnNRE0
wWRee/HvdPNG0CjGDvWsUy2C/RYDYrp1wH18SbieX/V8WJiAgioFSkRfLMsK602cVRB1gq62T5i5
vRZDLDFh5Po3RiTUcYXs6St/UHJ/YR4UcG+M75Myy4PfhgjIl7iy3yCDmfl+tNHlIvahWW3w934n
VqOtu4ZJIkXCRnxyG485Brns00jGuLBBBCXbajEWhM2+V9Za5jl09u+uqCZliqH9f55L94Thsk7M
fJgk0hoTs1HHrsCURgTAnGfGr59T/nBgtO98dByZl4iyzCsCE4DuvhXlDPyBoCnBtNW7gl65jaFc
N3mHmTNsHq70goJuMK+HXP+qzzr0MIPUXOyQM+iVw/zpQT5wMgxhAGoYwgZWk8XokdQEeMqNRMOg
NyHY+eRWHXviuv7Erri+sfJCviTPQA6wPMuMU/pYbv9rvgpvG/0XNiwrwP7qacV/hx0l5IGD7qNo
OhuIVDguQWrbQDGCOlL+OWXy/efckdCg6EX2LDNN6jrIEmA4FxZ3vXacBup6xr5XnJfYuQFk/+E+
ZcVJEJkun4ci+j+nAzYQit52EbXLxHbkHVCxVJg8jhCA5QVDMVW+GniCK/YSF/N4LoQmngAr3OB/
D0N+Nxx1NUIbmHhC57/FXKw4HJA9JlTbRT5usDXs7A0shPZyVDQGZFCC2xU8RmlyzH71B6JB6c5W
2wxvBsMuNTwzbgvnzs1Sw3uVTQVV7u0bvM8ByVPbA2xFJp0QhTPe/06GFvDifcwLc1HV1O9vJwa2
4lw6tl+QXRrIbsSs6WUOY/Pme6/ZIvLLqwwG7w8iZUR0mG+QpG5ntQ6lGTf52gHfUe6Ih4PXc4aB
2V5tRNACAtqQeLujsteSBVjw2cgKURM9HmHmbXnPpR2eWFo1F69rcdJ5rFATRBHq1FoB+ZI/n32s
AlYG/chZnFRIgpOu9jPMjQ1m8hrujx1AZI969Pq3u41F5cdKI4qqnW+OVEln4WM/il0AOvkid+U+
9dI7h+wOCuSr5D57TJD2hGTIvuYNLfO1HnBW2doM+Bjp4rC9VGPEV0ccUP+6g3t4XMK8YOwkOw7o
0RZOyXNncuI2nCbkhbRPBcaX/yl4uk+SZQpdm8HHQzZ0OU/RD+wH0Gygf+0e+3+8Ye33kMQRo+oL
U1b2bWv6stFoTdik92TG+OKVQHe4IN6+blByIsP0yTndUe7RySSku39oojtufTLsX03aUMfkOmBc
pV0A2moYk5FlBqNrD93kWBdU4+rei/0h/0lv+wNbYQPP6zcILPQfk/cvT1wG1G20pMxsH3st/MxQ
KsNZ8TaNK19kE/DAsf4iQg6bF3mdGeowc1D9VWfy47iRe6+7h+ZLNWJJWyql4I6kr55IbC5nJjzK
itve99rqxEbjXTXUuwv7RFBpSKi33kT05GPRRYGTxto7Jgovc/kuoqauAebtvtfpoU6nGcXV7eAB
pWyXE/KsEFtiwiRbVMdnScWHl39eICH/YMSZqQq7yBJTWq9Nc9pzR0N/KbML82g6ZZh33qtV/nNw
qTbdWOU9XrfK2ax3/05i/dkTFfydpM8UBL5wuOSlykXV0cAdnXpgiOB5wjjJOY+chALK7LOSjJUx
HCN8nYLMIQlPzhLhsoIWItqKWBGrggOKRJHmXmm/yIU/NbYnpEOyuOpj4nSGxblLfg8ylmAO/4hK
L+GYdh/z3UI/YWGNdGVps7ifFw67PukpA1xc8SN2KJjR8hbOO2aRLhhZohjkYmTIDspeaf+QvIvv
77TWNMltYIJrEjlBNKWSxF9d+4+zXWMDWa7MPgIUoxIoIQcojSBaAv41I/7cVDkM+O6zo4y2bBeR
vXoOrEddgdITMNyV55Br9YMUuOui03QilbB8l44qOvsAnAnByBVDbF/YiskXM9HvQe+cCpf2z8O0
dizvy8Y3OM1SPkBscS4USAA3pRR66iSGe0BXF9C1qKdOt6YhOi3pL8BWXRytTBYuFlNNRxDDq08c
Bnxfvbc3tQqbpHkIMfnG7H1+EWM2SNn73l5/3FvtwLAsy+034tG73Avdn/8tAiF0t3+s2JzHHXbf
vnlNa7GuhNq8aOu13RbCBhpF9/+3WPuskzPf7Kfw7Y4NeDqCKUWg6GC3bY2LrD/lpUCQkeJHlJDF
qtdlTJq/qbaCrz45BsCllufmSX+fGB8+xlG/d3rZKAruO7zmJOZMZYY+D/Y7SfpsGGh9VfLctWuL
JyrmZHV2OF/Enrm5yYULgx4a0nIY6mEKjbi8g5EUt0CMa37PhQ4taOpTRRqa4/To8cz1jOABm46H
sXHKutb8m/ldwB9AcLtdiA62BtQIJek6xWn+XYrBJRHe4N0xCmypQ/cFukWArmCo8toOjsklDmY8
H1P18vFZFcFr/ljP77diYLjcy015sdxEbITZBZnH0EbQNUphV2wzNa8ft+LgFcVME6SM8pYKC+pr
L8ePlynfjtv1sj1azdzPWJPBUojXVsw331tXlsV9JPoOUgEwxAh9f6r2dQqbNhI58qzujn9lFfxu
ZA8Vh+fblf/c/PDgXgtAzarIhoCz+MwfbGSscvy8hrT5wfhn+ii+E8fDG6X1uroF7jRYTrhgGpIp
qTAe8MntRawCsqpGrPt2KEGp+sWWr7FsQp/WghRLLAYFpenOBGnEsWw1+8N6ryLGHioqvx4LxGas
kS7XrMAHFaTu+92E39+QEQdzyh7maw//KMG5Ak2uWHBrBZUx0dn2VUXp4nslFC8sPCdyXokybaMC
y44Iwvz5Q6gBeRJHFIaQ1m9IeFld7RlVWWKFX+4XFy71Qg8ez0BZnIema+doF8rNFuQsEafQWZyR
8dVEy6492LdB0gvRR7f6BaI1xk7P790O+lQGCdYDM5tmvwrHzKTjwJp7tXTTgM3o9zvNRpG1nf59
rujK6nl11L3TNFA7y2d5Tzh+pPN19trpdTcIlabZY/181NHdK8ZLTQAzLW7kiZPVBEDESzfKB5H0
sQ7+eevEOWq/MLoLZaL6Y27n4h82AaX8AxdXxaOb31BosE2BEM5NhwUf/Oh3/hiqbeWPOKtG8zjZ
cyyWD2KoKIjDj0JFy0wqDRWNhFbaZ8usUEDg0SjJ/fIZ3eUzVe1sYKjRCa+7F6+xHnF47pWewc0U
sv9q5XaY9e+xmb9OOjC5MVPo6ijMQlPQ/6vCvo8A9VfkMJklxz8sKPZnIb11r7MAeZkn8nRXgvAs
q1FQthPkrng9ZOgya9a1HVwMJdb4uKlMJnawPkdvb6k/QsolaYsWqzc8olez2wgYOjQgYOYUf7Uh
o3wGrAQLGVeFhwAleR3ahfJnuLGpk+vS3vcw+k8CbcN82IaBfkVm/sQkXgeO3H+icEWEju7GzBDq
LruUVRcXUm11FVne93NyTH3mXoFe2JR4RE5lcAmMumP7zHPoUOuFNb5uWCHgMim7hp9S/wjfMj98
Em5j1WbaLkRkMF1myva0TArt19e3xqvsCAbzMCMgM7qFEVcoy6yTtLIwj1Q8YLVN4mEC7SjTWClB
hdMY3rO9Jc+5f3WtAt1n/Dm3KakcoGWsYMetjzbokO+9U9XdzkSCPBKU9Cge6q0S4GgyHmV6UIKX
zaJW94B2jJ25w5IN0VBy27oOWyR5P0vHFsIyRx0lp6z7bpgnsGizq0sYam/bRttx6/a2rYbSYoLP
ApWSohIbhQHFzNiWFyLhfCckeO0EMKumLfhOtdBM/WW1Txjk5XSmSMTBP/cj6jMKPeu3sfwR4wyu
5Ahpma+Lc8TpQlEI0W4yVNEJj/xeagkqCv9w6aGc/kBbAE9HtWInnb8pr0xetQ1rQ2q32M6o/WyT
B8VDvU42HNbnhZP6ew9H1GZZCbI6JobQo/lBbfif68OJaLDTJg5bDuQCoYWpyyy1ilV7uPZVSKH7
HswCbgHIaPB/Ivd3mRO2IN1QpF2vdloqZPBT81xsnPa/UHjkC296RJETZIQtn8l7HrIxurlMW1Bg
5CwVZr+rDEBMYm9SQKco0nFknqJvK1v7KuvJcNGb/nagNGlJCBA87ue2oab+Fs0/DWT+Qtu84UO/
kJOvj31APr9Qzukz5mQOVo+G+WkZ6mAkA1YGkH+gcVY5T+vwt+oulXSmO0/xJiWiwbwz6asOZwFQ
hFFaVeqXQeluk2+F1j/9mG5WOCv2Qdn7/LR7EmYrlDsIfbCitJ+cVogFMhomY4gN0n0QC2Fx1yUQ
oQQxBRUH57FMg/l8v2MQrEjr9bemN8b2fdviheTDdkor+33Y3OF8fehShWfpXhDgYD7Tt61XDMLY
VaRsG5Iie1k410zxiwuEHkn+pjsgKXUC9IOCzi7gD06mrrD5O++P7pskmIIMPXvvjeZG3lHkp/8b
mC3/RT5/Hhu3Rfqe7cm6qFFBLek8DfXOT3rr4x14cy6fXxeqzMjqwICPWNb3Jr8tewdROZHf5fg6
R1Lhis/CKjPCLj4IYnk6R7G27EylFyvt6N3RI4cm6ktXjz9Wu/e+KipKtdZqNsBPIoQU2ZEgiY2m
qRAkeCMc5cQBNEi2srGuScajEvvOYMvmfJm+kb7wZBL5yPz6uLnQCmcSDjuD8aeGiAHAlDkrYBKe
IfdqClb9pzRwI7utKvLQNZoHEtVqP/E8uSDCHpQLRLJhmrJAtJtcrapJJfugFmsCyU87iqm9ftR3
PTCbH8FVmcVU+7LTOfkUC5NlFNoWOCd/MP/2FofGq6kQ1i74XC4z+RBIS0wP9yZcAupANWxBmoks
sp4e3s0hLUcZOlkXFH2LycAVUHYmG19K2BF2GhiRBQb1J7/2VW05jqHNxk6MKVwFqF7xhE0krNaB
lIjWtY5juGyoY0veVH4vYidcostMxDS7vwB9Qnthn6ZdzBkTyH1uf/l6eEzE/yIh60bxnP41xzKL
Qftki8IXkrCQzyreEesYH6IgJ/rOI/4cNflxWFUQW4vY3gbwhrsd/6pK+tpY/+i4wSQGL5DadHs5
D821DVRdC3Q5QK5rjbRhdqoxBZfg2l4CpGmFfVUvHXouCeAzW1dAKo+DMKu3ZWle7M9XlBw6tcLD
jUS/MwQ6llyWQEhzvLKaCRHk0NPijWmB2bPLFqgDLZyflj6IqkUszoUxXfagrxwcOcFpkZm/X9/R
4dLG/5nzsdL1GxoMHeoZs2tPlG55tsOqhD3BMk/HvzgziiAZxe9pAtUAV/OVzGNSlrf8Yf2EXGEe
uFt7p3YzWDhsYsFh2iWo1PidgKpO/hcufIF5nwCTE81jYL0L5eAqZ/LP0MQ9//9nLaQ4sBmIoKBe
bsZtDxJDfph+it6tpnF32To6LtNF7PPRl935bOtWJKjqe8m3O+pvW3PQVJjWfyi1dULE46Hg6yzS
UpLHstFENbhpxEUyhxUPiTCdgi+MvIIosUcYB2cERakLoW+kkxd6DB5Y7m7fAdl1qJglxJA1dWWV
koSK/RNm660lCEE765vMmCM58a0pqJ3uZIEVi26ff8RGaFdbK7w7Ogd6ysP4Ia0QG2c6N20KjfYe
msBQxiZ7h87o3XK4H2BWbrrJgDKuWF09/Kq75e2ABQfjxwb/+thsdF7L62/iFh48Qmql4Ns9eXlH
fRZnu1xYMm2mKCrVlY6TY0iiXC4L1U0agZ5MitV7A88+OILGxM0DrrPZZ96P9svUwHFG5jtVGt3b
F0cUHjZJRFK3LBSLUmKiOU9GND3kG5ZP3iah+GKZQnk8ThzQ6d3iinapLpHJBxmzA7QpDbC8MOkG
KegoHClQAJ8CCWNp9rzWB0QKlJClp4OuonqcrQtps7ByKZd7vaP1zADceLiRzkY6B+9ciag562Av
CGWjmyXaUlwfRifhS3sV+mGLqe10b4co4qt1XcQR107H7j7wM1luwpIchSJib40KPTKzXDCSnFlp
CR94f9+pQbXs1i6Q10nnnh0ndFy65qjOYH19kBb0Xc0rBSIE4VMxpcbOa7oQehS+mUN+ho+j+u4I
H22bDTCBWMiGZ9pWgbAf8aPhXCV7KknP27ukSnyQnkxpSNI6mkKh5sMSMjC54IDUVhZXT1hHPv//
toWFqD5fWz6bSnauNLkDucyE2t5aQQm05+mx6tBbw3X7uOCWzu3zuPYOIg6HTDdnknRCZv6aKxXL
GUmAO+TIA+iswqIoH2wrnt2FMGpQm85MtciYItDpfy+aFLwQFZ4gWLg8ywUnG+/tBrN7KHtghkMf
kKS9ZKg1YNvXdOAkb+bcI1y9ykh2uPh9pNLxFC45m9dF7uedf7v/YXoWmQjb3n6fEL1dIE9ZAJmW
8mfVcQasPsPEgJWkuvFotHvjMkvqSMYiY5GC6LGORWQsw/JMSPa/BCASLwxUq4xBuQFXcmbRES2Q
24owaCmmsW+Fqv7QfwJY3sdlUBCqy7/jReU0dLn7twq0/q727AOc6g9fq3TI7X+2B1BfIDUANk85
YtHsKBFxVCBsSzDC0KX+jvbwUO7ol67vkg/+v1k+RHGrAxwc4zZ4h9AWDM2/M/9NAUjfQ7Ehzut6
wwYDzXgP/kWyY5VSxGmGztfLQlWGqfDxoaHsguElaxzIB7HK3AhWSDFsLwUX9fJsPaKHlzprIeDp
bhFT3lGwPBp6mxMoAmXKr0rHNe5dMRRJf4HkIIhQgOAAhaei403ltC8ylHRcpcv/GBCFao0wO4V8
bbpTG7xTmvbb2rBrz99fZX8hwSTeWqXpOYA/W2KPsbEhgSeeVgagqPytQ0NNfVVo8zJc/w4lCQiq
NU90hKMTzQ+YGUnLeZbCn3plIn5w0g6ztAH7Xfon4MJgX4mvCktL5Biji938x050KoPNkXOiP/gl
Sj61G5HWkrtpiomfaKEIOLz/QjTySXSeK025PyXAZqVSfPBtrXIrySkGNPCuUjNxdx5960WcSG2n
0gNO5QrAEAZA/6ywTIjCXfD/7+bXoCOCfsyzPkvlTh8RZIoHX/UG6e7hgOBxNTUArz7eyypLKGrr
iaHwGNAkbBGFT4Ch6AHmLPboUuqwv7HfN8xDw5fVEU6wAXEXIGQZ7XYMeGsH7QeHXaFhUaQbZolm
U2kdf9sKlprJq8u/2NnRMqKD1FouRr7W2qeXwrczEboJrX/Fqa4FmM/rdGEqALW9DoNQe2u71TEb
W8b15RF1HDbGvynZLEBkSxP2vFk9AGHYFF8U92aqZlG1GfJ/OvRs/5/H44SgGdeplQYJaF/Lllfk
SEhmSMAYcJDnu1I8q1hwbSqy4TWCp/8lk3QgFks5ET4JxiU6LfRhh+KRvoDeysXLtY9ZAOkqx3XC
duoeMJ4+tvFKbAsfOUTmxAcyjDYLbXwWsrrOZ4CjoOC3p5QEModyqAvM31Qfu/DZ2iO6yRj20QwY
1t+WCI9Bxc399t61Tl9XPvum5yjJuLBcGJXrUyjbaybumGQHLZ1o2wDd94XlOSHgjwAbfO4gorAS
6rSo0jNLNV2Z83w8Fagg7azsCdj8NMYtaPuQ8Phb8puKUm45MNawdw4dWoL2c9CnjpWWZyDFtNre
BVK8Wj1rjZIGrbX2Q15m8bJHh4c4w5NBCt88TQLIt8VuWm5YAVI81Treqx+6320T1dqx1tOyy2sw
rm7hcqdoKtI3H0GD2MS+P5sfQpz+XDsspNL6VCddQiIl7jyWkKRNqSv4UuhZ3fT48PUVVWkMbose
N86T0FQljOS+kLpBxK8f6wmlsjXmaRQXjom9AbZVi7coO8+jOwQldUzfaZkqgwTkpihRmIb9Zilk
pyIN1S8N5pme2FEXtxXTUQyOnBIKp+VtqR8BJYLuEfQXb0XyFlyz4Jpe+94/85IuXU0vBs+yP1p8
KMdzN1RZMe8Ksyob3dkNj/3HgNyenWeH827fctJk2OrB5esEET9SLBh/uosPoo+7IrEnXiqDBpeN
5OjrEu1PlsBcS3NJoIrVz12S8nnzcmz8UCjrxEJqfo5fW9m8pbPbThzHVszzypgMkaI+KX+d5bHz
HJXKE3poU69f8H1rlDqza6OPe1JFPf6u12lXDcZNdL+GIkSmDpLKZkZyM2mMcfV9FqwVuNX7QnNX
2hrshAGdGikU1bR/O1z9kdAi8KWOhtsR5lZbOrS3Y6evJ+l1agITGX+uyr5ZhabSVr7s1xfLnX7S
jHGZmQOB2gCtVrQ79S/7VDOQosmcJM9zZNNN9dK7u21K/oCgVMv+LlJexQ5NpjrHEI1aRkVqDxuR
Q9A+69JGU/4rNxVNlyOZ5hdpjjiumpb2+9cEqpn3oQSIHKEGfVTUN2h79B3OeEb5pIn60B5l8i9f
aa/YVRsQI4i7z1QhjuzforXyuAYyCcbyLZ5j7E9MpwZwEmcuX1OmWA+srBsUky2ZsLCBKzOcHyUS
Wju9aZS8xX+yJ70WQ/gnV9GRlSbvHHEoVuv4aKBAAXa0lYHOlP1kOg5L0lb/9dXXQcqzr1jROTw9
vRJWApVULoTuRTs29cEq5qtsHT6uo3xwxPdRsEfYdYI9EX3KAI4MmW+0JeZdKfYqPizbHeXvjtVQ
zZV4yYewYrJUvZ9WuvWBQ/JlaMpF4zalftAvSgCeDlZQIVGkfZvpGZ/2uvsPw7eFekcziQRg/TH9
PR/pU1j3F7czq4QRr4Hgdu+IxtyZ/NiSdNF1yTpC7EKCbhKOUt0R+znbFFJs9Se/qDr9KjQdEU2S
E6MCt9GCF0fq4b0HkKBlZr4v3wIB07XK75L30gpTBdsv1Lz3JTonWsM2ueockxTHYE6OYvTWZfRU
D0lKA56BHeuE2gxpKDLJNSncKArycXiPAjWa2pHYwLf1OxdzrzSm3GI1xRh1JLUOYzAeH1WpfUnF
s+mY7CThu1x759d5DONpUyOvJ2K8qMBqCuqzQiW/hG2h6fwUUWhaZGcJa3viJ6dNozm2dYiv2gjv
eIL750HucmlVDhn6WM6Y2TW9meKe+h0iOUAXi3WxGVBFb9AhX63nerfV3O+DvL2xUiqHxYUyS4er
GS73ucr3nCQ6TWSWsnsrYhmdt+6WJcJc5fnUtvvHCzELfu0iGrO3XpSSBk9s5F4Rdr5VykZ86Hvt
SWHRU4HIYbZ/h2p6rYoGFDpQ7Hc/3Q8/naICmaEMcGkm+2n151aK1BCPjuMpeyUCkc4ofu9gv0PB
piLN3XbucYNpf0CCaxEXVYyPJ+n+2kOsWmmpug0mVzq7ZsKFUJRQ5Y+tjIBazsDmwksAq4Ks0d+x
jLpREhlle9MCW+agbdUjB+LJvNy7OvpYxKjpwZCChYEJRhVYNO1H9i6hd0peDl+/ur/Ex32igl8u
GEJDioeM81gpcBjjsmPTVIuhxahckGNMSi2wDwYE37fdJyH8F8h1hryy0HJeg+c1fYE2Sb2k3BxK
SBb04Yj6BbSgJBBLrBt0iFiClGlNoIj1DACgEn7Hd3nkRUGkeWhN8z2ouemPpQUyccDOzoylX/IL
lXrj27HFYboBr4Fl4OACYMYKNIQ1Sx+HNKSdkrO9i19HH8k72wZFzjF+0cZHTwjK6wtVGQ9f9ZUm
N8PtTgjYRnuKcyDWPxlMJrU1vd4OvsOViVpNaw4+7hHjufcfaV4OvPv1Cveb/vzOKpesviBQK7M5
DZ2weK2KQLKVHbpw+xwTrjZJklCxPp1J2eSA4H5Qo4L0zCThOw5NmNo+RuhkZUorR5Spn7paOEJO
7YTu7gfHCkXXzt3jBUNkxrJJDmq3FNZzGJBScLjkbgqdsrvLxUiXdMRd/pYdmNLMMSRhR22tk2b/
bQ7MpVHbm80ZKMUSHClR0GO8oWd9Fi036NuS2uLB6CpPI6/un9BB+oeFZv0PZKMR92Ox4krfALZo
tqKf/3Iw0X1LXlQSD/ndt2O3iaRNpvpkoozZcGTh9PSuLzKLLyngudocP7Og3WN4b5AzDJIZdidq
JSeCCf8SGm5IKTdq8VpiHDk7kROs50G6ZSTBPbU3y5kgUEjP3s2jvku2XTFLTQmhG9ovHcrwh9Ra
WbIZ43MEJ2FGfLGrkvCc5RF8PLv2vowBieAjjjFG0qwsELraAUcQt6MxAEkj2JiQKi7SfyVMym3L
/msdFvhnM9gUzBcFzStlbpe5UFpQXky9H3e2BUUNldPOz3k11ytJxIhOGL3LWskpt2LKe9xxksne
rYEI83OFVuYJytwKnbgveUnHdpvRwQSFLbxvOcBYbxc/mfgioRNMAXMwzX6MfFd2wajsftitmqQJ
8zhQnSduprbSFwV5psV4h2hzqL2B3PsBhC+u03qmrpsZFNr2SKHECjfqUbwOh+mEagzNVl565Rol
X1l1Pnm9n5cnfKIbNpGwalEU9Q28Cb8uBBRFYrzrq/pfl09QoUniCui1Ej64n7ON/71bHOwvpyHu
HS5/g/0u94gRsRrSXy8wtdex8JPeflXZQH/ApfPJDov2Qq8WKsHjb+a8a/c9Q/Vfj1AvfZb3dVu7
92KlKB3FyffiT6OPP9MkEa3P7ItPBBeczUhnuQ8BxuDlGuH65T9BzlIF0H2NGmyPXAynqa5JnZ66
f0eQCVVKROVTQiSfFXqzgswgwAhsqOZU7jGGz1YEP4BOlL6RAH4MFuXrppzSXBouDi2HQJomSXVM
W/r8DNskoNrOTK4A4VGKxsQlP8/02uJ3qa1HrBdGPBipXUcjcQH1chLyS0/NjeylrcE2gTeAUfpJ
HePOXMg3JbZk/cHrvFVBh5iaM3Zgzanx78R5iBa5h/hRW1y3h6uRVHg69yvvxDujAnHtUqwKxWYk
kfLyDhl3manU3GzXJo9oUvKoCZpqyldowXQQfC/xdAiJGf69cbwsdDvoMASvk27elNPFp+G1fESA
JnSdZBIJfBk1x4FE8vk0Qv4LmXnlaArnNekDr83H8kpAbAy9xIIUv8yplnMbrPVWgGqYXPxx7N5l
bIP198ygOxG3yQ4+Wt2raR5FDAAGmp9Nq2gKU6/1DMcHq74AHn8JOisTlPWSB4N/quo6WsMpmKzL
qMtIHfM1buXFtV/NSVmLcEN/wiQ9vo9zu0P8zMVWya7zK++LtCdZ3sCf8rNOpiDrtKeFfj6xVbTi
wRIWDEP9lqtRWXsAEmsv+Js9oeC3r5lfCCQ2orof3dv/PaA9I7xBugBbrOz5OvzALZTkYYuPoWsI
NaDAbMUSf58YXc4qgLXNkPHT/rmQBWGR6pqejkOAOmRNxSUUXpCCWbN8lSNNUhx9eLk7dvtN0jPD
91qFp7XPFKeGGeSi4yvtCDOwy34Tlfsei+q4N6AJgGLptMk4LkJLcMPbwQWSt7FtIJb32gYY96SO
Gkd1JVI1oQ+jtjFknDBrVPfgnppL+dYS1tlACJ5MmHgHH9pNpePdmwera9GjBhTKVLLBR7F2EXkQ
rA3a5h5MSaHPgaf/KaFUBkB7SExmwJmGp4XLKpIVfDsKhW3E6gtf03Tzxwbq6/qpj3H6gpnU9AnI
H1fix/VskaOB5IOFW80W64W9752qiaAr5O49ZW30VSuD5juHZasOFgWwvskufvid7PEsWxK24NWP
aXOpE1/myzTuf3UdBIOAbCvpkIu8ZwE8P94AwAh5UdHT6nrk8buuudPzj05VYrEYNS6UzS8rXmwq
kFdkTS5dr0ZRh+ZSU/oZ/4gnplWOXzMAVRWfzGRAYU7/fJTDv14A4+aY9ODVCYWE/HjP9Kxax19b
QjTzkRpmxaTP7G/1k6SqX/x2UQs1SQNvb/VGLgAgnuMilJ0IPGCcixT7VZb65EMiDaTlJPEDKQAe
7bdCIEZcXazKEE5DWgC4wm+Dor06o0Vs0Sg04rdAjZQPni2URlyeepzRsBWG0f3LQxLlyZ31pace
eFKGx/ppMjOkJgVpki8bUK00Ze8YNx6hBUDet/eIuMrjjnWj2kIt8qbG+mTEEzpXrMPtdgxi/jDu
5rMMLqjkjXH3DwDXRabm+5a4REKdAHcQOQDRuThxl9Ou1hNYCiFHs1waNZjRSetD2wylfFLEJy8t
I2dbyJ70FKUiJ4HkAaC1ydTpEEVG2bX5G3ajEiE+lGN18Arx1+3paplA5E2qUaUBhSU1WzcrvcXt
PID9M52hOKFXQG0lz3RkUhzeNNFZ+a8wWSJUFjAvOf5pMWq/uXzpEhkDtjNiG+me4/OKYGjoLn9i
FWC/93w5jiD0ibL4AH1ggpq/d0nppqKP6G+madkoUdm85ZEmSuwGDoL5pQzH7o/5Ebx7iIziqqXM
tx7L1coy9Px621egLlaObq/lac5ANuOz+a68KEIKoHFeSjVz/knor2jNWdjSy02WoBty/clb80eA
KPQlLVW2Ve+wZIyiODlmbNpITdRtSRz571DiUQjP6G9TpWoUJjdzSX/jHXu1UmE+2yfnAp3qz8Vm
4rM+TErE7zNxNDLJlw8bt7kTjn06dZYbVUvqT94QoNWRuvZQQuLE8We3tZoQQiOc/td61cz5M9Bs
i+xvsID+vlytQkjgDJRHTcLguxM5PpvHG9viLiayk1T+W78i0T8Tr+DMoUKzhCvTO+0CiPu1iEbq
1qkH4Kykxy1aQNP2ROWmDeSEXEmIXdK4VeVbK+yduWGXKb9miXbtAS+cG4t+DreaK9+hovEQjEme
/nNMAi8CWrSqb5jCGjEZDv8fKYFi3MY1D47CzHfvD1kQwYrTibmtnsyVDdE7KejhHfNpI8sw/2sW
8KZngAsDsNkp4wA1c9Obd88mrZ8xZ5oNxE1oJ9CkyrTAJ7FTkAahJq269AujyIYOHyPkgGTeAJw8
wm1paOnOPDY0DfBKlkeBBt/1KPa9KKHkSmyd8dicfc4HD9i4qFQ6kj3+IEfOqY2ey9Xd9rrHgWEH
dU2UdpScn7JcEC+44NkGX2d3qxmL8pf4yjqzFXkqndDxtETUcjYQN61eyaPzuNyBew3NvU4Exr0U
Yyrh602D2nzqXbJmHHpQceIF5Sq2arPkqDt5xQ9vi1U2ECYwcpwwYVRmmiTNMSAiCAQBwuSVIk/t
MEGooQM9CZFjJaXR6LytBky3qqAA0fEqr2Y++k4wyUe+ZOrAEbU1e4MxbbfTTXWf+aIG18JJRdGf
cURAveSBWfLTvP2vYXGspavCupYOGZqaAFGo75V0JKQvCpFeknT5O/NmcV3tT+tCIpCdVWL2DR9H
IQHeLK27Kny4AIPIF5nlvPfXCOAa6AoLenJS6Yg4DuM/dpg5gyMl75/plKbN607JcVamAz2ggb15
hfscP22TNEppG1NtlVPe24uk9e0ZEIe/ONk60Dyq4frY8uceUAtEkXv1CqdbCbDauafzKjmAvnXM
iIjme8IZVrZlopSFr9eksUVYwALTKZSwfZCR4S3wGNhlYZE52v1Qp2hsHwt0hoPNLpjGkUM5LJfm
+rOJXsjtLNOZLqnQa2BCRfXlWfNGnj8Zs8mIVZa7CvmFsRZu2owPMvzdjm21tko4R8N3Bxm7wAJz
1a6JwsSWvK0Hsi9x3ScAa5cyk6hlcuSTTwgv1M2eyLqZpJxisPD6IKRaiYiBhy1Z+/7mpvhd70g0
UIA5vD3GmnIA60BUDx9dJ5FSz6Dz9wZrCM7ppNmIUU3WZ7Vj7lWDPewaVpQR3tUc6xfru0Vekv8z
p5KvHVF98NGtwks9iilJjJFiKacEH/enQQ/oaRy2WAQHIMJwlab57rVw9VpYU3iRgyAMvlxcL/Zb
LCcb+fcQCm8q8fixRKcS45VjEsGd6ohIKrCktj13IyY7St3X156dYV1qIgSo/bupQ6BsgVRfwYUX
6Uz/mBk3UdHc2dXrl0ywQAnqrcKIDDeiSaLHQBixR0DWWdLGMLea8+st22yTkHhla22dgj5rqC3h
/opUgIEQeIzDi0jx4FZ4DPfcuTLTFc4/KXwj52/C4ClN6qPPFzGU7OqxMMYX3D/Kvk69YV8+t1hy
YlT5JWKO7ANFsq/ue8vkUmanzacMp05PyzVcB8uuPa+NBHNhpiT6r/AL3HCrZulxbxlUllSH0YXG
8lmzs0PTAqbnL1FZXsUVzl7NFblibt+zyZlP2YNqZe87csMZNEg7bkYiU2Zu8avCivLGjRZ2mDcJ
Sezjv5BpYd9OOuDNB3GCkrgojmU3s8LMVEW9i8GVPRJVAocJ4jDC+tXTm89T2uTu8hX8Fy3x6JiA
1O/8aEzGxQG3jarno4PKAwTmADxPXssPUmydnn5tpNN0/6JmjCckxn8NFO2LBGosdJcgYypOeceZ
cOuHsCVwP6lbRdwxMHXDGzMp9DklRM9fbBJ1fP687ZjzCYa9o213UQVwI3Vg1LyBE4/GooIl7Qmd
U+HcRakAGVeEdK4Qcq0XEDg3g2Ab9t2GGewNmpUnpnTkQ0/vEydJV/YksHiOfkDogUWHD5Qxyb5J
setFgZ0PBtI3YTG7ACxLMBnN1wfnC4jgjI4Xy79OueMtE3tYzpUqu90xARf/uocq00ELATkCWk6E
nfTXdxVZLaRgz3wCYAHPTp01lBLbwSACekVjevnb/UH2UiSJ9Us/dkftSmrgmfJahLzlA5/Knhx/
eS7ZK9EFfLs+LFIanjJg6j2KSCT4Z3iLkty4SFfijerueSKcdHM084A6RASuLd0eN0OZhEVhL/UY
RDByOZaSFKSNVmzCZiu3DjyLPEOu6N2iGfm66REfgJgBaZpu51nKY0xdI5XSPZyf8MUtpQFQOwV9
tcSFcQltRAG5iO7vr8EC7XoULiko5awftmc88f877Nj6PtM/lx9i1Ev8c6HpJo5nt1l5s+LI0x8I
Zb9+jr2L3ed328Quh1trmodH/qUAbMpQIZLSW1woN19kR71YJ9QdNblBhl9Ppil9/GOTT0ls0ysy
63d0KWKWaDXdKQRBY4l/XXzgE2r1Z2ekg9SzVAuNkIga1XWZast+rVe0LPpVVxYZuOTwpxjXkE5D
GDS7pvO/u9O4QrnIH6UzLp/r73J49v3Uncf/ftUI/01U7BYi8V7aWIMuZxSp6WfE5wWXGeewLsFQ
XIjPIlWw6tHKGB16W76Wzzw3vnHAQdf7Rr/ZzD/ShWTG71u/JBFQHBMRNDukOyfwnEsHtvh7BVN1
quhD48PJVdt6+DzWX7UoDyea/9r1o048NYUuC3dOPxUlCSxPNj0l1Dy/ZDGbsZo8Ub1hDlo8kEe8
edJDjDoSR3zRJqP5jf/+toq2LyQBreLiiX2OeRq9W0QYuNobGVlhbJg6T/CTLkBk1IoYwfgTZD6x
5mmw0LBlVEMPhkwPLTpmQeZDyAaq4XcpT12YdbPxeUzzgn3GOy/lJJZ+dkmfnrYZ5XbSIvWVahg0
4v82MVVqRA2O4yAb+BvJMofZKlL0qW1ys7tPVL8/RGUd0miIwtt7S2YcfSvRffouNeDrN2TUhSkD
lTA8Mq4PUQhywoGM5E52KT12KUywtgu4vVx7iOp84fAZt7vGWQGvlqeMONu1sxjkvEcdG6DPNZ8G
TOQN2oCXe4fDlm2A1poKsrWVY8q5P97XcMzZilfS0hqy9G/0ek2kyO6jCpsz2aaMvt5fWzCbPVL2
UJcznx5wdVzeWd48aNrUbJ4PCe+Vay1t+sDjvCIV5E/e5AHuezbAW2EEBJd8YpdJ4bQGPAcloUdN
psdeNoiVbU9eQY1ZcDVjWi1e0Z09iEQJ3tim8LwHNe52JEnAVzE22gUsUjcz4gS2h4dAXhBrCj+b
ug+dd9BWxh3BHoXovRXBBvl6oqhHGsXI811vjFMUx3h1Dbz781AK1qREx/JGFsNBz3hpatwYVUSU
Qlx6LQw99uvxV9cEOmshuWiVHlE4CWX0/dtCAUFMIWFvlAYT0FIXLpREj5oyg9P9hDbCgFJrgn97
v0Yi3e5mfbIzD84KOeqCGAELEHEuLmJvmlem0WelylX9FtTV/jv0J5VeREidvd35ts0SP0iZH3us
CgIF+tAJyNOv3qqYWiLHqofHRXpcdnCw6gOT/iwmYADPDa/uraQ7eTpQ2uIAuIqyJHn+txRJyn1s
9uAr+NdlrYuMGHeYPknx+twrBeyXNNSnoA1rTai68gnY18ebqk/YvRYx/B0bf/CY23pBkwxG9zTr
QVsODjBdbqkf1rmtv67xvJUivaULMg0ObfoQ6aRnvaz7l37fdJWhECYxqyaVl+np6M9SPvMnpOi9
pN3i1sydukfCSuXFXRdPhN1olH1udSbTK6rXfVnWhEtmdjIlXhRmO4ox8LkAgM+yrP6fm47h+tEp
PlUHXD5dowKb0lI9VFex5rBePcmGrJ0kw/XuN+W8w2VPXFVFNiWCN7XK1UR32qGTRVT1OasZGBmE
C48j/vYvLRQvrlMjpsJOpV1o8m81+edazLDygD4J7QmblXRe7KLGyRAZAvBEvYSV8s1F9GLHo/GD
D1Qd3jSeLaGZOgeH0pd4Qa8NB3n3h/pmzgaXWEDvp30nAXMZWGjjcFjI52dgX4/eY4CrcMP4Sc3H
LYUSTmILpCrzdaLFidvvmP5P1OaL1Jow8NuLTB3D9TdRYoeMHqo+GuzQbqQi4jhzoEfWj186KVQG
CuxIykmfQ7VehgntVvozWOmVP5cLLhIeYd5wC2sg5i6OdL20muVOa5uyMJx3ygqhcmsAYakeO+sG
hcD6KQYEu+V4vRIag7DNBoWe7XT8qZE1wo5oNRXu0jR2hXdLBREarD40ci68o3dv4Z3hCYO5HvPZ
6fKHfYyjlV7i3kjOxspkUrL2oQ+EcsbIGMDNBf8C/VkGN/bKSq1jN0GLKhuNYrwYwqgIqHeHGdt4
+t5wfQIH5Mmh6Nh4WR/VQ01FT5FBko2dELn9ZrxPNhAZWGFuukRRdUV6nEjgFLozVB+EdgzM6qHG
WhwxIRyI22U5pdN4bev0iwO+Kmb0HiMhRt6PV6b98KNVxQTtBMANN3anWznwQB/vTMkabji5KdoB
Vw9h1l4GVcoEYGfei+24gkCbpOZ/3mU8b7R+N5Zl4nWjvtEIri5kEl5BkuxUgzviiHzNH8GqcaI3
3HxVvWYuncoR5kEdfdicw6uc80AYTIDWvoTXelJN3Y9AEEJKvVlb2/OZh3C+uCzcr3pv8Xp1N0XJ
vzuBBAw15blDQTbLKmEKL5zxwwR33SQmyIZyEswlPgChJhxZKewVLm+ZftqR6cgH2PMOFxZ/aSOr
EU9IOIXU/Q0skkv3u/thJq5jiCyDhF3nxNymWlo8BJp06KMvd0f46cZUolU7EZ32FnekUtfUyCqE
kTQiv5LIBkBT4glYKTIam1dUiG6ioLjm/WELm2o+i0mAoAZGAmMw4O0yNPfY6U3iZrTfhXZkHDwj
TSM2HJUyl7tPTpCouW+nR/TunxMPY4KBXpeA7+iHXtlHCJJWYbdcZ0Mk7LkPdst0OHZrNy7ASWQI
HlYJv5tVxByqhZZI6auauos7T6cWyhQ21KVFDB9SseriE77Dm7qnuEsb+yVNmfATdjmjIqsJvqCQ
KRRKi7+frIMcQ+0MTxSf3umDF3yN+eGqG4K9xiPNqfxC7bm7ijK0viUcMqY89FRvwHIbLrip2e1B
xXof8srHADnmXggYD1syqxf3Ui4cDenOCI7leI078asQdD3RGh007LfmirD4R2BSdR3khn/lEjP9
AAPNXVbHBKNyGyIqXHgMFrz894x6k5GnipRen/RKxH+ELSwWz5W6Fd/1nz1B9lN8aIKna1SfK/OW
Lj4FC/fozGjDeKw/Upj0J3gPKqw/goKnY7sFR3ieUDnP23K8L3o8qJEnryXHvbkhH2ZZNwy3G05R
CVOa8Ve5ehFFerqTweWOILB37Os3xw9J+55D/rndZP1YYjj+WJwOoZYKL4oQDFQGH+xREmAkKxr6
FhzAXE1EtbEqDQmX+2JwIWNVccB4YoGYRBLEIdvb4in3L4OXy5aA1TEP2Z11yIZ3YDoUfirsbwS2
xBvxmSU3M3VhRi26IlPbtF90sIB0sniHsNp+SyLNsR+OrsHWizQ9LDTmKiGTL7A14hPP31ikAS7r
UboJoq7BlSLpflEonAtmd58cTAXcZTKrdvueC32IMEO4gPbvFI+B3RNm6u7yYcWfGsmjLnQwM/D0
JYOx6o98ta1seMIK+yJXXBNv8oJE0ZSuE7IqmPgBu18mZ3ufAXr7tsvU5zcRtSNND9stTaSzyAMa
R9r0FMgQPjYfgwxYa4qLbowmV/h26U5fgsq+XgTjcIcQgCexKKpBVpDFvsDbOViNCS4P0wrKnMLC
kTG/+kwcKVSCxa2lvRi/G2kg9QwJqcHSPqtsRXN4GB3crNdInlcUePQM22uQpJAcmcJa+XuJ8xgM
Oo9WgRe7zdX86thYzPfm/Ns0gQ+tziATtL+B70xwPJ8FVbbPfbpsgUpyvnI+HnCOUBNVev6X7S12
KWknv2M4iaefUyDUmYVGjlbJv1MssLnzm6M62C39ewEOkIYwC7x5nGXJeIlpd7mwaVsFUbpGigX/
VPt4sNjDu6Oh5aJqeCEYpnxtujl+yO3odQhsxJtstwk8EhgRIjaeKfdscU9vnnqBf3OEyjAengIj
AwmKo389sIkxAzImEf3P6HciaO7omRVndGTNgpoeT9DTC7NSoVt0UtYL3Ld+aFvuoOcpFGVMQF+I
iC3UodA+bEC0L2v5Eo2vC3C+HerxDi4dQqjYmsA8qxt69Xp1MTTfJYMsnqyldiNtD1l04FeaIgQK
fmbcXAKhBlcfpoNiwg3/aNnMQxbqMl6kk/QroQgSjHOamiKuTgz+tAa+/W9/BUsDSDpxi8Fc9nLi
DBdDlERwL0y3OF53p3BHnw4KYHO+fPaY2zlYPLrqKzzYe/6bgyyzvs7Ku/h4BDLPff3PZ2KyYTu9
NrLWMtdbnukhqbxqfyZNXr3r5OrGCSSQAtu8TKt/82XsGIHXfthp3pQnUp1EIWxswH9s8Uowjuli
Q40t7/Wp4a+cu/CrXuqsCxlcqswvgRuNKsMZEMHAo2hGGE3z+QT9fhwuGliT/C+j5bUaR8pfqsnx
esXMYxmrAUcZ7XKR5H+iC65bSZGCjfjcgrumSpBuli8+vRjlGEL6N0oNPW/SC27lukobBfGIazQq
d+5XQIMwrR5Gpob3RCSLHtqR59fj4JDLhkreYzw1J+AcFXC/2zAUtP5pLX4X6fd5dPCqXBbqC+pl
ff0vpGL+4H4q+o8XO61i030mijQzFHY7U3e8BX+rWx8mra+yN0OWrm5ISoHBuBsWKssDDkwRei5n
qk+Hp7irmjAKjQnan0CF3+RkbxSFeL/6B6nBMt/tw1XguWDtuoBpdjPKuOAntXHPUusk17fwp0Hj
pKku0wyMTP2UvY2PscMbKTmJOzv5MnDdIVK2YrH6nOH5+YQJvvE2t+cepNf7kKAPX6UMIiqFXjhI
+/bU1ttgtvJ/RvB26SEb/NywtHeDUGZwS3YgZe+tUXevUfD/FjNAuwCB+9M0S6ENdImlHkClYC43
AQ14SKOy5r3G6SKS+hMxZyyqZISfiockR5jZ99cF6iAHZYydUPm3DiPJSZcNW5u2EVl++V8lyytI
drmVFS0MKodn4iD17kg4Ip0G2RDuHkaZLfVgbEbsGY73O/SWV+blQrd7bN3b4yz/oLkO9LKcd99c
eaagp8djoDlAsmwryER3Y0EMccXr6ZoqdE/AdeZGwD5osnzwq7buspkr6oq2PSOLW0VAZdd95SGe
cUTzz8uaLnaP24Jqy3y2qeIOjcej5dKlVO0tBo7dOKH6ruacf89oWjx8M5czORihAqyN02gMXnEK
2zMpEQnCGY72T4rYJ4XuK8Nz7LlghLp9CpZwqaiS0XQofUeAAFq8FKFyMZcm7+6QIoj5zcx59aeR
V1nswbkU0toDMOUoXRioEiDHa5E0zmv3sJsY4lJQfOM0SH65cVlILoLun7+N87t9D7L/23+9pTTk
q7WOeksphfKhm5wpdzUSwFK3YbcOGB+uzS29GJpj+auozRUVFzhV2zurT82OW5P+uWC0V07CRlyU
RmL1GaNfmD7Zlx6YGNfidhHlz1277p4mvISR5rY/AmUDcpY7tWYo2nYwYi2/NPXUWNRpXFKS+A8o
ChHT1jIL4Ls4lUHi0u85LgpXUnqAEiY7UOwKcI7vwOpG4bIqrbTAYARfwUfkPgE6tVaMNSgVfgPv
3dgxQn4tFsFDqgeJeYcgePkIgqjP0JyIyWfpN5rF1bGzFVcAk0XHqI8bENmlPkg5w/kyYnWLWYww
1uD0xnJQHgc8pNGokYaLu+QQPV/6xyxhHp/HgC1mVLv9QpJ2MAgTx9JjtYT92u0xe13G0DgNtGey
GRnvlYwjIkiusF03fGQxiwyRiODAIb1BEQYfzrGokKxjsoaXM4beclyySoMYCQ8pp66SU4oPOFgo
QfRdfCGteJyhZt+a8g/LepRnFsPgsN/H/HE40pvp8ph25jrYWKfptcMTGm3teSUVAkWgyiOIQhsv
qsSyb6n+/SXnELYpXttHJHPPQNyEKyD5QvtXX2VFi+u8QG9SFVGR/myi9/gViT5DXsIODhgAU+BW
kQSlyD9VHTpR2Y5si0n30SZh/4c1QGuXrbMHLt/u9jwrJbairG0zQaN7wK+a7izNllTCvhLeAon9
VNSFFzPmXck+KiYuo0HA06NHKsKz9wFloqys/vhEO6RXvQ2qdRjJtnJi1esCvD7EJlUdfweVrGwb
YkmZtQjKkAbCTuxq5+uSttRGlIzJH22crgjmckCC9ACEgzmI4U3v9X4/BCBflcdt0PQEvPk3fj4J
NZQkS/H5gxWfzjpZp6MRT+AB6cnEa2DFbfSnOtJ2RxkHZtEwI9Nlwz5ZwNufhqy+wrVOBovFZam+
nBxPa7ae9G8+a0ymLSHU7GnHHmgNCvitaRshZWCRb4dp1HOX5xO8kyxEUtMi0f+JY+Xzl2pnYyEu
/n1vkWFgn45eSgXuiwSC/tae1YfevCKMIkjCxoleUnqUdozdEhqpxzjV8uMfzs7HavsI7pTO9qb1
xDpAndQ56nS8i9wXdW/oKH/inkY/CJyjxL9HKKEes5QRY6ZwC+7fdXFi62YxlXeqdxLFb+Zwr2nQ
E8CK77tpwqASFQbhBDzXTF/HCFZBPtnWjYhM1wgp5oncrYjAoBDh+DCFRw2JYn00IMUfhWAzMVUc
mUBFQwvYZoykbeihzJm09hd85Htkv1pWWOsx0QT9cBy3DBczbIQ/0keZXqgkg7tSiu+XIrbWC4IW
seNCYGy4hEDw0sy8XPeryDGvxrnHe+znOUOnUlc4wocNR4J6Z3F+xsgCe1KsLN1GONskTnAMxzQ2
qXCHLu7g2PXtTYHr+f/lRe8IgZEg3xOAZ3RIfRcD+rZV//aEeZBgay/nuNC/tgKhdUAgTxaNCVOE
B+8IutvSitU/+/1uUGx+yPMqBmU3OuuBifgVfNpEToK+QSZZ15BUvIdXxQLWB9NoVqC1Q5Cmt3iN
clGre0DdNxv0OeK722zD94UaX4Um6x1H2/5zIZxD/S7a7RzClp/0/kJRblVjySws7+6iAASLleXc
My7xJiTPf6bx/AsbN5jZicq+gY+LR3quCky/o0B5n6y1hlABO5bTnxE+WCnBQPcQZ1Ar+oRH+d28
zfJqBeKN6r0quzJLFIbGBuYXmGYF43scArgOBPhgjOcMD3UW5bv7GG3HpsHjF4YLasv+CovRLWXR
tlMGtcw67jih5zqUBEuXet3LOtdpZHBLqylCzRJwFBJfUVRsJ/QtNISgCbp2ChY1VAfKB2J3J96H
TOPOmC+Tpv2M6BM6J1Y/xuwrNIz1DPxgimlDuT793/EME6KEF2RcBquOFEA5GRAtO7T6PSBo92ot
F4sWhiSDevXZIbEP8LkezqxzCSW82OYTXuUr2hVGvTdhToIFXGVxT1xQ5kXcIH5BPOGLN3bdcA/G
6LJi1noO57UUFR6V/UxFtNHyGVXVze7+SlrfY6f9HIH2Xe4PhXzHnWjBLnvkxVZogE9bYhZYkCdV
BFf3PCxOtO+WHVkBL+DkiTyr0JZr18FNP8sLaceQO/rJz/ymRn2ggOCOqaW5y7zcXf6RfPQr7P67
VLrrvJjM+arzrm0Zbam0IO+YVq7MVYqCdJ/3WQvp9fhlheEK7T4kYCYp1vRXvw8aiPAuyZ7zH/Ym
8mopmX/qz/qLHpetxcf8rFqobDfIQQ0N9b9UwKmf7ffvSt+rT6jTCOaLpwuWSmCivDoJehznPMpp
gH/Lxg1XJB9r3Y9/pA9a1Rk3Vi2jrvYTovxUavA9+Vne4nVSz2KLiN1Yrp1N681PpK7ilOAZijce
6Kei618TJ4ZsiFWLhEu8yEI9z15qNjvTkBy8FZ5WW2OZKnS3o6t/qUCQGgFi6MtsETs2iXPc8Dt0
uayLJnCsr7+RHyf8N2aCxUPSE6R06NdrVUKOqPSqGDQoZmn8EJ5gqeMopPpEJXEHWSwcdh1t/ydq
cm645kCKmFrCtIGBjSST69KmdITuFlFxi4JEv4GPHcqtQ1yyB2GO5MVZrXUoi0WMdYVGvots5yyG
tApREOiWh8vlLaL2791Vlp5zPQmfYx/dRlnmAR/tRPKdaHflGMFuagZCxH2lBwVIo+CZQC21E3bS
rd9dbGimBdX1CDYPFwEXF7/Fuuf00iPQrBQ4Dxp4IuSb5TOWsPmh65Oqkm/7kktYz0vt4QMs2Hle
4rSs+BhrO69QNkbur0o1Pj2wVKXThrxVXBvcz4gKqwfnvetu+vy+fBoMeAS7Z1m1paL/ES7Vlt+0
looPW9CshnXklOxUyp0ir6DCJHhX9xOXK9Qb+pba9bTvSrgBGpsAIXf7B0Sfu9q60lM3bP6Js2av
83GyWLAGQuvs0EYcA1GNPgIeCYy6rMrpUg71zqwEcGDNT3/PMDol0NMVQi+2FiMVzHLOMEBRVeak
L4ZX/WhFmzg2tsav43Wf7hjdFGaQw/yQBBj+25t8WqiXpuqDvSqD72hXv1/ImQ8pthioHqwC3LVL
D02N5NcZ5nBAnntedE/rXGq4qRRPBdGN7RWt41ydfrD1q+FdI1bT4HMHYtOzBhBO0ki4vjch98G6
zGBe+/LRaJj6fVyZ0YbNTB2yCdBpNh4LSPm759KOEN3fStTmzl6mEo61Bq0zjt8DNe6/jqm8+B7q
o/5fu60F+rwcysQDpqSw+LOI5WqOezgwoJLsFhJjUOFOD3n9ZCYRE0TvZ66XL/G3hXulaa6042lb
zmz516/0IPQ3pWG0CCq5zPc3VSm3w4C3qOUw48n+QUxyiooaL/R2ZWg0tSDKxZNHl6lfeKWLswlM
b+4dlmOv5DhRNL9sAH06Hp3HAsgF6VBQh1vvrPsNvu224kRY4S7fLSZEs9Ho4vz04F9UM7sCDSSO
O1UKqsAdF+SHNNqJnXP7hNvRX+iW3kyDU2KJtd0ZOr+GGXuRS3dMkpXWLV5szE2d9hDqbSI4sx1n
Ng5jpr/iA5oYtRGgURs+7OEXUopg5Bftu75+m2QXJQblpZdzaOkimkIzXwtHb883ugiqUurQPK38
C4rqlpSYhSEpduC8s40R88iqMYEI8FjkvmvR4h1B0ugMLDi/hpU1OOk/E27Lv1X1CDgy8wRcZpW3
b/QTBen/ahzO3Nmtc35EPftZlqUkRC1rko5c9AmvNtT+n2bEZpS3RdUpA7OTcIYYYveHzpOHjwkQ
n/TNA47lnffYHlqPClm13pgYA5HBccfzcFAlMnZESIN8zX0VrLDfeCr0tqjbivdYBgnPTB0a3RtS
PBEaNPgDVu7A0n2BF/ExUwCfzms5tI61BAJxqixeQkotgnJhwvuiFASI1UwNXrPaNRgWxjEqCCad
wx+FTMV/U/qdYYtcKVDZNELFt/6k1RO4Bvc8o0/BPyBhCpHNl7kkDQm6cEc7CEdWRrQ9n46yx2fj
LgE0/l4JyvKkclgxm3MJmGAU0RUtHNBLrGopkTwced4Lo7wPYGaAyYADwBMfpXXacLVkg3pFKn5B
Fxnfx2vI6iiHPTs7S/5oDMANdDgKSahX0J5sSzKleDdln2BlguxPQM5vRjSfjYt/vEdS0w0i/VYG
ivnkxEZCHy6pLIHlUeZh1j+y4r7xfbUMW7GQP796rAgb6A+MAEHPR58Yf3S5/WKHIGh0tyxic1Lh
75qhDXR1y5cQP21ceIRcNOyxwstvzx8qaZbatsrfm2ep9ByRkQSBFgBDyG+WoiUs+/qJqzyq/ekp
C8ISLQ+dIMz8X3pqw8A0MTk8hFm5d3jsCafy4RuBj+bzP6+73RBcrAeSm/mAEt2iV0q1zDhcXjzT
hRmsUxYbSQ6fU2xNO+nM5poV9Kg3Ou4c+1sG6PSD353lC6dRG64jobHBkZ7WtpYoy7qd/icULvz0
IFqriaIlT1d8yuqksEIi3Lr5K9TPyWIUmmgD2STF7jV/4y5X8AOBlu6PKl3C+h3XWTULIQnjV7RN
oldhHddWLMYQCU22Vh3/daGmV13wCwE6zr4LTabOP4AV9bMi9zdT4BJSE+ykHT7AlsuYoAmLEDM6
zrDp4wZ7weKkchOKMn0RQu/P7NT9wGnsBBSI3oQFaOVJlRXQ7dZY1dJ9xJXhXgrhMeorGsRQee+7
yGLkdfB//iAfrDHdxCXZyTR5OA0OMMToqHFalezQgT/R+lMcbJ83jlJUPqrKcSS9lwag2XhKjsSt
/pEUcOaKN5dVA4xE2/0wh6CeBjdClm5Zbq7YmnLHbmmg+gD86ONwiGHnLWCnHNCasOI+O5Kg/2hA
tVbyGBmOtSYo8io11W9vyytqYKfG+6gHTW6oEQ4lfBmEU0meV5HiFsoyCvO0t/YKJDd71iyP56s2
/era+Xoleu28sfxYNcgczDEeYdzep71aloZ2gcGtuET67IDUGIMasnGnoFszbzfMV7xtPsjOkAEB
Jk9Ypu7cSvBbOUg0On1U2hmS8Z6J9RvJVhWp4H+PYoo7cA655PR9tKtLTtIqf9Hp2lTDMds1t+IM
33mE9o9g8McxqPfXcU5fUHRTj+lIBudHhkHR5EBYge9ggWQ//LpTy/Kk4/jvj+60yd9zJl2mw8iv
U3wuVWl+V76FwB+LKK5+c8ikz2+gvEPkLd/pCa0govneV+GYmh6w8LZCoCObdzbBRik7rZzCl2Jx
i1mifHmsrdQIZkw+QO42OOJHs3z9QHjQTChLEEXzNCzUDbURxp708J0u+lURx4s53UpzkdIOW30D
4RHc+87JD80+ncLsmeB8LYMLiOl4/hcQjsHYt/MY/mz6Kyc7ENe/Dh0hKH1WVrHAdOaB47AWp9Yk
WFzythbN7w9YAsIIDIjX7ijwY06BMkqFeHHtvQJ1S3X2BoKX2JzCZDYQ+c25kQE9NLDvGtsV3GKZ
pPGaUuDxozsbkfBZHz61nGGLGwKOfK6G7KZpS8cEFTstK6UuBd1MfUqFFgdldU6CVklc5pJCYkHS
VJNf74smMVPil1fMnSgZB9kE6EGz6yd4D/bE1+6uM0DO2F6Az4hKDYkpjF65iUeR4eJRDLzebtlg
blq4UsVvlL+z3mnLdOD+5issD9qJAlnX6fa/cvOKjH10H8SOud4/2QaBTc2nk4o0C98loK5DpPKR
/6oh/CfuSH/1IqJFHy3Km7SVVRT345fa272SjF/0uqop+a7WhFtDGlrQVn6W4I34bvG3gK33kDxi
Jpa5LKiOr32P+09n9iYl69jFSdcjs+eUR7a+43nACKddPC+SEOxLc82IOHwrZGyVxARBzp029Up2
ReESd5/B3ZoUwAYMj+uSWMH3RGknRH7CITruwsjivo5TTlC9ZqCaGX74OZZaQi9MhL2NyOKcTBWe
seei4YTVvp0Qy6z5QTHYmxKHA+9Cy8AcMwuoeWo2TPYoRTjE4mHWjRRpV7K86d/VW1XrQmLf1MIQ
pfGA+fdB7O9hEZMv6y/imwQ+KEjBhrOae4UhWLGiRatb4vTwDxLbKbRGTFEBBtcdKGtU2qe83lNp
evn5lmjSqgYdXGEi4Ik1eMDc6AS6RflfNGv1rFxetp+iWo80VKBU85t9wD1923tupn2DNRcwelN3
F3ciAQDQ+xTe7KqFwuP4fOaLA6yRojbMDVEbBGL52dgDPIF8uzOp1r4HFaMHt3s3f5RoUKvuZJ4j
+VMVPgFqQ5VJfKUR/1hL2TZbKiwZLP1DE0mctmnMRaIQpIqoOgI7kT0v8eIMBPRYyPecbzoryuFY
uFJRNC9A7rery2IfijEcgXXbnx3EZ3OGJyDTsppkLRWknjtFcZhjV2bF5GTs1yXceDmu+0D+CtJR
SwWDagMmZx1U5B7e21b2ZeKkwAnTLfS2XXKp9XVGV3y1DZYoANIpgvdaOI/86fEbSqPtMs/S9tc+
tOhwhPiF2npF/F07PBbYW+27S49KJLCIs9UEGN89yODKRXZ/tQZ7npx+7v//ZbD8EXYCT36WC/b6
r27Xf25UMpmyTxet+MSxVZUuB1hp8iZWBC11TCBuyWKsJ9A1j0HFqZb/PraOrexbzIzs5b1+W+GW
7y2Zd+YYalVCMslMsVVvQ0+0YxMkRK4stxIGEK6IUgPrTlM/d116Mr0R7I4LZsL9Yzzjeg83AZab
ABSXEuMIy03glSa9NOrK8f8bxsCW5W9HTuB2lD9r4wSWMG1q2KSh9b4mF6mjj4shK31U3y3iwgt2
cEOGTb1Jz2y9xrDb+62r+1MswA1aMCu6TU/uhokpu0I/GxtpvdU52OXFEVak/hcgLYL93RHzZPY3
p/7bOri/OZGR191YrCAVXaKtkPh2cJJLOS/IaVgzf8c80m4rhL3kfmz9Z9oQkBYrtYHlnyVtDECo
NsMNsL2BKNcerWJtO6bkYjKa01iBjKh5ol1sWzAWSNyCazhZQyU8TRzLxlbcvx/okYWeHjTZckEz
JnYdqM84vrd/0xOGZYY+hCBCzcmncOl6S7bDbiPaMdK7NOtaF0CXIbwMtryfWbyaCacwv5X3MXDF
e/UmHBbM/5t1/fDSDHAig+JP86G1me94ttl6Pac0ZS+47P+ATI6lCvKa0W6yUcLSJPoLKNGkW4rx
B5GPtUV3D9C1zbPbju0OlRuO0AX1nqDfqS8hT/PO5XdT4oVK4dCz+B5Qc533OlIrxovXFsyi5YV5
TdjkHMYKAyggcIo8Gw67Y5jdQqJ8Nn/T2+EzaQ84/6vaOfcrp00Q8LM62XgPGl8NpydFch0UfpKk
8jKq0tMqvt/R9I4dqNtCIMi/s2+ItNZzVXXa21bedw7dlUnwBwj1YOoEf9Et4zyE/F11m8AT/PS8
sAaG2gyVS/minlzhhbDEP72ze5dxnobMWVjmBu6IEUmooEQuBttR/GV8D38zKb4bgogSEDaovk1e
qImp5xjoXf1P3HbqwtBaEUfjYXQDTSoaWTiPhq4t++0od6dhGF6I5nqr78Gges+ucBeaJp3YmbGn
cj/5Rv5ECVjse+G0fSXbfF93b9uT/yMsILPfNWPVJG19PyoFOTqLlHvgLICAL8p1Zohuuay0eY0T
9ZZwExFFWf/tV+JuXFCDhYmtgNk63qjrtWem4VPccS9ix2tGlrOfF7GQitYruP3FpmHpI7zokjAG
fDB3NOqzFKMIzhSwT/+Mj1qoi2jdTK1TRcMuqz67yp+TcJrItNExi5qjX8UfWm9i7yGeOeX+NFby
PSiHky8zxGESkYFCBR6tZa+5FYaAGYg1r7aPn3uhzC7TQsO6ZzBaJQCI9RDD0xThB1/XiherrvXy
312zKdP+mQUZ1CDa2i0LaXKf1REWTlmK0Cp7EFzFVbkCqca/QnXyF4Z1XzNPpXHXn/TuLZjRH+Bd
bS4Dtuic8n8L5/TJCUWKZb+qF/yULdmnAvGHC2/vsGIzZqDMu82W6qzI5+wa9g1E7mdzp/JyqXtS
Zv+rWVjL64Rz9YRLNbfGB+7DvJyLu66D2nyhiM+6ZCBBJjYxNOJlsllLCXJZ8Ufc3w3l6/EmoVvk
3WElTlNikzuI/mNht1TRjTvoY1vSxYCFXqFaQYySI429/yzyfeaAjUBhym764R9b0Zq8HLBykreh
QqlTzzBlrrdgDmgQIcKcs73pCpzN4DJEmurWgJ+VLSK2pzPX/iR0pe7lBR+MILAy+6+s8QaQhssZ
tJPKqw7Htd+pleD/A2y4KmD6P33mhcE7VuBHvode6zaDtetMkviQkAaFIvd08BFGwniCvBWZH4Sy
UbfLOnNHDuTlL5+vbBYNZFBmF20ewiOrDFof/RGPhTsItc/lxg9e4LAvu4BHOaMegbq3CsEGB6PR
7M8qzThAp45afvqxuf+d2cF7kecfSwBOHglbA7X2toof4M1eDi7UAm/8M02/sLPGIUdyVpMZpPb9
wjOESqdQUdPcQl3/oNsXUYixYQcbL2msQgM6dx8WFqdvRgraJt5pTX2VLI2+MX67SqNxbNoK7UDD
FQirVDbgBNoiygvVQ2A0+SPMEnOKFPX8HvE1RNifDmaN0TF2OW7B2ty6hNH9Qr02xZ+BGUANFKg/
mvY9Ug/1ORvpry8IB38Z5nHR2faBUiwJIEzALC9fxt8Fj6CV+PDh1mCAoRWV4b2fy/HxFkjHqssK
hMZCAp9lxF36tJqtzXp1q7vb/D1bzSZLt1d0XiNbHqFks9YOyjNrR+6PmHSJiMwjPExBffExa93v
673Imfm3BB5+PXhCHY3MQDZiGtcOYSXHeQ+LoSiGPRhuMO0/VLYcHYzKhEfFJaSoICGemg1xubJL
nNNsZWkmXdkw1euAhNPHzZsxWabdNxI7kuihSRHN1IiR8GnXhm114tbeW5m8Mj371nSIktkdT4Y5
2nTzl84zjZbCnvY4iMagOsZd5j7v+Wlc902E9qtcdHxyndo0teIzUNQBFe1mJN188UiTAPtaebBx
Vt3Vy5mfU/EOrERk4OU1Nu9/EzxE/4IgmF3/VqxO+nz6RzQa0BGjcEcFNt6kQhLB/+qn9VmU4lXE
FLDn2A8kKLrbdfGqggIIzzRR8qBPVAulUSOiavlHCLkqp6blsT+ZrDxOgOZ28JBrqRk3N2viLk+c
NOylwhx1NDVMM6PezXoiaDtqWWfZzeTChyVyfJBwvKtDUW/bT4W4e7Uy4HEFN9m2n4CuYU02XvdE
T8JzoSSH84lupb6Kqezws2T625A2mbgCozmptxEmuDffujUTU+c9ZAbkU6Yp2KTjJDaB9gVjydB7
ucAF/iOJior3mZLkMREh/T7RBRPCVOaTDHVd49hm2OOV5bz6V0caufPuH8DhxtOyZlrCWr4KU+h/
BvNvzg3jIkM/nQCMfzVUuWUSTRKRBUBcA4pBJH0sNcRb5g9aItTevwMHO0iN4mxoGLp5Tp9cn8Cm
yP/AqwMpVoApzR81cYSrxrlL7B9QZ676go9NR/fzJWQmmtO9HYHBgHsP6Ng402BAbt2lHkefW2sf
g/SPKOMpoo2FSf0E+QPvthl3QBagvkCppE1QBwhCY3DDgMFPKIFHozreymorRzDwGR6K1tReICDh
fpITD+54iCh3vuRLuKv3U9nCT0v0e1K1FHMnJFz/LCvQzaLKLBUxIx7sKi49hUEu7ya1/txh1+g6
RbXH7E9HCanzH5vT4opfyMzJMQotK3hz3o76sWQHwJqjfKSC6zqTEUu7Ywzhu1M3uPgxYLz+gCxm
TZtrBimPg2TBlpoRRg2L3GFUv1SKMu/7JKZgkwHdLO0A0+USjkliewQMMRZvl+D13aUrl1NN348H
07HnaOTLRf2zz1++dfrdKHhjlbswdALFZoJxVi/rC027+5CdSL4q9vh0rvwBsX/PzCdmDf1qhRix
SgPI/NJi95CJKiQChirz558doCCmapUv5o6XuttoBRRcMQi/T6EyXowD83Wrf1y2bfLMzHcnd5PB
3mCD6LPOAzu/hnvYhuKt58EcwsLX8rA0r3mqMGWBvhOEOIAtzLkiadfihI7HtmMmhpQfSqY8O04m
LmZnFly39GIit6LPTHProezAn6Y8PP2hoRWzapti3BDhD1GdE866liAJj3J4Lc6jTAsVGabyw0tN
RIh3If9tD2A//9vJ2FyE6OqXY/z7WI6UuvLWHd9mWiCiqjocYFECLM1COtvez08/CWmhLsLU5D1Y
1Rlfz8i8IyUZuQKYknxWHLrnHB7qmre7h/T4xWps87VB+JamiSAr/XcrTEqTGSL3y90GtHgDF6So
kBfVsN82li8toZSJayVr8IBl/KpuHrqElnIEfFq5KUY9UjHiYZGFfOYK/qKL18XpAvStl68FAS/i
7zRr6JUml9gxBU/0XfzAGB1fK6w5wJ51BQ5aAyxHCE0mEGfIfildrzKS8OWNvqA0AGWEGOjtdmDO
0aqcghNazATKBVZm9+Vh/hvpCnFX4UNLskWj4rrvEj4WarFfeaH3agSLBUP6a6Xm7yIOjTNV1ZuN
ni1219yPWT3VlLbxKuk9OTHBIxMExt07bo51rfIsjdyrVqMFFS3qkn9XdS8xD7ddEO+GaoHkop8f
pg6kOtmo2qvecAVLmUhxqxDbsMjwRIkDf9rLTfZ01mZL3oNzNiCiPVtiiW+BdjaohQnCoirNOdpL
Oqypvmdce2Xtj5++WbOIFAoi6OMbfKBZ/AJ8rvIsgtmZFImOBXKPbw5i9WDpSt/aMREEuswy6HPh
YMpedWgu0QTduKvHtIBLbgHvkNh6BE9SaW7haS0HgxZN+wnev0E6g94ldg5HFKuMZXepno3rmXN9
+Hh1FQ852omwsF7soJOysVibOs+iNb/pB/fvcxxZOQmEDBD8hKTjAbiFqxvqmrFvpochNRKfu0h1
6kpu+kpEN7U07WywqBKIgTiGwzCbwiUyPkS7kBBOsVBpLuAMbKOTuJPJVc+dOQLd/5bHoOfuFPoo
iwOAFrmdKwtKAN5C/C5yQg5CIuUgJbXJPp/EjSrt+Z95/+NCgh6A0PeRoXyBpg8paj71M7sMvYwL
xxpF/3CGcYb7wfx02GR4Y9cU4Z+ILERtMcb3IsrqlJR2cO0qivfpxc++1CarPMy1aQItr+0DtW/a
2HIPWEmwvb4vLeoAbfxDOsNPJPcIpdD84VNMpnHvQQZbIs6HQ/VHMlaCy0rqUuITyStxEkvd3oJz
mHuBbWSQFnnmuSgQ3wjSu+h5WWDbSDZQYNStHFvetB9WvYmIFUnWk23cvrEX6wna6iGjugwUKRR0
jo2i+fZJivIQ8z8jCeSwrkq5vzXtY00jZ8HR+KTxjcxdgVLX5bPETOMap4I2l2m1Ar2QuH/Q5VKo
U+zWdjhUwvEeAtM6N+pyrxyM7sW6DDE5P8ISzcGbznYT36/3T5G0ma9b13Pbs3844Zo+lVuOt6so
ar7b1hdZZHsoHTuZI19ZC20ptHy0L/XVC+qQPSU419hX474Quf9L6lkpOKfRkhaK8Mihmban//QZ
Eix54FUchx6Yo2VV60UFN4dLigwYvqC5/gFu1WP8XnBSjkpn3IUiP8OSDIf6vAxARkNvRDEcmQ1+
bgWwOsYqc6RJOk7mt5uwqo/8rB9wourAtwCKYvlIYiR2EgYhPo09HDSE5TcsWJZC1UXZPzP3C+3W
bAYMM/navspwOdlEfaEkNZ2+MUpMwsQurSSzG5izpVoWJF4wMgDgwN0DZUCSEhU6HPG4+4acmFjT
Lch3PxfnIRmj1n5GexGB4lpPPTjNBf+A51XK5m6QJVEIZLHY8Mx2BvTZ5kBfe5zEUtDRYGmWfI3K
KaTYDMoYubj2qC2M46xJBBWMOlXLRBkv0vMZ+ucynh+PJUEzPJv4PxWaK4TNVV9kLAe0dQ0aRBaK
rshFLNX+ByNk6Znj3KklD4KeKjoUh0uDrzr4sN6i+Urjb6ZscBwf+k4LmNZueSSw4foIWPQ0Tmdx
DrAIuRzDrsbnwAundQ5x9uvk0e0r1dbssMvx4ZQqz9CShYGmkM53mSM6YMdhAA9GqwN2NYKiLhio
WqEMQxrXGUwCBtzExOhFotXHtqLdCOcgV7kSjgCaM+x1TYgZRoPO0FTm4U7KZ8EITmN8rpc5THR5
pWe8cooblTxSu+JctNaIqYHhncFmhGG30wxZX3doFv5wxl8hGYg/q335qEHivRd9yk8tOoYyHsd8
uU3fAn0eSYl/wN/3R7e161SjmcnFqlGVtwpgvZ+6V21nkYqjtAFo+qzFqVq2gOwSpOamHy/6LdGq
AAHutVZSJoTFd/uy2ptZKGXDiGUqa4kba9fl4Xlg43gjZH9Z0i0ilaB6wdQUzmElJd5qwHx/FKEV
I3hFe0WhF3zVE3waweE2BIoDLQXefauQe9D4QcIDPuUCvw3AdcbwYqA62USZDNCTtqULx7jQPrYP
J0fxIx/hkTuOaJknk2kkZ1M4MvAn+VI7uQRuYfnN6xDO0pimBIjU5nVFplUtVMf4AupxE0chpyJZ
WyI/wf7Olxo4Oyj8l8ec9a6JANxiiAVnz7YoRC3i1E2KPxZ3Zi/SCUULXrt9d0Kmw+8yuGVU+t3X
2Wvk6QewXhy0D2CLxfSbuYJYhQUlj/Qt8iz8k0/VhBipB+61b5amNfsYw5ZQNOjyCxc1CJAD+WNN
bV9SiNA7aoDTzeHdD9vZkbbR4bWWkIARGNTeOAES1M8SX88hj1FHLW1jL04MTSDL+uu5S7oNib/C
auiBKG5M6DWYb1H5X8VYib/4NJHhK9wzgZi18aHoUFp6ulEdE+9gE5DjX8DQtWrxFpFvLEvyIhw2
sQvW8XJsIyFrkNO7hVDyTH6Js2o+c6iscadheIQ4cC4kq7l1sFMgXDkPGmu9P7LIsMp3+2h+uIlp
mFhmg9pnGbXjZQ2q6q8NjP1N7wtp0kn9O4WmzYug5N3I0bUux2VHGPIv7aa8hmjKD2V5jSjPomlp
b2Q/n+C1BODd0q0hgeZOtJQjsEHMPjPmfjareXKmMO0UeYq8xJ7bk/il7HoTAMg1RUURMtQX1Nrx
M1AIYg47UEnTn/PmT4eFZAjJqTpSfm8R/2f1WChI7vqtUUyJf+cJsnEk8rBdWlt7A41MPLVzj01U
4PWbnnGjEOJ42McQvneIQi1Py5lYFPMGY7zNBwqoI+HCHZbHS6RsbdQE2k1+XzsmB+7uQehCMdND
tAejP0i/I7fCuqX36kDgLzawhs6HBMCVg0XxqirFspA53TCsNEhrWDftqsPzINfdMxOpquSQ49Pl
Fu24sLUnpNgQ9Jy0D273mAUzSG6ib2oJkH8VPgfcInlIhhIbNDfXbyBvG49jbbFZ+pj09rcL2tCC
BRG5xJvCp/j4JZEs0ivgyHW/7ci8uclIAyZLPCt7W3gLK7rUNyXbSz51YiGrVZrmvt8vHWYIJgVa
uQ9Odhpy19G6u3kVtoQ39FH5yaOrU/348GNMCVyxpB5OvR23bTXyVb0xJUQgq/lBTwTLvftsVEEL
N3o3SlUy8tnoqETtJhwVxD4R2BObLCBxVkfVz4c3W9i5nwYjKGih+5pyiwZJ3zy3Ze8WuM7z1s6J
xX8V9YQOm9u5muQqXA6G02LIw2X5cj2XubRsZRmtxvH50TYVsl+CVUwfpQx8LFBLlDNxpaHZyIRH
XrNvBGbYJBPBnQQEfjaT/UPvoO461QRu6dRV1tcy08aHrE3kCOns/7tOsk2OpshM/5bpaZ4L/0oO
atL9RsLwQTSo41gfgM29OaFeX6Ip07iHrspIdbBNyOu2dyuv1oSe8vjXWkOk5tmZYdcUqCDOKgQN
dBL7XasD55x5D9jtv1V1n4wuelBkqsIlAnQcWJe5Pkm9GxhzAnGjwYjN1nu5ZU+e/HbgF8cJSVpm
gOXuRMTpVvYnPVjJUlJwUHLrVn816UtBG6CFZTV9q56nZeXxZQ0qkNkA682eI/5B2JOjoU64BSNx
pVcROYkdccCmWusPZahlicDasCDaSUv7SsZMvzLeuawH51GWlQ8hlyQhPRgQncjsXRucDCPEB2KI
YFD+kE00ywZzHGUzO7+NKWatU2EgXLx98d+ZOLxM8nnuWctLRGphyAl5FLEbETOwwuqgfEIOcpoh
5f2gwA7xMx8YezjyVY5LbOegg3q2X+0Yq4PTMA7pyb921LaC8xy/zrVvsXfPG0lPGjJdec/L02PZ
0kOg0TS/wNlUPABpyQNBv6FL8/1gVkkMZJVIPrBrDLJoN51sBFVs+W5jRln1Ub28/W5ntYP8k2vJ
38CrQLG+REFvPcmQozd6nss6bgcLwXcPzrt1qu8v5i/jrojpnMegvfu72yZoDgG87Xdq1mT6OMQy
piM2nf+kJzdjLCnlGHqAdcJXU+hyCJ8fLAns2mCS5ecVlfcqfs7657/KMVFQHYUnncgYSoZVotcm
xJID7vwEbWLux/lNGU4UIyvRvk3D5yznr9d7CZ+E8FGHnLPWYMwGVWcYb9gkiD73WjrRKFR57L6d
6o3kNj00EBsgpRR12KV2tbc+0u9ONwh9bOFa8UKGHlWUqqvqAnNtd64l4ST8/9wiT0P9oduNZsPr
MYmBIn47+t/7YlJJw6zV1o9/oyEWDY9gHMwDv8cAX3BUcbXlLSHkj+sEdcEB5Ms9LLO9pcUGF4KS
IKokDSkETOCHFG3djxy2k25DU6wBFgK1R6dSWFiSmEUd5lFm3Q+TWLg3XnONJ5FvOZGLyLZ1+SQ7
MW8W2brngvPuPzsNw01Q95vCi6OILAY2z5vuRN9GMAJlSQ6W23KHcI+CBeZfIhP+pN4189JUzsNt
ekNH84toDg7KfzWzZVYgMo7XG3WrScuhwUQ617AKFswPVwkctKJXAPoBQZ97VYSN/iv+tjFMV1WZ
mXfwAafRxBZSmUKhzApJwVEz2pLxR4oluE0Qohro+riWTsDOW9ueDv4exvP+f8CHfdeBpJydG3I0
UIjAzCsJhVGc1Z2bu9QhRrz9Bc7HRnWnOrkzkbSVK+Jt1gUPaUTt1G9p1SGpHOFRB78oWwEKOGD8
QJfqgZxh8KqAtwLmLwReooYd/ZPRJseOZjW1eomRDEbLOVWQ+7vFJH/BXc2yohJX5rTQbpRGwDKq
2wTE7KgGfV1pUmAZbJZVs7KvDNT0zgNvwsyffI/zi1rZ7T00nYcAg22f5WbTMjvYeaj/J/03Pm/c
2MZOa7tVigzv1GqO8TLaMdwcrPvklbKd66M7G1OGBNLP4AsE8PCZTt4WFKt+z2eDMhqBhhGGrm+i
mkqMA2jtQj7I2LF+fJFgdkXM1iY7NHTKGtn2JoZdUypvrnZdEI3yFh4IkzeORDnlkxxs0CV36bi/
RbcTIJaNx0vUNPOQ2AK4pTCr1pWmPpVpNRQGc+wUCvhbXR25OX64R56zS/S9W0IOXRKr4x9j4kZZ
pExMQfmtKCsvn7qwtTTKnnav6fPuxsdBQUVVMhoESjtlR0r/o2L6TIazrTlVk1iVBB5X04EL73vM
sTGyKxj6YnKcP2MNPxpr3+thOURT/Y+6lLt9NviaM83P1gpnYA9E60XZ56MlbIjSv4eagXACAEbZ
R0hEKzghfy6aP530ZcrBWBAu/Z5ba/fepDxbKtziiWkNKflythx9Y/4GWxEUkTmJBhhQ+Reb0ND6
tBmxRSrVnN/crwdeAmM+tQWyD3/zcrmBKU1Kp7mjzuypNNx2qvnADAqhajbf0CnOPp2bTgtNqP22
if2yLQ+Ee5NeLgLVoLO/bsXujN40pi5Tl6EKSaE1kaF12luVYK7FFiHOGIjG2rAs2+snncq5KVr0
rdXr/sWF2qP5cnbbeacfdAIwqX8kSUJO8jWxRKtmbbahR6sO61PAtsmwsLXPIqmSmeekV2P537Ig
WQ5XKzg1LQT0Kya8N9wnufnBXSS9taahGc81MDEWfmPjG1WpCwc3w5srpGX7Ft8IKd49eX7Wu4WJ
1RDkIAr1epExh3NGDPEU/SIsNyksPA8j3xERriQWYV0iUcmUe61ONjbXSNlNvHqR+y0ooSJe30CS
rMii5KDqUdUSxvdBT2DBXKZs9xqZ1hc2d1/Z9LRHahH7x63d31Veqak3BNj8N8nQnnnaV3G1oFA3
W32w7VvX/A/GZvg/rr7S9/AHI5wrRuSOteCvgLxgSMdJMpKr5Xp2oeFIVv/QIdSbhJFVJG2Gl4wE
mEvVUYYjjUsVvVr+KgGCCDRkQe5HpWQWA92tT3nERA/SaBYHpoubbXEOKNcTT1KtllEDSGCXiycO
zaUtCZ8Ge7Tql4QijZaN9DbP20aDyJ8dPRZHXgm4BEZzVGwkXpeO7cXoHtmdLONjkfYaCMfS8tY/
/YdgDUrpEHC8WASnP7SFAZdtixuentNT2BzgaBJzywualIWmghADqD8yEqPL4zLs572iJ758e0TS
aQrkOlCLHcsYhXRVIq+3ZT3Jvvr2zbgnLKESEizOCA/HsJDMqt8EZPZfubjJVk6qRGawhc0F9GSc
EGhZXMjhkO8EAMZZknmb4TZH8CpoFdwM/IHhT8iAPGEppdUKu/Rm19D9HECdBgT7hihdIDD58wUb
H0VP5mcbUUpxI6E+ZvcDb5BLqq3s1XFQ8QPRkXuUmjSORR+a41QW9CyN6r+p9iTo2jQgODwn9AGg
vvUANmdT5Gk5E7HkrC83+C6+AzvAbWVWdzkUP2tgk6mQlfRpYPYi4Tgi4uRSX2UounFjrvopB5ls
NlCq4zju4IZ6K9NTFzSgJ7yDlGp0R1AzA6cC63gMhbpMB8JWwkor73KzswtJFZgvjbdGmofRHl1Y
9PoC/NPNVEaVwMlrHQiLjfB8gukFHcMqioLRMGPeHwrbEdQ//U1RxC/k8nvkk7pJPybsmcFsgQVZ
agZuShlGFpjLejUf6uXyFgKPFf8LQe2o4eTPVRX9fOT7JjhaaolM0Y584syZ+1QcbFFOBAvUhIf0
taa2gz32XBgL6L5yL2ue9Dr8fqVqx/1ig08x81MP0Yt3M4O+cAy+mYyrw6QJQsY0EmrMaDfXz/RJ
ggVNS0eEkJP4VQVt0cTv7dmxnwszmdi0KN33vaGVOBrXrMqeM7SdBCnYfSES7yt4XBmNTHYEUuX2
z11JMYjro4ymjAwltEbjGbE7/QCwICNzv9ICoEAlvEodvmn7N9M7cQ1Zo2sRJGPgZyg4jhde94y0
Kl0kzcug1arc5maXypoMNMNvIUEntR3NFvl6orn30xEGjF4fD/UqCOEaX/ppdOcA41h6LJ8Ucemw
B7LbJBQTQJs0qFOgb4qo6dPvILJLbfE1gNqXGQP9F5UjaFYhF2/N9qzmspZs/CwZADSNVVOgIxo2
RNiphNttKmVKYT/HCjIcXpxy+0dZ3fwZ4I8BRBo4sKWKjTrD24gkdAQIiw63Joq8VDxvcZgRJjBt
xCEd/XxXH53EpwmVtYcl1SvyjDyhuIouyJnkzA6RVxecoVOl3lG1F3/14inFNIvTgj1ZoPx153Le
Ti2/i8zjJI2jbI9wlOfwDqqx6ESzIkZa3d1GerPVqenTZzO6F9xLFOQvl5t8Eg4I9es0TnKtoqez
6B3oemTfgg5fmkr4r2UbDGbPrI1Vi7mNREwA/nFkY2lnsY7Ln0k/lVT20upG0p9JustVyCxsI6/q
tg37dKM9VacEquRAATs8nTHfbjOPgXcFDvbSKwFfFqxkxVlC/t7mWct1O7t/Klq1CKy7IUEQE68s
9tHOl/A7Q5UODG9ux3mxcD1lO6fq8vxLncUh0+DtbyitolBgsxMykmukMAyvVJvWRvLIPrkXAX3S
IbtsQsW4J5Q1/fwpPQABmqjIxX5Iq1VgkXLjiNH1gdNPz+gaBXnWuUAHNvsAmDV1Tm1yxHUxv0xL
HnqIsFEOuJprxnOc3Q9gg0DNIQg8O1Scb707Y7beTlDQkmIdPkhq3qIvgr/b4dmIcwVEQX641jnv
+4gc2c53mDrKO3QrA+ts5EBA+bfAORTmu01Fo18cjvtAKIa9TF4yXDSA7H2xuBVGYPszI0Ha1f5/
HaTyqrHm3t8OYigjuqgwHMF9E3qH/iOOd8IQ6Hc9BffofNVDlj48e0WvpAPS29yUmaUmWVNedvNO
HLjlqIGBNZMS37Hmhh3f40NuIuueefaw4jqaqQJ41CZDbc4FXv3Sdr0Kw8jUGt7IexgElEjiP6Ew
U9o9tlOUAUOU5YrMmyZKoGql+6agPErTHpZw5GmpJGJLUa8fero8tPFLkhm9tumHF90oKT1QvbDE
eLBYF3iRnefRbfJg1fO2LTD7rlYwp3Bsy60m1MFa/uDWUsLZJNU8CrfmtBhyDKC8KseQEbZTLsRJ
qClm0L4HQtZVNf8jJdw0oC6RvcJbwD/68LwGW8wuKC0crsk/0n78o0ysXV2kgHZs0MzCv74UFXJo
qpsTqWIBGA8nZ65S5gwhqrdgSE2R7Lu7HpTZhuSK/ryEVeG5bpCpqyF0/x0AYUlmhkYaods5CBUl
g5yYInbkBDgx2uciCs0FVi5ssoQghVC14Iw5fXqs7ayxK/B7IPYnHT3ZnZTWM/jsbWxmAsdQsypV
FiweHWo2kVg8u6N5VP9sjzKQaEbSdhhOibEtGcWg5k51BwI3uOAWdGYztvBqGPNm8yoCl9N73PWb
tKEP9KcSbvVzGh7ouWkyVNQJaRu5ys15yojtm/OqtuscNmFz+0T2DzuJQXSQ4v44ydH75wdal1lW
66JE46c21liOIf9XNEWxcUD9bYLlK+O9Ns/ISTBF4CwZI+/dC5Z0RZSqXcjq8E/SLE+GthYGCjKS
YeBNbkfZxadRgBM+IAy9KiVEOTP0A3/91m+Ro9a/sFsM566xpk72aWU+nl+mghZ90uUZIQPwW8/M
onUL4vic6ZcLZmL0z2Hqiz9xBL14xHfWQSQuXJJYjoWzOt6+MicdgFgJZHoe2EQAK9Yx97KNVdSt
5tfgCBnXrSHoJEpaoVr2OBAGVz63a2cVqLMNHxJpYVaL6gQwIlqbffOXaO/aIO+96c+QSAN/VXsh
MiDdNQM+HpW2SFuCiSb17or8mtdQLVYbRBfKyZt4ACXGIGj8B8E2mIDiAr9zC2V7vo4wlF7UGE+L
fyllmnmJe2kE20Vzh2UJT6Ck+Wl5RtOWtN4BiVyjXFb+gCuFdPdhZFLTgHMHqhsHBkAdF6x1U33H
o0BvoIxJ/7EVAXHSqA/TwTxqvMJtFC6/Q4nD3ARFLMH/6kHIZiUt7PiR3w9XDhKn7enNr9hGR2+x
tHeWRFPPPbRAlOerVW+NY7dYoM3aLQ4RUdPb+eGrQkVN8lgHrUpoJdto9/PRCaF/vRxerH9zODAr
DYUcaOb7JXarRubZ3FIzdZ04b3XbLXQBe+qRTCacYVZH920s6EAanVTNObcxH0h17t4T3mqN/iGa
LRYYqarAaZb4cna9Taouy+i5V7r+o/R7O/5nuOxLVyV8DVmew+aucrjCwYjW6vbiGRjz00nrr/qP
fZsGNsm7EZoQwgFiN4ooDsL/uE6xOYnhydFlfab9hRCVk9REn9E2WXiaOy5xkeRZ7v6Zx7s9oKvw
rb3QnTzSuUaTMz9lgiSVMxh0yJKYIDUfa10x+StV3Qp8o7L6osNu8tYdtu1EPZ5GCAUXy1wSZuUS
ks6o/Yxr+e2TV5lhCeDZ8m5W2LrLGjaZ1+bT69SsaEKUwXchPV73/Kc4l0axKg0ymx2DKUnX6+ry
YnHG8/HWhB3WnPE26SvDw56SjQhLrcJ9MKZtZKcC3G3D96vd8WITJUEeYvvpMV5yaAfn+DcGD65M
cKzGID4NozFE7crTjV3shGdoGd4mUB2TQggDXk4qaYKu/z2XJa+BKa45O9b7Zc0tqgNYCKgzI9iu
PWwXjM94EGynkvXeqU3PXgJEiJ7KcmbBuY6dVsPTToI+k2wD7i+Ox9QrG84F148vi7Afpm7TcEzx
jj3U91Yixqu5ad58keF+Jk/lS67HvuZlXQTxKc4TuFgxofBCfHKCzupx/Cr+OTJ9jQrdpB/hBJ7H
6ARgVbsq7Cuf4ifl3DIav/QrBeJlYjsjLg2J5vg0D9SzFBjC7p5U7yMOEiH6sX2TNxlVykA94ER7
uykLoOnXfA+pZsRboAxQAHElGrmwW56tmG/gE8gcpBp/QkZq0nldxBy1tUrRwliWw+Y5HykufFKQ
O3h9l6CmK8jxUO77lK/0dmyAVAwqTLwoqzNdMb914CosJQEZrFnFwhQsuLiElH3i94LQU9yMy5YO
u39oLplQ5hXX6PAW6GDZA+RwCe+rqhXbEebU4SFAngDczSPqUSW4KxBRro2bTfT07AQkdpO902PW
R6DYHD7VFLu3vAbP0jVa6tA2iC/fRY3qSTPUXKfsHcdjqqDOo3ISbQLF/4j27sKaXsvC7M81kbUd
KCKsxc2gPnMeX7+CfHSlU21NzCsn1M1TZ3sc2VoHdgW54MExfs/zLwe8YQw0odsdn3gWZ3lLRsHz
jmBWgr9C1sW2po4veVFHnnjMPdV1Q7kBjF353CiGwqzVZ3jizpvBrr0RcVlE+MBYOIwdf6t8eAMI
dJHTCA3URCspd9X3peqK6/Y3iww0+OtYP8AkQqE91hVHjXrE5MpnVs6s3vaKUqW+v9i0Xja4Yr6X
KBfs6W/V54zcUSxKNuCcaRBxziPd3H/EwjVBgPxyb3ywKuaY4LIe+XXHyfFsbzg2eNFGGVjzWIat
J6fMTM4jJFBmF2gMTW65dI8u9tFmQEYU4kUMnbaFwhcqK2XphvT/JtIT/D7Z1akIzw3ODd6QNwV6
oWxdpAI00QRCnGogxmdrmoz7Ja2AqW5VohlMLLHXB9w9/D1uM5r1IieFbpzCGHVDUgg5vygk+W4J
AX44Lv4F/JqE//AFROdbaZurr0S2+J4/BD2ZK94dnxvx7TxjRLQ2G7rM/9+ZZsCf4jniflCxRjiJ
k4boKRfu+Nb4oUQMGm7WHQJtuyo55Gfzc5NuLKp9nUx5Yvk379w3ajk9FtqPR/SSZKS52t086ZOa
YFytFQtbDGRBHY2GQ0KGhkuihoi7k/DOmpn0YEc9KtLR/QFnRHHDroOlztxKB4jST2MCX0KE81RM
rI+INaPtjJtRk0AgmD1sPUaVqNP+afzg0gepgZHa7F3I58iUBEt9gzW+3wu6+ca9LgOv3nJ1RuqZ
99YrK+GncEufNGaFz55OYgUtlnl3vnVJKxjS0SAGtNJjMh5jh0h6GXys9ydNWAUR0goP/RGetHHo
IkA8tDxCf5PbL65Nug/U8nSiP0Di0UvwHdKa253TVTmN4G0+qfD5yDry3+iUt7JKGbOHEfKayayX
ALZ/wWABk4tWLA2on9u0hE0yAVW6LnQ+x62rmKzSReXGs+46iGhL9TwBTZ1HF/ilkKlV/k6UuUbN
cnH9/oI7RW1k268VfemE9n1eRYf1vQxd9FQ0Kkp2hckNGUr2R9xhrNLPSTfMJMFl43I+VFX/eq8M
6E0KIC+tuUo+GjeUcrdFBV7VsShZDibW3KCFj3E7HsAVJDhrLc8o0bS/pPc95moV51ViR7ThsAED
c86jatAbBi5Hhaa9KYQ7BEjzsLENfe7len65qnS7LvT57Oo2loBAJMSHO+Th+UTCM7Ixh11+0iVc
1v/+mSxPHW16Un/lSKdIzG0zhFkGSCsBaEbDLhHHHMbzaBwo4SLygFTPX0HSJhZ4TBsq8NmYQlCT
bB0rBJSF4agK5edi8tasWdvTehctleYaQxyKhIS5CfEOI/Z9ToOJrj+R1o3HEi/YxtNy
`protect end_protected

