

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HkvkoCL0GWrNz7UZveLW08/L6sfDm0zZGNFYNcAn/nN//DPdCiitkWZaJWtNOusOSxOuhl+sv0z+
p1lz7dl//g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
krz6nWvdzbpcwbTOZlkbRdRmwRVOtCA4XeulIVQdqRCh46kKaQ1Az7t++QIQaaeY+GuPXRG5f+RT
/lT23OvjNTfUf7qRgYm7gawbEeSl7iLfiLygAHoLsmNj+AH8gs8Hs0aW+rBlNMkW1CiYm18CYdKe
BMk1gzJz99beaH3xgaI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S0rVRcgWQWVr47wX9qwnY6bNCk5yWX3QNuIUM8LuaX8hn/SFQmfJmPcNes8Folei/+/6+LEFm6Vx
Qdmf/pAXoMlDqA6Tk9J6e0EI5j98K8SO2xXJ+gzU3YFj+q4fP4roFCd0CsvGnNVnvR9QSY67D4GT
hyqra7o7wYbpUx2mTiv2gaLMwnoWnT5ZzsGdEf59HajWnwkeRTiguJpFlA2id/NPwWgZgHvKZ76o
YSHOqyB8zjfPqIPDhrl7blVRoBZvXmfF2bfsq19DFJHfG7UvY7EZPYFBD6y+qNjbBLb+5dGFTo4R
zppTZwWHLFQj7AvvDn7yqC0n1LpKK7npCeJwig==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FWYznElFJatYtjlAAT1QGN7C2Fn0bGHYIFjGBmEoLmnBxd4gbSui3fgk6xjK9rjjplTgHc9C9c6z
TaKY9/4GWl/7UJ0kugef7sQQoHIeQF6ee7w50lZjl/t7MzkZrTP5lkQthyugzPF6QCmhskF1nRLh
8U809RlH8O1td9E+1vzWR95+g13/K5/hcQtfJV6eMA0T69sJUMfVXf9ZGpdTEe+8VgstiL0bspGh
nonmspk+8f3Lj48HEmy9cJWNiF23grWiYEzGAr2f3JfUuscQoAvyNZKmszKrqZ+SsW18FBFVcMMR
aHTvY8YDuc/AQzYbOqTYkc0p9ROnWPSlq9UfKQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
l2MUNe3fletgp7klnltItrRM3tzG4+89OKOcJcVRFyluXO3yMDNdtTkvc/SDua4RluI8ntOM03dS
viHFsuwjhwYJedBAb33tsrvwg7rG9tbt/LEG/pDQgEQsMWzKwbaNYxt96yL1pqBTCXrawJRgzhDf
3V9E64J00EAhc+Oi7ns=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OwI84vg3qgYuEbxZTTdCAx7VKjyk9xG5pPpZRLX9rHBXg1TaS1COb9wYAyuUkiMaNfwU+43FnUYR
zPr+xswATVVwp9fQM0Trz2CcY0oNj9FQu4CbQMbwQTnIOsyvnJwIujdxNq8gsEGemveYYjxPfj8o
WumIWJs8TCPZgcTg7V/Igr2IkCv5OUXoa1wEoiQnNS8hgrskPdguRrE0QQRg0ky2cZtAABfuiBng
oKj2VdTugfxBQIi1J4RVAb74Pk9k9CVJDv80IQ0VWrPTk5H0XM/u7z1dp2SYZUzGAyorho9pm3D+
vSFM5cFHGC5DCvaNPak36o3DJ+oTWzbx/S2Y9g==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1lsEBCKB2sqDzwDdv+Ksc4XOO4/Mx6iEV4rMgINzaVZhDq0geGva7klDVIzj0wbmLz8Oy6aAf2gm
jnjEr0kr4HwkpIFY6bw4gHSiuL42715ss8LC/IamaJMz1UyvyuflZZ5+w3WnVQUVJyFbnT6PcbiJ
iJr3kzP3kvqWO8h1atovR6OTQ2AeF0M57F5iLaipkXR/+ybFxvyZ9/Mn/qb/hckXmTrKdKyWjYzq
82ZZ7bsguLRLWbUGJAR1Xf2ACffKjcMtafkrD7fm3SKeBuj4CCaR/XIqBQ/Vqh0CD2XwAVxA4CgU
ZEl5yQsW3u3xjQa/H8EYOKX4ui7vrtobcsVM+Q==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_11", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JbNe8kbb6DVzM+tMySGJicqHJ/6WO4jSB3NMMp+SwRzyNOEwlfByQCraQ3Y3nQHUREYyNsKKEufK
sUjuV46dEokHCsNIUkveT8nCh+SboPES01C1eQx0/AR8CKBy6y/sWYwi+cSgLOC//wf4MVo0NRlr
eZ0/T4NrY4XEQRt4OBnbRuWmVqhfEtKNwQR7xNIqFBEeEC2O+ol58Gdq0+YRgeRtdKiHyAVVSxa0
bMzI/T9jTTCNMKv0ckDJ1cbw9LGyoLwKGWSWrxLIFXUBt+xE59mdFcCOcJdPGespM1nKJzWzlXnO
JERLLXL5nt7hTwByS9AR0qDsi72yUzO0FxCuRg==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nIxk7DmB875soFV2AQWrZMt/6MixO4JJ3i54+8Qs3fBsH6g4tDNCPbpBqLlDed6dueueFUP0dHHM
RB9QdEjaoRsDWcLMgii2yco/P0MgRA4zsSUGcovzMhypbrSuZvmaTEzWy52XWlXwmKs7YM96nPq/
+TMw/n+G5Le6vtVfxveHYs+NHPeqVuCWg70NBSzkoShfjtC742vBlPPhAT4TNTPpDbQjcMK5+KMb
7KckSUrXtTbN2R3+5LJhQ0B7eVbv4QRxFhX3jgi+lsX0cRB3GokzHZJA8SZkAZj38gyTfEqTEmuh
NTect/sqzLJU6IZH233HF6Qn0DElnGjCYm/NQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
AhraUkthYzkpa8qcx/8zKGRxCEr+sehZfAZXAIU18LJlDG5ps/MkIN9BgW8OK/CpBfXUccM+f3U9
U+CSngm0wUg0MkOYWAKqKuFTIXpDxKtVNNlEsS6TidXUOgG7AAnyiASFbAJXhwcntBIIqwR1pA8i
loMRd1xfkTrCyW8+8G2qw8mE9H8ykXIveShR/9PRp8YSBev9A0M5oB5x7SbxIBsjQm/PtNIdhzvV
LIoane5NWHoE9Zo9VSCFZVaTTbzlQfvfKMyk8D6q6FmzJoK7v6WLdOfJN7byIKMytWHgJGQhgMAX
pyLpkpwFTKWcS+ODH17/r6Lr3qkV7mCOsdi1DP+6S0wjOjKh3p0i6/0yxP3M15zVjNUWCwVRTzcZ
DeF74RCLGxwb9+WAwv1dtQW6h8lzdke/5xUX124+M0JP2rDSLCZPUjNhDUyh3P0aCYKYh0h3A8Mz
wfCeZDxC70WiyhNf50uXX6a6/t+aW7eALJMzcK4T7d2N38/1ivw2Z6cXieT/75Hr0d4B6mIxeDLW
D2mpD1Sh9VsP/rG0yrer7kLc8Vq5mUCjvqiZS1QD/wigzd6/jpfJGwtKTpL4CwIMT+B4KVdTjeJe
jDA6UULsi1UhNNSCpP0rPs2h0RSAn0xQOORW0Roq+5Gc7zj58CrbBSderEVzb9BZNSXUTCT5SydT
2WCTpBOYRC95f/ZpiEmhhXW1Akxtuc/YN4Q3cC4Z7eRqmrbE+Sxk8KxHTIt6uiMzv40Aa58CA4Ct
k+u6t15BbFf1zzE9EPlyKW2I1uhZmHLVUZ11b69863+D+xBAh63Kl+81xKn3N2RbPSLQz8FNAIMW
ZYkTZTiYtMLrnRLx2oxsT1g7SgsDcvo9iwmuLqHiOCNQlRu9aCXVF/+k0FaVCRORiwFdbllHJODL
O3Kk+24JhVfC3iBcA4dSA/aphpHf5aJLj2QlAMHlAezHJ9yPciPEMSeILtrPGxhmGr8B6Tmke0FJ
Ab+Qkp8PB5jId1xxCdKZJDKy196YExywpTvIubKhzMjgLAQvu6xNXYS5/UqKZ6h6dBgUgdhHsJbj
WC/Dz8fAJoBczNVFygwAHYs9vRWMOBpHSFstFmF6CV2hipk/z2hL2JnQD/1T0y803k3yTE5ltfaz
9JdgmouaZM+vIRNDuvtq0JY4vr51mTHL2DVoN5Aaysj8RMDWPxPNvE8xkIMRBzKilHinViWwFjGs
FindHSfOEb6tlvdScByfD6Fxo0Fds+tBpjW3s5nK/g2jr2bA51lEyCzdIGHp5OAUUBsQGxiHxP0Q
TSE+Efw9IHonxGS294qxxTVypotiSOCa4aRUNh83XwkippKbkm+tDZ5BVpBl8X7u/GTSgbQ7tnxb
5Y9JDwt1QTdMRmMV1tlgWtP90ZBGkW4RAa1vOcMzdIjRqz+3TIuMqD6dPDyoHF7WkpySanDLAE1X
u/fEEktP66zz5hlmWzyX8E+NnAp8eaMxahAbMg0v5HUq1SeknVP1/Ny1BL1wxLshSBa2YtEiZFuT
NdZRwStrWJMvhp/dF9KKoWw/YP2DZcdhQznHfDsZ3C5sHp4sD6CWJPN/wrD2Cv7uXIH3ZdgHohWi
u9fQch/IKjAyx1nmPD05w4R230NRrlALN96U+HsdzEQZORXy7D6HMA/I4Oe+Le8YhVM8HK/9WTne
hS5lo/sXxlYqeAvVh4vKjnZA6HDlyAORre6dHnfotW/0Q5ZVy2GQ9wXdu00UQmHzlB+NxsX5NCax
Xjv3tfqWxZctHo/M10UwDMkPPXtH2IRQSUj2bbl8A2916auhqsV5sIFivcOXxR+r68ABMXja1POG
X/bl+7LIjG7z9KY0cb98MRpzAs0PE05dkIf9GFYUvZn8e2XrRunQdPXqqDnRQ+UAAMA5zWAgdVGf
PtFfUNFJOyxBWq5f+wMt2CLuAz7XOnM2XumMEBcdujDWJb97ODRJSdW2xZHDFpTm+p2w8xFohZ/e
xZbczO+JuAyq316iVwKcoe3yOmK4gsspk0H7Ta/706tszqtUygnwty229ubiW9vWyYi8wIQoQno4
AwzyUZs16GmTfjOE+Hm8nX2F1zPNBGFriVF+FzhCoPZjScFMGXD/mQbMDfz/jj+RRsuFktsigJc/
DEgT8XTmX9BBqFqKTN5QyFU6FQQVeZ6NcjGO+mJp0tDjQMQihkIMQWJ1Vn/DmMgqwYF0NF0GZQSB
FvdvCLyAvWpVWtaxaVJ+lsYdLfrWu43tZ7ABq27ULp0giYm6jk9Z7x7u2/MmbYjsFg0rasJfjJ23
HJyx6PCtBf5UmoBbKW2L83JAQe+bfXIxl+XEqrTtuHPWruQlgH+LRD3TBmUZGyZ9ouJdgnLeLmmn
9AfWgULAmSdhDacFUIMZ2zeNX/Ww57QfOe9uVxySD83ROqkOIIpRjIfdKLxFkqF7PFDBlHyvfCkf
eVcUWxcAVj/KKqHj9pVLlmoTeBw+ay21zcdTlIZmLBnb1U+3ItiUyxSOuWxbWIabnIbfNQrfXjuP
NnmLhbxmPN3WUsQJb6x3SE+EJf7b3Jsc9QVlLLPQInQrXQLCiWI4UJ+DF/NLfKTXVf1w/F1tztZ/
b1FfeGnBVpk8v62wM8L9Ot0evgJAjeUQuvFnLXIZfrXxhrjvJY+TmQpffKBYHrS4fkAWB4e78QGr
zQ2LT/H8HTcrM347O2O8Uenw+eZE6Tha1yOduMnVMIbxdZLLQhNI4V+Dj2y46ydVMlZ6V4nVJj3b
3bOMvh2r0lAgmznDpclY3026A94wEWDx81t7PQCBxM1nXuTCAhxOoLw9QgdV98+OHTAFER7i+9Cw
QDWEo2JhsH8H0z8/KhCPlBP35h/v1u4yXrwdFcURPShtn2eHmjQh6gHIDS6ASv2ayV0wdfwlsv+q
7oTvsvAt6P8WWOXoy+fm9ffo6/tP6qwn2WidYcT00awx3Yde7IMALQMqQfXaauLpiu3yh3CaHLox
ddehnIq6HvOCxbR5X3cH6R82dsDK5poGE/qVK26sFkAiMdNhXkcGSVksG4FsIZRYx3F2OxbCwRr1
g67662Fv3+qFEPDBLpY2v+R6Il1sl5Cd8ouQ+KK/gXC2/HEFCAP6UPK8SHm0D+mOUM4r7QFJUrLL
XOGRttKWybIeRKbJCaDnW+epZpwAh4oBn7a8v34u3oMc7Gmpt6LL0MVNZaLL7dLgH6JRGoAbaFQg
JtNRASt8iHEphQdY4uBfwy4PUazwWsiIDz8pcoIZOHwEi3Yd9DaJ/aqSlluFewTInCzGXQQFSCkL
KhjJe4lr1ZNvrBiIzsH04wXb7tZnSr+V7itXrVACIZ/9P+i6TKWMJESxfLlGiiL8UEuOId2udbTM
R9XvZj0j40Z6mwbImlrgc+pm2u0Uuof2uK2tIIGecpJEB9lk4+IvIk855qflBWD8vH9sr7p50jUt
c3/LFulteaH8OvPCTlqc9v8BC/338Akpc1CSs5vovxB3kCoCi329Pjipv7SvNsx8DZy0+ah6GWh5
rTMz4/JJvYt9m990VoGykv8fXIGaCokq05Rl957dEmMVRb10RDw8kaI1M/g+NHCFofke8nuSottJ
IAz8jsEMmY98Q6hhy/AM8qkIPDXmx5ID/qx3vuIW4qD3CO/hK53+d4HJvUUGaS8+4US61/0DQvnC
EAEmP1wOVIvRHEv7xFYbqi1vHRVCpiVhKtxCSneOj9EL2i3/YduP7hEhwjPQnTLTmNVyM/h2MbFE
DCgRJO1l7ps8I4An9VRtN3w7V8FvFxxwJEgESZHAnLObqv11kFJHV2RF8WPKrbJmp2xV6QbHXDHE
Rv4YQxkzs1vWj18RYI2xCM+ge2ljbXsNn1OQNoqep6gLOI1HFHn9abXScR15jsPk/lzjepwNpMPS
EkuxYjkAwIEy2eJwmBp52HVhpX6zHglOYrUDj/MqT+PSn9vjIEgzHg2K1as72LHkQyg+XQUtuI75
qOh4fsbWMIkKTXAkh0BmnokZd1vOoYkuzG24t5VmuVv1mw/l0h/6F1J8gXQRAdOkkmy0Ossojnxu
md3pPf3qdSbcPsgCvRYVn4e2q/HxPIFbt3iPzjplyZ6OfS3hPBFTiS96L9cbnX2Nw6xQD5eQC+Wv
FstXXZlhAnJqGhFsX4o6sWWBzbIMePcbgR483TtPdyNLDk1/tkBOsRmFaz9v/yXRIiXdt9EqxIy7
oaaOWzcAqfCIVMC/DryH8fXGPtFslXk0tgbgrLGb9AFvE99FIT03cv13uDrPO74tITBPzs1za2ga
nQ8bQPmXBUM8JrcNJC+g2nA2XRtBmrZivC5y3oZKdsvCrn4Kf2VvtKmSTH6WGfWl5vog1FnsZkzp
L+RnywrqweKHZpPq57Sl7L40kyH046IgVAANzloBq5qxxB8VqyIrZ55bBh1iIDXgxphAhIJ9bvaD
XKcxx55c3jcy/H2PjKceKsm9O7URoItkU9clSbHzzx/LmeUBsPylKO3mClMYTg0cjm8BlaeNhLTN
aVElEPC04bnBMrU8V+Ytc/Z9lr1ImHUg7zuufLoh2I8tp8e+0H0M0R7BxExzfWU9YijCGD7A6ukA
lIiMhrOvzuTV/bBbq7Td5V4JpBEe/F3zTXN4qrivXNxNP5i9P4LctvhAQGQCNmRNquPjVVqpz1NE
wB4ju3L2fsOsL0TTTLC19lg6mqj1YVVN9QaySdN6fwFm/AVpvGKiISIKV/dLahXwuBBaUBkBSiQo
qEhvkIMKRvH0aui4sCdLq/dnHDqSjIAVYFNV/yvIsY0w/dB14qALXR01E/tOFFcq/tNcDRvORUl+
93eCrwcMQ/s6SjfdDvz0SeqaMvZ5ythOWq6Hx/OYozHGIxra1geFS8j/4x9oSJjd+mU1v6BIQwdQ
nImIv7F1pD/xgO6p6k9YpKIkgQVxDl7kIG9Spmx3U1GGrmm0+auVUO+yx25HJ0lRH8vSQqTbyuKS
viwsvlj/4rawwFJp7SBi23+4bkVIJzSTjSmW547LNQVoG+CV/t2JUH1GzqGudalEP60CMmlm2vtL
BVzt/hywQNuAtnJAl0pdByxzVsFdhy9QA2PKACAzkPNXsCZQkmzOFIHvVcBOPks9PNVvvZV6U8cC
ApdMWGAu+WNcyvZDoDcms6IK41jmO340B45jtegTmXR5FH6mS7IzbTA0i4tEX0V+yKqfZA0VG2TR
/U823M1ZjWqns/Mjvk4DSFJzRwQJZ4XfSOjRgeay0fJBj9lARoV60NWceK4UVSyrWKgU/W+PZsh/
sVhRp4+lsSVZcPXaXeHrktdJ7X/p1hnPxR7EhiJMnHDLOUVOOvGJflk5F2b/ucjvlMiZE7G7i78V
PU1f0AaaOxCVMnFeGSiyvHhBjq7gYpGLlZBo5GXE0adwmrrL7e5G352fQo3J8rKJBFMD6UMSJltR
CWs+MaZZSnA21PMqQAUoHLnLkYw4xvCJH8PZFFqYMW28BsKPKOEJImm4hfQ0+vFrthwb3CIstjpJ
oAvhrHcCtTDRk0Suf3eCrsrkt3KB9l2UasUJ1Ei14SQreZvQdhd4OlJe6O+zvs+lop6dcbmZKhI5
5vUEinJ1xM+R7z6OfRV06C2Zuds2v8WvwWWzViR4/lBED2uPWBwVRVU8J2WUOdBWyg6jU4z8Y6KK
brVKC3z6HD5yk/oSX26jWosxh4OtIqxfFJDN+JzJHKnrelhG2f7IrN7n3eegOOE01fAaVNmncLlN
+15ewLuNTCQecFDXi6p4iRqKqElORJpoXAHCg9Y8E8/ljXqUuuK9iaQPm9OUzHp6jDlkWuoMKVw1
9G+NRQFTLO4V5pjW34+0BYMYSDXa8zLY7cnTFHu+A8CUEg0bzGMx7rYK7hpym6CIiTQzkzrvAcuR
KnmrOaMvzWCD/7Kjq9xPagrFpxMNYRqQwzu2USZ5+j6OLhcDsmRdhCTL7JDtRSIoVpBIPMYaPcQp
KxPRp55baNqL2r09qXrfU/D5Uh5ZcpGDt+twegGApMtdo10Z9sZbjwoLwFRNvMTF9ZXaHZ96uaYd
f3t/PpcMiwNeCKw35fXDXyubaimuMI5YuExCAuio/YG+pURTAM9eva/k4nBYWWReuPmSC54LzH0i
adoGKqMfKs092lFkvNB9DlNrkj4N9V14lgyku4FIZuE6ESSQHQisVgv9DWyIsHZLK8g6xrh8hszx
TaD9sb0G9fIitLgHS0k97MHFQO4q/Inqpu9F6MyjaMgnx+CNA2Pk338SQngvPDO7GMW6ZD8SZzE1
agMJ6/f6KwWfJNMKFujsrBn9fkn/yLMVwE9/1lvWTeNLdGr+w7rsg3rD8NXQlXJiCw0Eq0ti5h4o
VGSqYdHZHvE5x5j9cshOW59m9hX9V5EMVzl54OvNIXQlC8JebNZckgLTGrfjqUwi1YdGruO9/qWw
DjnRPYgB97V5ZPpMBNdvmcIUGo+Hfi9x/7ZSHMUiog1kwyXKvdt6EZfM73/idJCNlcxsveX9uxOw
KGHiAJBHiIKIDpdr55B5/j9ctCQz68YBxaVoUI/E2SCY9GCcew/Lg2of02P2k5gJTuABecAHhzG/
7BBJAUgLM5ONp5EqI69QQ+hJLnIZfWBbi6SzA4AcS+gO2D9hL8p+3dWhcIs6cdE13X0wv5Cms5NS
N1QBsT/me9jNBrucs5Txs2ImsfxVYQ8A+JK1gRMq9yLjI5z/E+Xmt8k9Dm0wvXbu25XqwGg2VyK1
eMadvQWTBH04l3Tk0l5eE90nMQK2TMtcNk1SC+djPEAsXesUgS7sd/+lV8gBDwAttaHGyzaO8QWz
Ju8jS4LZ3RSb648Hry8XDxoVmEhCaGADTtBpgN9RlUVHdwIjUIm1Wrcv6TDY2w8kyEB0KyetwQK1
xFnFlklwNvtWP76g+EeEO0t6A+mESJYrUNyxQoLuNwEUiDnpz3FZ7B5pdS1b8ubsTH9Xyz5UDE+y
x9gbDuhqwB4u4rd/vYopsd1549unqOAxL4oXFz0CGEcynCnUb/oLE3RjbMuaFYduumzBhliBqnC7
lyD/ZVl8NiKXHLuw1aSg1vCT2vPq7q9Aa7P8hRtGtFLINTNAR06/YZ7xVYCYOshJkYnX96cwPNXl
AX3N45rVfd61bA/Ny5R5TyuHG5w803ngJY8Lit9AuzQHockQRGY+Y8mGlUAW2CkKvJbkosBJg7tH
+n598AccHTtgkWMueRt0fOCcnE9/P0z1mY2LDb1YNFNkwoUcz8E36y8kvECEdEqFXgDL4FgwDB87
cniajc1S7Kv5GtFLKQfOP3EENMFXwQPQbQgqdySSKIgw6c73IxmsEQakkRrRs6zRYBBWeLC7LjRQ
wLfp6C8gfwiZfGOaqY515xZROBPwHmuNU1jXnOpMTI037fkUwbEsqA+NOE2ePdKx1Rl0rPE6sW5W
lDqIlPkfBz6FT/aVqV5FMuXTpxkCPnWMJkVg2B4KibcnDft0Nbe3ua7cdgCqv/Zr7XaNr7VWteFA
93xJ4zSm7D8R8AfXAfRMopwfBHD4gpfUIa/vhAMM4u7UYMRIdFLHxzkR+KEUZQSDKMYOiRPspq22
sTeTsc9wOsjjq96sadhHHV/ME95W88SbsVWsXaoYd6aVp8a10AVEaEpTIFI9u3mkd2BrmRfSQmjF
tRXwDscsQNjmAs+Cnl3+gEmnaQ4Fhr0koztcd+SKI5Npt7enI5KXE/0azkEz9hMbWIPaFBwQTkAo
5e5eelq5bv/+I4WGf37k0am3KhJt4rXnPiMM2q6W69m+nEh5IlRnqw9IkkNkIT/e/+EPrHQg2Ziu
4AY4+MuvMBotBASeGMqzto259y392u7fzO8GPHrLhGRiK4CEr+JMcTl50RB55crcxfotLDOPamSf
KlYzTWvMwrxUe5dWJlhwhdXRzOUr3vjc3wOZJiU7tFhv2xS3B2ckSbtObZMBM5QKed+C18sso7Jd
ZkDklwQNN0J7OEW6VIfRUq0BTnueBo20y8qa8KjZAiSqbNPpCyvY/AUm2/GTin4MNv7W6xZ/kbVv
zkxhbR0GvqGpm8JmCYQhOxq5EYUncNIli1u63+j1g6PqPxYtih2bO/x2u5NCT/2djxBnIefhsIkX
yRX9vMAuTWZU7QHropK4+dFyoKKGMlMt1RBXmhpBcawUVmT4Kfu/WMgLVvopSDniEJ8GiYyKE8rN
wWjGRmRi0CMp8iP/SEuVn4wPU7LxEGL6kKpFFQfEm6XCGVaQNABfgkSG5Hw+h7FPD6mJ6aumE73s
fMac83CX/3++p1wt5D4QcZgmF6H5Hezyup6ULyaFCckW7ribCO00RIgmnkLBOr6FZUn4D0HXbAn+
ELWCIboSZEVfXod/IUJiEn37ITyuH6HJLtwVWtXTVnGQ8FYqYtorW27MBCZPkGGnyfUi6d9De1Ld
HK1w//MX6JTNxq9Xe0rtStcE/lgwLxXk+424DdGJ5RL9KgEJ4q20i5ieCdZVHFjlVNn1JC2KxABj
YrS1M7UOteIgtlLkI5rHD5V94Ha55Itu8NhayAQJEavIk8JofymDXKItZCiXfkvU5t0ZhZ0TSaOP
2pBQmdUShdGIzxXRGtWfEArG5yiGHhQubyepTrozi0msfL6+04QLJrFZAe9U3u7/kyMgPjUqtPeZ
qN5iBK9V61R0p292PbAyckpq/z+NZi5l9IZoqXdvQ2QgV0CD6y4CXifcNdH+/D9TzW9vaeP2833l
qS0K+hu21mM+z0M4w0o06T+FvmubzIgNM7T7y9r3NXB3C9nmLBOEEy2dPAXtopBGhJca7bAz3a//
F66V87gfVI0vfOsn2eZfYVCYEDml8JqziaA4CtDzO0yWS6ideNN5AegomS0nqHpugnHXfEqBr3CX
lvRpVRfOssjR/f1fu81rBRBrDsbwzTOUEqdkJrsrXnSqptkGz0PzkToQYqKkRzsu18S6Szuf1g0V
ffAoLeqT5cNMLQ4ET1t/9YJl4PZUHlLMQ1cM6ozijLXL8fofVkTwjwGUU42zKaTeudT5c011zPLP
ySsyAaFSI/zKq6oMPrFMmlqVyHotIdhCHzN4d/gNaRLMTMT/mneQ67L6AC9xsjkaMYcRZE2jal7p
ajbXWMqs88FbpFn2zPCjYl/6YI/hyyUxJCu2KHY5ZX50GbD2LMAhoSx4kII4S5yQZKJNYaFTuOTx
aNNuczAMMT33JeHNmAaJS6km7JhF8vHkcFkJsBJ6/3IfuBJOEE2r3nRALEgacbiYoPUQyhfe0IND
fGeLeGVJJlv5O6ZpGeGTZs/iylj2JE03GzLVaapQ9v5dzXsDrCkTbm21jvQdC8Gbr2t6b9EMjm6B
No4ns+FCylRbbm/mOVNtLy1QiRL41yfQx7dkHE6w34kGZq2r/S3IBAkWLGw+vxZ9Xh2QRLc65k4D
FOHyRv7rYTyajvTVNyg6Y+CmqrshGi2Ld1rP7hWCNPi1GawzneDEhP1954riRQ7D2uo5Ci+HKAXw
dDnudZ9lops2zj1OkQmv6sRjWXSWXajw2qVOr9DXyF5zKnMwi5VrUbibK+rzUPQOXnX1eok69U0m
39eBm8TQqmwGY9Cxf6Iz5E+Fb118c4yWaOoXLs+CrCzOVlxZpw5pQ2PQqvgYwQkUuqwvjBsfemX4
sZd9Ma4Z9uvAXZ9AXSkB8Zk4mmzyvjfQLmrARlmk8fC0IjYtC7SU/qrhuIGhOwRCqBHiO4eg6UK5
njcTokblgh5PJfoijbzfPUdrFfaSuH9tX/aCFnQpv+49T4Rdr2VRMdG4Wic0wrkjBoWW4AH4jq1W
u/U5FlP1psC3lYDuF18UOfACb8KQ5WoNjWyAjLsWEVriFkah/kFBhMsPegmb5Dfzg8lmcr+ZZKah
HS9zR40Kkar07yAJyu0jBVgvF7uVfm+4qC4gs6/6ikeyoq2uNlJH6LHkeadPu8sqnZ7XvQ6fxJh5
DJo1VSYk1vpXzAkwdKhV2qHN7KM/XzpkA39YanxcVjoGI7TGMF7tS8s15c3VobQNlzrtuG0s8G3B
803L67OKEoZ9Vf907fWK641nUGzZbtbWcidGHSoGM9e6JpY7RrhlyGBOKObOFMdVvYifN1MjXfeW
+8+efBcn1/O+h7zL5L6/Y4NRXBQUVIScJqKC/KpLw+nI1pvWkbgoPNySaOQunpjRfJRrUy2qbebz
of6L0BEEtO0KjBsRaa2uLIh4k1bQ3ENGjZpupNM+Zo5NvnY7vVXI3ihhPZ//Jv6+XY+LQ+Y3q+Bm
MtrCBi6hIjBSDxBZifBcWtpNh8RN+dTZJd0lNRfEnQSuQve7RnhN6kfdZG0jWz+scr2jy1Vjl6tF
ITKuTcfqif3X3O1k+dGQzgP1FBLcodR/PlHluH/JfhxQbjnG2MwozVsH0O3HGVZTYue6XVTl1oTR
Z/Cxt+SNeZGa+JbUQqZq4Y8UKEcPEqmqPDWp8V3PP2qIpTEZ1OdYlwY5Ik8xtPatLBQIDJu1/Afg
e9/XeL7Pk0eSMZi79pCVsre9EayZwOr34hg+5Sf14KQnI+3Eq/uCPS/5cI1B8HwCErwpzxtoIfRw
H1tLEIKU2X5rMK+NJnajxHPLLsxYiZS/lxuOEB9A0vS0Flp/i3Iq8S8Wi/Pifi7k9coeCUgiVZTd
oIrGDE/MSHYv0SvCYHsNdmHNfl86rtSM0rwBgu+hcXdkYovNr0iMa4blIoaDoUqDTPzduuAGQMTk
WLzKUvdBxvCGvazdVmkrZk3Sf7ZjW5qldxykMLdhXKG1NWzDmGAaE8xWhKmlZeEYIQxsGPPhlad2
X5ddWL1E5QEYnd35hwe388gtM+niqYq5aQzdlFUhKD8Ad1lD1L3My8E4jBe5ZALXs+0Y3wsRnXMH
56VabphTRxF4nzd7OENAX2GuSuDiIjI4uKQsxUVtK2oznw6rdxuNIc/FU3vyDA+5w5mw+ml2Avlz
O0zdF+D4EPb5vxISH/aEs+ky/X3hmpZVpki4Mvtbc9c0XxNgNpaGQW+jOh7VcjSg3Fe8GB8oDRY3
fiCAKuvRL87xiVH8pYE7Q17uReqhcw2OPxkNGz/zRiaHi4iukXoEqTAifdUrcQBOks0Kg31SrUkp
PBnUqOXYxeocLqm3aHUluhpaTWlz6Yy607MZ1I7e8CYaRXBIIrQJi7/mF4r1KukO056R1/9X0mvy
lL1hDp8hkJOC9PFxEBGF5gvKaTI2MP1Faw4iSIK9Af3FV25g7G3a/elGmup3aMpihYospOl2hEZK
WNyU3zWUBbsBiUxDzI1utICKUUeMw9d/i6EJMyW4sgzBYuERLe4BCBVhAgHL207jekG8EYMQLLHp
BuvM0jgiNlQTp0G89cdaSbqgCInEToBxxkBnjAZ2INst0ehxqYqFQZ4KWGhfwC8Sj32UE+NIZ2TY
Tknf0CwMbH3Pqm0mmqyLD4LZBcGXLQB/M0Gm2tfcyGs6Ylmij1pdpGI1A2vkLmibw8RuQpFWOWfM
tAjBhk2katUqp5gxgPGfiDRcGV4a6ThTgVgClQ4vFR0FmB6LfMcJ+3rOeDozlz9nU4xrh08xasVI
UA3NFc5KJ4V6qDLmJdXCHq3K/n/lfaE2895qQ9OdEtr7lssoh+p70HfmVIT1E92QZu8vvcQsm1pI
t1z6rz3LzJnm22esa+RJIc4UMBzV3PTPQQvostvoXI8qgeqS40tlWEKa4hPKGHo4fZiwv8nDn3IU
ddyPPITXHlzdhHMR1azO+J+k8PPWLAD4uh3/wr9WRt52KXTOSgD/+iegu7soCTowgrItbUW2PqgA
vNtiXHc8LOqmnFPpJUzJn30xuYSnnKNRLxDS8hQMSmbtRr8WhpY0P+OWnO05zoUgML0ocaKGHliK
LOtIm4vUXZuHt6ZrTVzNZ5YwZD5PyuKQoI+Wzwmx699O06PYMjhL1bxlbSB1/mxFLnmEyimYyMdj
4pTF8F0S8D41/M/JEWN2fu4UyLRn29F1zoRmSkgsxI1felXPMxDM9a17OW9WPgUj/X2JGNFWvahV
jQf9HLxTEkLvVH8uDkmJ53ieWAB6S+rqcMYH3qA8rsD74MjZabOX1iL/DUfT8wjw7NYa/vDiTM1U
+SwBEHCw7bkOeuv3gCXS4lCXyA7IHwLqXCeQuWkFGcLOxYZTLuPlJ+ONzG2+Gj74zoAQO+nkXpDJ
d1YSsSeHMlrPHyU/rjPmQFrc+1gXIcsCTA8ncVo3wldlJc5WIBqXIsgp25u3X5wLPIoTzsWr5Y//
nbhq19k/5MJ6kW/ZullybO6ZeTJeG1pXUr/WaPqKRlCOVCdZrnIiEQIIDv59qA8QP2s8Ube+UIvX
8L3r3IXka/85mLX9QcrYQS/aZCwBro5bhHyJ7Y1+aDtdLaCpMvLx3aCsA3wJE5fp6p1x6EmgQ1m/
gLdJexY8VSmmgu3ParN2elP2hp/+GpdKBYG/PhLerLkqDlwDttGnhfzrzITCJXSs3BXsKM+w9/Rn
dkgR4g2pszqxxyZZ6DTfU11vnGTufjecQgcAMn+8eiVQS1VOWouV6KdyPx/jnEJuOiERedNpfqFy
xaHFJEZWX3XqooWvQWH7HrDsc5Z2TAFPWyUDKtP19LOuKSIJUTJ+Ab4kMaY8hkN0iGvrg9jYGBqB
qUdtrapxU/EB0/emAEwC+ASM6DhgdwtJEc5LjnGIpsDRJbj79IQheBKAloijDzG4ZuKB2QELSuzK
qt1iDW0uldh8duG/00p+r01IogTI3qpxMR9wM2adMZTENFAMQE+nXB35Qmf8nAvXOvUYgY9DEql4
DGb0ckQfqt1oOybNTnB4bUcbVYlUWRzxwz5ZRuXq2GtPY974oM91mUb6LpASwyaYI0RPWxjesGOD
ZGwiiEXu6r/JhKfgtehqCdFgyQcZtNPA9GlJfOyJzZ/gsmdaQPNJQ45uvjIlQacY7bAKztPfhWPH
O4ePH7QGhfvDqdamO3BMJoSW3E+C+tU8/wehG+mR6tAE4W9uBujGrGHcJl7/msB++PNvKQ3Zg5U9
Xx9Ej4Nz1dmYIZLk7ogPcPkQDc+hCUQ4dBAlZqKUDCtuzG4YzEhNoa16IDp/HUZNeXRTpSakcu6n
fskwUwaET05DuwcAnoIt3zvc+dz8I9z/+JDDWWhln7JmreFvSZzXFY32QFHQ30OfbqXEEcrR+JcR
PRuTHTSKtdAOy83VDVIe6UrdtD/QgVkAx6ruglXaV48PErBwWNgwDVIgdxlm7OIo1OD33L5nbVFX
2+ucXy2SyZr65PEwGsz61I3E0JsdQuBnEqPxBshrE8U2m8vcA/DnSZ9KmLhxRYLExGjrNWuba4fA
0mlVTgpTCHkqKrVpPAIzc+RD86/4ApDIg/FYJv4eigmK6L37gvJDP5FqvEYeTnho6TlcNnMa+J0V
XQGyqCd9NCT+6o+b8NeUuj//zOV/2+oXfYhxl+CAwAvk1iLeXlP9nSjM8jPJrhP/EgkyykpTJArE
5F2561qY5gu3DCdcyU9vJvmGRzDhltMAhbPHKYKBzFY0tcBS2Klpc9+BkCfOKvbUWGJpBcGWVXNG
BuIFK+B3VNuvcAZ2dad1YF5N87AENH/Ht6ZyLLzDY8iWtQcHrvh/+v2VVo4KojW2BCAAdHL4kBTA
9CUuR9urCICbzr4OItw2zGltIV5pGSa9zGXsqzmyd5nXDpdWRbWpgABzfO01AsH62aCHZpJLBkId
GGw4KeSaFCYLXZk14QP4N23vnX+Zm9NdOLtqFvUGNxyBPcv4gpEHoRweg8IKGaElUeVjBFaN7d4p
Q1MqAamPQjpTw7u5W5jpe+moNlldidD8cBw4W2zRl8+Q/iNdXVKfK9YuQWsjNhif9dz/ppVISB/D
CZ/T4n98PEHflpkBmt6CnLqNZoz/r7KkU6aMRg/uzr18GA/zYT12d2MXEb585SR/LAFqKQJc6ye2
HAv3AdY6+5dktvi95or195wCp2/bC99Kqeh78k+Ny5j1ANvyim+Nb2UP6RJRPyzPq+n854TiinS6
vIXXMZbSbnHby9oP2GzRHjgyvNLdmBQs1tzVYu9nnRKja41koGAvAl8XLy2aEEOz0pC4Z0BYDUto
KHvwvbShsyCaeArN/KGu1M8qd3yOBSdU0cB8pjDvBSvU2K/sAB4aep34MF0VqdOPeQpYFRwOr+HA
BOzZj1me5IDAD86JxWh2DTTgbfvPcl7noAV9YZ9ABqElC4g2wKgCBxPYko1GxmNbTa6chbAIgG7T
0XTos/oCWuFeiYXMBv9meva2Iia3lGzEiFp/un77nQn04cD5+PZaHgrcA282jIWDEAm7a8awoA+2
IgJfqStjkIEais1Diy0hKgzEEyMvD3MQW3dXdTo/m+Rvtes9UncFfffB53IFzcwElLBPfTfdYmMx
Xl1YmMLKNXCWeqIDoCoFfUnE6LtTpR6VlpEsyTBTG0ZOXKm//BfN+Xk6GRH9KoXP+kz7T63tsvK2
zjUcp8AKt8Pxn2vV7wzk8+ZJaezFb6Oe9mf8PWd+XIoSDXsAbkJMFHyq5+nNR+GaNMrWep0XFf/w
8qy0HXepk/Wm03WbV/dbtrRYosZDokT9DZr2VfR6x99jjZgBD9OyChdhHsv3kiR/FEdq7YqloI9G
RwTghfZPwE+CeaYAVIMYpkOLWi7F8HpMVA6HFmICVM9edxatwlLQfZyIEOmspjt/7nqhmhJqYLmZ
F3cWoTG6AQ224a9j1+sHVFqkflme0MQE7XSbnP/cWkXPDMiEI/dTzjA5BR5/MkrAAucJH2xWFVdx
fnGFLVlTLnuWHy9EUVeN7XvQba/XUTLb3vX7YGVqKAg2Ib2xvpSMSNteQkEiM0F83bf6HivqIxsl
U8b8rUkEihqEDiWhfkJ/f3Ua3bfTQOCk6qP8S/wWCfsS8dKbKULYq6dOIctGRIyS2BS4dWZX51U0
6Th0JNUV1i9V9F3wRF0S0qUefOd9S/GD/UUxBF8lNMj7NViMw0dH6+IcCcjkLpdENGKTqKbH/Mbq
9btTqjhK0+5XPDd0KHNdBp4hjsaS2woW1OA+haDUYxj3wg8pr1UYxZoPY6O92LJLMVi6S6en5oZD
ys72Q0lrNX4pQkbmFX/otHNp2wtd5Qf2zapVYSBe1MkEMNzPQNl4IR0jF/1krZhnlb8xZBpQdlDQ
nNenIPjtwgqDlmMNW3BJC50L4ahxJ993gXbQ4vCH2EHGHFz5JSeNh+tVenU84c14CA8HIMapRFpT
/Gqub7HhPimb2F4vcLQMSBS6h6JDsm6I646QtkVyD+UfnoLaO7yOxm/ZSrfbX8JGO0JJiGNkOTqV
0ArOju1ygD7h85D6Z+OCuKEOuamDsHf7To6kzb5fmWOdkbpKakuiaebkJlFzrYprBv5aU/T/Z1xg
N78ZCUeGWwvfHjTwbPa4gTrj+QEsDV6oQyIXPa4Kyg/3SxTlZCHu7cGqCmqu0/M3b7M6Brht3Qan
/KusVzvvJFGsFz9qjiI4E049Q4TJkmHHFs7432LpDrVhJALf15w5nhuTOJlGCOTER10aSnhVsZiy
KECbRs1Y72XtVIjKHA3/ulPzcqbMUsy+W0lPWNh6L+gZ/LUvSw5dcM2+xl8iDYJ+uzRyiXjqYoUc
vQGoZpfvQviJelmNQO+ifBzHrWDp3rASdMq+bC/638Nkck8GPAOy9KEZz222D/XHx7iQOSRey2Qm
LFKxO8wC0SR3tFSp/97FixaVwc537Arw/31GbheaICKMc2/OVFRtd+Aan5SMGCUc62Xk6IYEaTlb
95cNI8geEp0dNjf3Ok2BdtdcXv8iA16ztBf3PETBPA2c3r0BpxVbKHsXBYdJPeE2LvA3uN1MRa/F
oueJBict4KTzuBPPMwBmsALg1dJBwxi56TklhlCkI69dDALhgBkVJG/4rZH+juLlGhhnNE2qAUP3
/jbA4/erJjQXy+VW3LxvZTOHvchWDEQ9nRbiD9ToVnHCZLVTRIWM+rAKV+35JgmYqvjK5n8bMPug
yWRsKcKLD/SNbYm6aJ6Ujc9Kh/kFV4TkEoNGDxyEsjYPn8jcJNZMgWD1PXVRrUxoK5Ey//RMWkM1
AZgV93jRGy9oiWbVw7TIwoLOJp9MaXBV+a3+HDJw6SdjDvBlgF6MKv9yJA/9NvkybDDVHQoiTVUo
V1IdX7rYWI5u2e1yPGRqGGXRIoZdM42QmaicyNb0OE03gxaXWbpCNdI7pKihbzOZ1btoWfSZIsQP
hJDcEOViUM4cZ4lNTv8l4KNqe2J1oaiMEwC1I6DC+Jv1Gt2R3vwlxUerugbN3l+GFOKvaxAT7h0/
K8eSjcoJeQ2N/AX5b2+d3dZIzb4Yd9Tk1jzk5H64dzsOSTziIL1JRqFZK5TYEI6RIoY1ShfhHGl6
nWwQgkVLHUoVB6n31+HBICIA1DDCfzKVt3sL3R7mwLuwrfz16EGj2L98MqFNanHNUekk2w+WrvJB
oAKy9yCiDyW4ZS9thVJPxPWtJAxDf8R4HbJDahY4YMH2MAH4rPsFZLkMwCA3KOF4ab/TJy6qvIzZ
FWz4ZohbnMgOiQuXTKEihAVFBe3qnpoFf9bHEBiTHJlmQMnMDr0q1wHjX72eIqoBn0by0C/bpNgZ
ACz7KHVzsVGHQXpdV8k0YDoZ/nbmRa6YTWR6PZ9f/csHmSH+vvG/aZ91G62rjc/1KmVqk7G76eHz
k9f+2IVmu+oaQS7Xm59Lbgnmx7sXjhzk2IylmOPqupaV0iDHthO0RF+fZkGrnaoe0tASdc2JNwTe
D6yH1o68Dq8wzDoIb2jjoVqAPYV70NQGD3BkvS1p8NQsEKObWyafze0L4awVVGnB/DWYbDt8oyon
9Lmo1qC/yB3mD3uKDI05MO8XhZ0B3EjpjN6OrX+BRydzTPWovRf0LoPDWcKh+VA76Cxo9LuMhudo
Ja6/r0YvabUYJqam32faHtHzY6W45AERo4mCasY/Z7n65Mt3AjSs0xwWAGH1uXDLbwjsOF3o3Qxl
svzL2DLKre8aa2m/D2H3ma9aWFX4R8XgczKy4Ajfk5UrW0aaEOoMgjkI9ywGMqArXvqwjiifHXR9
vmV8tgDwhX1s/CxVzmv2JFb05A8GjFUg3AKIlMgSA+SIvtWuPb2Nmi1fmG0uLDD/hbtsbHEmGFr9
hlz5MEfMGE9JBII59u1O9F5ODqFLj89/p/0oz9NU4g+CL12xNs28cRNrVugxtmAQ1o4yNB5xI8Og
RwjMWD7SCCw3Ud3rLdoKtaiIHJsA3xJfvDSnuVQLqkj+1YFsWQe+6yV2MPaj/puJR99WJDKnDsTQ
Fvx7buArgZkR6r1vFNzWM26V6faEyuJGL/P72GmZdBzoAOJB/4T86h8PU1NMD9wRBoqIKUNoP6BQ
rroBlzZ4KBp3a7tAA8w9ijW7qbopfjfM3Vv39t4rJ/4l8/WkTlKap4kPA1EY7cdzwXkNTcVa3b3j
KmGCAsfz7b2fcRMeIKQytV9MjPNnXHERTQE7dEmrYFUa4KiZMJDVHfkwbLDiXnosIrAFRxlXeTlQ
HCNiIA0XyM0P6xx75aOlgty7XuagcIcPfIX1SIwjLqtMFNRU2AZi/UCpzUl+epDB8fRFWW6isljt
h9typ0EizLBXDNgPjI9tFXsFyCIhPXGchKXUIW4QmWsCyZT35mE+ObKuXDjeO4LW4zLOKmckdG0A
jG9Dy1yjqjt1RN9SEQzDuJvAgZ4ckqqpnC4nXvCzhCAJQUEmuqufQtliN0z12jaFomnN2p6Tap1l
I8jLx/zRABCO7wMZ+CPhNFhJX5TtEmulmorjInrlR7aj5oXyMyteAss8VAyFDI+5nKeH2tDMm4q4
oj4IBn7frxARxzD1IJd84XOxI9hVrIhelzfs1ZCAq2HrnmQkUYbqO1gADBcTwcEgWGu053Cq4V7L
LVoWH5HAGu055AV53CIhLK+Qin16c9YqgzrJrjkbSrA/GcIv8h2KcZ3UxaHwHMFvtMNhGM3S7iO9
r9kMoK1+GcFbQHayHB4ENX/Es1+9yy4wdtYZbaf2ni//Tv8LzqdmChBj6JcZEuqtKyYRpLdvM8wm
3yXeSIpSH368la6f4lZTSubBz/Bv0Vgo5o5f5ZpZtNy1Eu6nmRCJRfra9ZLDQboafkvzI9X+4qG5
QW2barYZOg6BRtay/D/+sKhiVPPLZ8WTcrOUr2BDdLEa8lcrdSzszQZnPWptXkw5rBCBz8tB1bBW
RRbNmT+gP/TXZi3JFxnOYbonUl4mOdYr12YGvEUMHINBQwve2+fk5eXbMazuwrBC8PII1/YlKuJ5
8uUDlGUn8mR+VfeE/XdZUjAkgtuPvMynE2j4vM8xLfi5E4aDGE2ME9fNiPb92eysualPkKqLYY3Z
+Y9Z8UAeggHmW3hQxcxGbv5Xa6d5+Tj7OfX/0dTsS0oT7iKkLPdqhI12ZZusKJxPpzC4GCJaH3MP
4DPoVuh+fK90AtoLsthYwN/9H1TBWymNe9F42icgchy+aO8RO1Iu6GuDrN8UHRn05B0vd+YtKQOq
8rj+IpuuuudGZL9qPhT4QFhRzN5XMUYWrsVgy30gjdTlJ9KO0GI/W/pNzijED+o65lx/x7SnwPR6
PpPuAfbztHGZeJFfIN4Soh+7JBdgQlPY0PQ4cbPp3kk+5OMT/gOqX4fpE1GtAHGMB/gB3/UyHwe/
Gp+STpCGnkpzWLRHpardN7Bc2ZNc8vBrw4KO+wGj5X7Sc8zOhHuyJty3563izFZGarGi4gGwHKlK
6hqAZDI5mlv8k9lo57Ka/s/OqTCdahC46fdkBa7aR/lGIk/eADuKSGtCkklrS9FVyZzZCvrEreld
LwSSNwSspTG6LBwQv9efknjhXiTSeAfESN9oiyOUPKsyuCVxpyR1wQmG0a73VSfXyOB/oOxL9Us3
yrVaRsn5/sXBodIxhyLNvyopdsFT1OEqKOiwt7wK206rhXUx+7u4TyepG/VlTyylNJenFkA0y5U0
K+YazXXXU2h/6ra5ErOR0n7+aEhwZUV9sqcglF35vTLze93T0lw0arQ/idyf3OBzIhD5F1wZfDcg
aD2/rQ5CCV8QBkFDYczMZw5XTpjFJUq4jM3GCzGyXrqB420y1XEhzcyu6UjwsQQREEagjdsGkvMs
/TUO7+sLYnOpCbKpr+PVi17/xPzrVPt4VUT0rj9IrsHzKqEr1cmPIsZ+1A4BchA5Bj+PMJiOiSjY
C98MdRFvg/MdsvvBXhDc9LVuEIZ3Zh94C6E7dpJiSfkOmyAndOffWCl/vzLfrur4TOLtCNDKD28/
wq+pPU/jmlAzVWoRkYOGZag7CAdcyKutzjxQcrJ/7Olc0eoNTfTIxa17SZwEAEI56Bnrax1bhsNL
uE5UCwUg2DAG7jzuehVJKs5Iv2rZQ8WR0bdbIAaATyDWOmXxzMSy//Tu7K7dVZebHqLmW3+ha9/Y
3qh9VxJOl8NoBg45uJTEpqKzh7SCVzkA20SLaJDRgPtSaq9buTgVv7EbuuQb5EO2WX+vmJMQRM6/
KLQvNuy3LN6qoP5oHtQV1+cA+hjMgVLFt1HSGGdKH/G/ZDrQmT+CWVMs7PbcbMJ20RPvrZvB3LLp
RpQLJiG4tjq/7S5+cnLEMBCpUJiHZ7ifRqHvisAy0XttrTNGrcvPfXpN5BqyLwAfhQuxd6zxudrI
3yhg7b7Y9D5wS3f4FZ6bkRIUwVYseX9nscsMZClWoYX5vWBbiDHCi1773ECxmHzKTZvm03AeKwBr
PmElXcH9kUKx8YGUlS86NtNhzR8bj0zuNHWDLksMcjgO2PcDyzDuRO0sl2I9KMm/4aPe7tDSTqWR
Oga75zUzuWgttDudnPnWqFMBmuDAa8D1B+0Ozp5h9nopmLDa/2qniMVyGj7tPIzmYp+ckXMkscqi
fuCTKG2cVwz2gcRxsQ+Ep8Zpz2PynHgjp2jfIvDI0tHE4ikCSWvlqGM2JkjWW8e6hBTi0ylQpkT/
gCn6PhxrSNlksjBZ2mU/0Z7e7N/DZSa3xw9g1TiZj0Mn2A3FufaQIydQYNPjMkxw6eHy98tAZ7uc
nZd9uqmrKeBRZUAraeBRAbI3rPwfi4+jgpIP56wWD0XTOlh/eS1vBJAGmSpL3x23usp4qKcr6rf2
wRcT+C6QX3g1x17p6Xv3A0Dr6l1tGD0vMwA9v9B7J35v844leNQXQ2284E7wlFgcbDSO0oC6QB6o
oLqzvEuezGG7DYKHSxO3G/4hD3Ic1xXGHCg7+yaiivKsUSlfyhoNHAEUoYWnU1I8OezTk4qP0JO1
VgIZewoag84fqZGxtbaQ3e9VEawLwZVG/LQE3qEYIduNmorwnm46tOYcrQ8sx8L7dBQbtABFP4x1
6Kqr6il+5vAmPje/3ZBCY4LyO5VHsNXv/42xVkgzrOQRyfM504gtSKXLYvoqdvuW0n7lKEEegURa
C7SEvcNc4qZUQDGOHNJSFzUbRfVA5BZ40+q2Gr4gym59reHAHN15APVg47OfFxP/JQ4vWe82Ctvy
2u+HIqd64Je5d0ZSaxi6gy9E8AjyYRu/HuC7AyBtE8UQnfFneNbpQPgIpZB9gbnuhTNcirafWO5i
3N7aaaw+Z4mazhzpO3PWBv4Zq9I3sCDkct4UTM0fdR6u726m1L/2G/TqgPVF967O7cFoMOgrEc5h
Ngg1ROO+uV9pZg8N0jGUuHsuLmaZXtFG6pJpAxZ0plX74wRtCQQh6QvZxgewzsZ0r0kd7nTePFm+
IiLv5C5qIPYswGwlEDhnllRZyKkAe9gZ/qqiTokG/iGPfnh0NW0kEXreJ2xoGQJUinYtpkB+Oo7L
hGSQFzNWlskNgSXEwCyHA4/CbZGaqw9GVcmmSml0lnPDLyiOu+CRe2k8UeENUr7OpCsS1UuysDPn
VrEZrpEsHjZEdLHILH+ySydk4XzoHI/UF3bxcx2Ep74P1SOD0tgvDHtOJ4VBezvUJMgxaJbyu8N5
XgFhceJmwYxU6Eyxd+GrdjUZXa06Frd5QxlxDSvOoLOCOpByRHJPsZBJIOEX9s9RtYCkHHoD6k/7
oGHcC3AN+WrOSsQUNXWp8+RquHYxrB9D116MQcytMI1dKTDOHpSXBwYWfyCvW/q6PHuLPNZ0K2wA
y7K2hFUNx8UdZ1t3pTTkPhkc5CR1u5DpzC4Ylr9XrmycTrUbOLpPFpbqh+H6Rk8XXA73sngJLefX
NM61WXwakFtGWDeHAUqO1EOqlEGlNBM/hQbbYYVyCo+7DcL9MZZ3nZszNn5KAoVQhna4sAUYcIrB
aSwun1Vr5EDEuS2/L1/2bv+iyq8eQgf/m0rCTDGVdaiRCaYLOBEbmJhAh+PdBz3SdmVgpcpizmFi
y+trwQSPXhq39xvlhaxHRr3CF2QUK2iBrUoZoObtbrikwQhhq1xrcVJrd/6Fdoix6BzoB8zn/ydQ
n/Dk8KOfKbN0Y0ac1a/+L2f5WRL1Yv17mjjCDTEyUf6aWnhDOxlp8/ZB3IzDVIwIvIONSoRi1n72
INFyGK6fTdrLV8HJktB55PsMFKJd9QZB0oV09684FdiXMH8BPl5ewlOogycKX2dv7XQA26aUGcdJ
mAdZVCjKBm8uiFzNMBLLwTqJaiuoJXCtr8h/PQ0+1JOPxfIJCM9uyMyt4kSypT99ekTt9fXy0TjQ
vRD0wiQOhmmpP1yHK4tnHpy4TbwnG4oeQJmBw4sfo3aWfxlyxQNVFIxMFfzCvGXI2np9cda4DN9l
roy3q36EZa3FAXh93cY0kmfdCUj/IQi8l0bKpbIXicBKB14QRiopkAJgQq7WXpDx2DcqJrEWSxdD
B4StfH/yREXfcqsVwRmvSqKP+iliRYG/yKSceP3SfbTHgc7foaDVvNNseCy4APnCCIPZqpBUgfxA
SL2rLJhk+UyKOGefmKGsQjomVt7ZxXJFl0XVz/WSL0EHXGKc12pB/bfy7nOWgDf+cPfV2V6I2KEz
swSZ5E/ExcSTh1CBej7d3ZFEZEn7c01hTIpCTmpfuOe3TmAB/vsgBiRcjxI5GDC2fYIWisZO1XHo
7Yaizx/chq6t2uWwKLVygxqAQDPt7cG8bJQu8qjAG+R6pg9FDldC7ycg5uMaEKEsupNeCX9sUO4e
N5QcN8yT1LWLov9s1RJhRB/pSUuDb571jQZ4Q3EcpaEiN170MUY6ryZkBhekkQoWbTZn34zhT0ND
vO7gPIogAPBvBdoEEuiDNHq53wfzE+2OSYOOYMPSrRb1WhO0HPSJhbm/JcpmeczaC4Vd9eYRze97
ZI0UTiXytEFAMEyzWp+hhUC2bkgar9Sl+dEO5448wVNAVV3kd5925JidgoTxDWVHvkWGGH7Tn/IK
MuS4XFQzT+qVJJH2nlQ/hwlrugvGUEA9kWIhUMd6b/EKYYBUC+eUTw8cehr8Ufplvnt/jSD07zNs
hdf9mOdvME66AdfV42aXgCqr5gUxUqrUOF0yUoLFTFWbeoNWbSp1BbCX2nY5PlofjWfTQ5uriS9t
IglgJwaNt34jrQx8zre6mK5aaTcGnqaBNlq+ur0+IrgAhR9tyYTD+7RlQpXXIbHyVfThL9q+gu2U
kdz9Pe0M6c3vNJLvyTnqfIgri6KWoL2m5mYgdzTxNrEJnvZga6dRCsKUQJeCHdv4x7LQ4IunYr1I
aMSjWtyA+PeRPWeubAn8jjJ1dqurLg7Rv8pUNEEjFJCVe42SZ1mNPNl1VszEp+7Iy4nGztPC7UTs
y6oUzu6Fi11IBSM8qCHM64KiGFrzddi5ZAiRV3sLL2F8mM5NH4u+/c+0EsYiZmNLy8yNpf6Xos9x
sVmcKSI61FqFQQHqiqz979Ni/YwQsPBY0wTFTHbIfiyTR6Tltn+dkjcRKKI/t4XhJV0T/8erVsRn
0rChiLLqv4lAN7WjXlzk75ld25H1VVlfx4VXUFIo+TJ7T7ocWQFmdEqS6DZZeyiq/0kCA2/1QAjb
RyuY+33GXqCuJrzedts6IQRI0GZk2WdOpS4KHjsJZVTAj+xU66Mf3nc1BXHVYWxQ5f5T0GaWb3Me
oDIUyRsOw795/+M9iFtcfu6gaiE09aKEQniwc01QtgkGgdMwnobg3yLJ04aJyeknMYccclcsEten
8kkyIjfxZf6hkIf0y1074lZJ2VOWN3yAFPHtFA1BHw/zbpeGNbEiY9vJ1itbcdOFQ/Mkrllmfp3l
ue5A1lzoIeUduVAtbtT+YcJA9IbhY7KMJLIaM9yQ1+5nZb/vfIobKbw1bQlMFwxDMajFVBiJr44l
7w0r3+4+WzM1nSJzm5Tc2p+Bkc4haa4148cJI4bQSbve4HCtDzxWUnpO+52/Ql9NvSEgrrjxbcfo
ZPS3EG8xgDzMlTbTIiL8Ek/02VL+avg9zg9Con9fezUYfuDaSnJ8JCX7VluXrfjAsRbHFzwtIp1i
o3LBQEJwzdRVBGbVTladzNn/n3g3+9FPmxgsgCoJYjEtnXxTSsX4S5iDZimr5j86bAQOfZHhiGnd
oHcK1QQwz/DFvmVdFVisr1wy3Xy0uGVdIsDXMge4T/xP6aE3cjpQhN3koNRhChMVBbQSLLfpedPy
8E6eo6F2/ZVEWVkv87UsLUfkKK3tO+rLcnvYfhXhZ/Z9XaAlZA5PGhFBubPZlgWzrK7XPfjlcf4w
mi7dwocx/QBbQUykH21JyXRDmt/IAE9Tb8sH/o1bGE1fz6lGrnwEGHrxYUXmas/FcgQKkeI8W0YY
8k4F/Yoi+tp0BN/ACyI5+q/puOIYoi4GkKfepIYrXPT2Qw7M2cAEfeLGUef4ngOJYTJpgf9pq9kp
w/4/jvIzrvcVNMUlZCWA5vEOVWGR3AVqmDVKLiXBErbbE6G+EydDD7KxKZUHLPWvuq2QPcwNLi/C
V1Tyl9TRrhyiXsP1JX8tDE2zfkU5cdZk82IFyEJMYgrprtkUZKGPUvuiw5WlcWvMmuZRi4T4gFwV
2LCtSvNG8/BGgGJW9QfCmyb7BOScL2IBZIzoXcG0lt1+CfVXo4IjguuttLMYGdqkpqWSTbnvmZv2
xv4ZDR9Yntex5tdrzdF3IRnj/exMnlPSYf53UnUk33MACIWnI6Zt8szzprajvYkW8WabOgxJDW7O
ZcrFyQqtTuvX+Ts84GmoG6FG8qESrmtz9uv6Z56dbFB4yoOtBNX6hIoFNTIDwNGTrBnXyKirWwOv
u7EX/wisFhHpwI8Jo5pRYLsGRVTeiIqWHMaunZgxWNIiKvUrnniLxKYtqVaPw1NFES5sg49DGqcx
NdX/kFN/nhTlo7lBcSq1a5SK4rWvZvEG88sPsQoKuSOz3URteeCbkc7SEeu2NMBXmTb00qQw1lQE
VpJ7uoPl8Qb7JuzucAVYcoiZR9sadVw65QUw6LOFiEy831VxquhUrlMXI/vb0oZ0Encxg4qbPorz
/yjXvNomhcJrEPi8qb/I+JTQhxnLm8hA1DI42BkCEvseILE7OEvL3GJeya6q4SMXRGCgKkKPN5Tm
fqXTDOjHhAbH3/vJZscNYoV1DUbSsVhI3hxC58gToVrRP5V7KDSoA8YNH3m40uIGqC14ETqE5jMB
5aI7zWWRPMbg/G8Os4c9LHL2aYatiKbEitr79YG1Lud5z0Lrgod+NBcX/whv4d3ZSLFInH6atVE9
UyDsTTYWmeNiuUabns5APlQiPfSYkgFIOnoa9yUj0kOVvHLqaKI+IvPUu6UR3qmjD6M9gzabK7pE
GGkqJNMtzlBOXEs3k/TGRikQEdAvTxzAOA2BOu1r1dHUS5kGpfVSisjLMAIS9SXFp6Gl4e4jQJKP
mQz0vhekwO9EFMVzy0DEwI2ZR5cERpY3xzqbmo7gfciSqFiXUCXsvVv8+IOUTiwSskCBcuIjey/N
VT4QLpV9544xoo+8EqTaXS9S7Yhvb6nsUDXoHKmfXzMwkbTtvKwygnY4kKY5JqeUEA6mh9LHHwzC
YnU7U/3u+vfqngPv4JmEPf8ICWM6FEN0G4KsvgiB3ynBdXS4uqSJIYHiNzvZugyx99yqVFmrQY0s
KzT2+jGW/4OAD/a2T1C3AJyofv+yTGXdsqAHR6mR35VwT0x7g1bMx+R6aeMoiiUt0oJQjm/5yGJq
HP1fD1HVUeZMH0CrR0NdAuxc5oiJmUKZgKghAzn8ej/cGzIyeP5/EBAejkxlAiKz7pJSi4SBZfcp
LOr/y7UASdmr9ZMzGG0lcyt/1hpiSv3Z5/Zs1BrkS75zFC7n9htu/pe67ymnFi9ox8+IJMT0TF9G
gXC7Ifcrn2Ld6DMpWnGGUtHk7OYsq+zyy1ebwS36foJbRKh3bTrrW42jQQFaMGpV1Q3f1+ueJwf0
yjaJc7c7elYSKz3t66tbEWEIsCRA/vMQ1HVwRirQa74YeFahTIPi/sfoT6+O+ypMy4hix7SwDYvc
Hm8cgvPOdJgegmAmwRjvcrlK2jGLmVGU3AvirkpweydxEr+Oc3ae/bEIssHTvETA2DnYEIm8WokE
D83oDPv7GpPkHlg5wj1ny5QwW3oQ47m5Z4XheEHdPzwwRORECengDCdoBYsF/tVVReTvafaclwpJ
K1/2wsp8ex+jR0ukhgR4ufgWgKXJ8vsPZr2VzJQI93LSVfDXdxS8lFtESKTzjGOnpNhaujZPirkU
5ybC+90AWvvPlk/ZyBMSbDufXMmPscCm6VvA4tL98xogDep/wcuzefQaDqFvpVvzj4x/tzhCtdQl
d2WlDQsSnr41wKalL4BE/F8fVGClee6v/7GVOYH+2FHdf3CyYsG5gxY4MOQJAOb2thAWztNwtsdR
UirtHf2JntK9ku4sS9wi9NnULpr1KrTkXUfNKg3n9wxgUbfeWlRYzege31QNw0nRjlj4PUdiHc+X
BvnNyrrclbAwlE8qamctPR559j9Q10X9dxnDiZE67F4winrx7dSTAIpMcJxuaI3HMaK+JBqRBvzw
zfN/+sWEE72ryJPWjMk0qiRz0lZhnCbrmpp6dGQsncuSW8jvx425sg0IkMjsahBjtzLpZ8kp04rI
vhrnA0NdS8+guGt4yFEdYd7af9EULHG1fiDkKmqkKraCY3fNdWW2scGQh077S+Tjr73oeW643DV/
Y2TNx73UwSUQzLHubEt/XHCcfTrZVKbBZKlqlTQ2K+o/XFUEmTALEILG2EXj3WTbSUKnlniGSGux
tMyyzkE6+bnGQR9Q8tX1dRUEM2bZZPMP13sJdzZueEaRpxWZlVFS/d+Ro+d03pYpLcv1wfWE1Y1p
1F2AQpkojttBNZkv+IicOufWXMy4ltcZwHyQVdoLThOQoNVIB9c0alLHisCBqJ7hMpUsIO4k8xUi
BgaMREHZVOKBtcaqAJwG9PLmJwEgwMHvB+8WAgHXlWpwt21LeS97SntB1uivPw7ZBAOyG64V+wL5
9ecdp2VTGWkTv1OwQCr+TGqirlxWIGa47Qm1Gp5FUmW9gWTRwCB8mGukXO4TeL9ZpaQ5TZjLrTxq
00DMNIMCECzkTN+QWetnOXvfGluIvTQ/AANV1ps0Y1nozSZPjmus53RxbaIuJuZcRluZLWd7aakf
nixss3uob7UQ7UST9u4LShEgeoQvNu+yM5n4OFiKZl6SRd+l4mY8b34mA5FV5oSuQRKXsgNZ90vi
KrRo0KUwNQ0xhQPI+/RlWrbJXBnogamC/Q9FLdufYJEvaHpKQ/Zwr6JCUbaonB7RnBz43XIOe1Rl
87A2FOs0YO+i4K1+ja2Q0TXdJO5y6PHEDhNJibmS4vaEpqSWbQa8L3nGqT8YNzdCPW/nZn7umX4U
FXKCdePqTr42II7GSnxHsKyKYdcAJnKE3nGD3jjcMoHOSkQNgxUmJKWHQmizq0snLqenTFN+Jsh8
TacRhT3OzcxiVELQJ0X7vcHaleim3TRGarberqTgEDbstZSvUPY7yecuT1Mi1ju9CnIZ4O49Ms9V
ee1DHyxxzGztnQKz/0a+gmPk5jS/C1QqtP1kkYgbhbBcXMKTyxFXIl4rnboGJuaa6uR4bPbPVxOc
r5qXj2Chag==
`protect end_protected

