

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IyCaF6+6roRR/z73FG9YaF0d7dULyJHX+GoNBLXm93HBP9lCLRfrto6vEw3iGCXzK5VqUo8LUzXz
LNIjSmykCQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ars/zU9oYJUMCyRasaGmgdFnCUXaN3o1oQ0fks4+dXZBJExbjObt0eQ4bTm1Oe0kx7bwkjVYQOv+
UQ7LSA8+pLx+dSrw76W+fhwmbjv8NHk8HXyQr62gS6pGtiXKgK736w7+XTNBA1vQ12Yb/XlI+UNz
IEXEAHZPmFtNRS82+9s=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ypT22bO1Sgj7GXF62sjMcbzRg1ae280bxZhy4N2bQAjzULe/jSsJYy+PGhgDbzqrDKTpXiyDtZkt
oD02eLDdRTGllWcMLfmAbMcheBPHnKTXt9HAhXv063PgOy3UnY+4gioTKkh80haiBvLJgatSPifi
YQpeTG2uJk2s6avI9DDuJWf5ytesbOIq8rdjhkKeFXOVJkRrosfyEugTvccoc1Vbfz7A4F2wgM+D
zQAdcf6ITFXwFESPDeWg0jBH/8FT/oGTumoj/JU8XybS9R37MtI+EqSG5OCB5UPfR7kygCRxMdqx
w9C2YvXXr8F4xw6pVMAzGqjHHzZitlsy10wY2A==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iUt+lAN3QxnHPLXCGVB/8iLwL0mQDxrC2eKEtZRQ3tSttWm8FZZIS+L6sXzOYBFdcvxa9yav+Skk
gH0KYhQwN9nPnbBmvq+pv0OWmlNAuJl9BKYeCRvvHDm6ZFmplDtVldoTwk3H3W89FxmDdhSnrp8p
y+EZ4Sey0JKCjHzhKDLb9aiV4K1RcLnUYIHkxt5NRemjZPNHJtaHYmmTYfrufApExkwl0g97mMJh
/9bAzlLXFYd5iRY8cWYOanmNtNy8XdgpYQ9x9FO0bReaxTyYk8KeTd2hcuaOnipXIq1dnLyNcsQ3
oacpKj3c+OCD0yKkipipeAUExSzqLkMixzBzew==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JjEJ4N/hIu1WBDUjIMq9s1GMccDmtrtckrJO9KM4FgsQ0FVnrvs7XLEtH7w3vJEH6mnZFK6gx+Zp
Z6sD/j5+c1FsEF5qvoz8DFaJv1SA0e6R+wJt9JWLiNHRgEY4FWJuMy4GeEzK+JXZXpK3GXkLR7a+
1Q6HsnbRSckp2PGMKP0=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KZqHvWv65FrttYAd5GXAxNF6M7H4sPlwsazq1nKQJNzvqECgNuEcm+ZAEJdmD/ayAjxuoA6PeUTI
0DfZA6W/dyVpZBZL701cNaCalR4P8jm9gUNIdKoK9h5ACM0wpchU/5peA9dkp8Q71W1JfJhVf6wV
Pfq6P6zpkxEHamzXVJgMfDIbIUtVkFo5jpozvANXGvZy4NvDF+IkDqh9n1WhJSFw2vSTSWwOc6Os
YPCyiHHgK6fUeo5HsDm8nUZX9YA0YMDCcn+IsvxAoCbVnB8MyuhCLYXxAuS9RlY1JV6hAzEQMCpq
3UPMC6tAiYJyvnJO2Ue+HpfWovjSQbxzMY99PA==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vdoPlvKWn5Ji3Xo88zOn99MOAqtEoxjAhuAza+l5LAfqRqsliwhzcGFkAJK4ugd9gKm/M3nHnHPi
/PzAE8cF+f+Utbn8D4EMwG4W0Hif+wOLC02e4qH1wSqAV6WWUm8H7NgadjCJBzXMdZZG7gjGozFv
hvjCKrn45bL0EmR7wl2Q8vZe6J7uihKTYiousdVwB8VF1FLUjPpp6Af2cQmPK82eSrVw0IFHIKqJ
Y/a7ujGEnXPRmoENXb8yibx2IfMb6P5x8SvBxbWHb/Z6q10od4kw4eQyCm6rPn5iaTS1SDweCTJ2
LVJYDuUcJm0TAZrXENpQQfojrfHxe1bol/kUPg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_11", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lmo1O/nWVfjvEnWKtJ3RCiwGaUnm3M24qPwY+KlvzkKo4sOFoccG5hcg/sL3BguT2Fqs6upec+/P
lgkR9EpxAHK53ySSYK2Gk+/zJ6wPEAQODMbLtASGTteC4atByoS7g+bnqTV2RCzwQJ8IeLVm63oC
q/A1HmQVWMT63Dha7RRPAWhUKfbQ6Gcxxbrt178CMgNEF8fK64fGKwpKWWGSTZdOuCI6JYCt31CH
jLLgd8XhBzNkjXVlUX1wvTnpXb+ZIkY6TeEL8T+DC3/ZFeM7LEjbf1gPEnDR55V2FW99uqAyh9B+
/sRPnmh44cDlw55G3HMOOIAM5c5/ybP6C+lmBw==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ByXNDvTKDI6gFflyODyOtNqLQFU3tDtRuDnI1QTYGEkfXSRy0PtPqdzLUwZOdH6S+7qVRr5I7hia
BIzMOSTXTbSUeFMET0ea5G6/osyZGxD3vhMq5mc07fbIvonlLCBhXZc9zsxWxmrQIUImWH2twnpK
slu9Wg50/fudlPoBjMVmVGo1w8qzoBi/BwnTzF3og4Q8HdJMlsbKVZ96oAGGsWVhVVGjpde8xZC+
GvqB6jQ2vMmNZJNkyZ47uC4C7nyRet9HhKhT7lFrpKi/HydIDNj30XFaozPxFCtHrnxgGQ0dtM+E
UDFL1fGQBdh4xbe+5S2zrlJKxZ83MLUKUmpM6w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 506800)
`protect data_block
kwxUQJS2Hj+s1kscEYt10lYwwcGDOV/69q6MNw/cjHApjLtE5p2HbmOsNC9XCw2Z6g6+mD9Gb5+t
GmqRTTDxRF4b70GtPYfnUOLOzmEYtQQxwh4izH8BS+l9kDSfOXj0XmSQV6bVUnhLp8FCk9WmCYfo
c8BU8snkWJ5NvyJpbciJotfhqVnSyS9nZE/Vtp8GbIFUbc0reTx/o1iADsEkCJ/CjESlRW8/UDmz
qJFg2QsH51pTHaUv/c+XiPU3Pm5NhvycxwDTuzWADbWzqDoLP0L/NITT1elSateJcU5NkH3PM7mK
PqKdqnlfehSc94JrWM+nPIO/d4CDEIapOvf9CnlRdxgBEgzMnvFoptIpXMgZhEzjZH+XwzKIC3Oe
wn5NoIpGVUTN2oVaMiM7h0Be16P7esZvjUjjIF8RSw2YXNmFnN+G2su08vkqxgi8pjSeYkY8equm
kLUM7wz6zvOs5qnXs29wTLVtDXQ2ArZXu2dx2uXSM0qN4j0YIJcS/ZatNU2YuQbgNwYgqRx8YO0J
e/GPQMJfQqfKuhAeiwJZsG0ayJdYxOJrb9CcXIHxhkKOJPuz8ONdotHzVb6CdAfYULdczvTgzPew
+VHuZCZVkV3s0pVIQWIrvX2KKKa19o5Wkwt3xEMbF/n7nBLarEn3wm7uLoqiQ0rmUrRZd4VxFd+H
KAXC0nIVSx/Fs0fsWcYA3Soy0Ms2T/46HCScFzbFRFCDRblURul2+d4++6hpIh9+WZfHGlxoElmH
biMFdCRTBgtjVeKM3r4ntJdWvHozA7MrwlNKg9O/Jo4+npyraEZ1usqM8lOMnLcM084iS8oRsecf
pfdiq8340rKdVmi4AR79QnvUOpthgio7ZyLJN7Hzoy5Kx1kvfiUsw4clahr1Ibj4tlUknniMStZs
MhekMwRzyoXxvIRTXZOefbsNCH5e2yPbecT82O8r6pGjbMLhnu7jiCYUxucY9zlb7JeYYbpih240
Og1gYWrsasf2aOIi63bkn0p8OsATJZFySWESXBh6ZgouBAUyAqN36Wv0ZnQ2sBSl3/UluaJwWh+C
p6MH00K2BPaqoek6tchzrriCtU7WWLXGTVu47+zMHQyW0YDhtk5QEWvcwsgU0GReGGqzKmNwddXZ
EasODm9UwZakocyp+/h0xfrneXnQ4K8QUupaIKhDIKspjVVprfkhFBBu6kFS63/68Cdx0su7iJfS
1ybhDXtZ97pxE/RWENkPeDfiyR7yZWO/WIpjIrrDgfQxkPcENAzWAjBYbxCxWu6aj3+eN9jIBe4b
2M4zFfLvtnrctUynBOTfh1T4XR+k/YbAHXizNRR8oKiVR5LeXkNP+OEdvcD9iVoNTf0wALcfw3ew
sLRUghQaxtSW0iSaKnRoqQ7klnnNZr1BkYp3n08iFicJPHiJ3nE6m7IziWhxUhzruEQ2orNpz5cc
IwstMZb/Y6cY8bDdY8uBnwIQh5+zziXifcmnxBp5ESzCXOyOS3eDiMw0dQjOIn7T/R+q6TVsw8ul
167rPuK080Mx2xBDDGkrHbA7hzZ0nC+Uh+eQyK4noXls3yMDu41ALJpjBCAdHiGnHLK74KFY+H+e
Yri7tsu0FEamRwuBzgSWQKi5GmFjImgqsCNMo1x3z/DaGNIhXTb4MSS1cnbD+H0hyOBYFz3UgBvD
UpckbUS0sLr6x+/0SPe3AsVk2YdMClbO1Z1HZj32o5+hs+J+8iwktc7tH5SBGyQg1czXtNikhI75
rxg7z/qZ/xoLlqdTLAVoRjUWSxSTiRentqRaljRdpu5NOIrQIck4D80JnTby5Zy/jlQXl+/TiqYC
tzmqBEDOzYyRy1NK+QIrd8rjhhPd4OdlnU4jMJY1XMDzVx1RIcLVeCg5zXhxnaqMqkxlwi1IjfUL
QLKjFesQhckZ1FxwLz7I2u3Bvdf0xfW2YC/PEbZ9D+XxK6V3jyWlniC8zD+AOwWPZsywPynHv2/q
R1fJ/afPSBYvVyKf2gqccKNGVRF2ZwwLzsBQP4Krm2THLg+enKt2KRv086A74EKbNH0AtHyWgCaK
RZC8iQmQieCgNzLhr8hH6mVT/l6T6Uy0YYNbVq1bESDdWyweUATtD57R3pMW6g9cP6fSD1uGDLlk
CdMO+qSZi7rWQn9P4qm0XuaQRnvyBXjSyQUyJRWsKhfFOq4qa9HScSRxn4neL6ntRqABpWFvtcds
mCsFvTR2ZD5BfmfcrgFqScrV0QPkK487HSi84Hh2KN8r3W424YPvmaE4U/vniadhMbAqdaUYklsU
D7csrAMaKDjqTLLFU/LbvyFmKHrmFo/q+2AVhAmtKx/G4yAS9lg9OjDleQyUIoN62LRpx2frAu6F
ppPHOvhSn5/NnyRwxYfdC+xUB6OaUyOj9hU4l4s/1/0dKGxDkdvjywKROMd2e+IRJzQGUxhzsc7G
5NzOy6QaanoheHMhx1HEoyY2RS8dYmwToG4D+3yNVbMeQvL61TRNm0MpM4r8KaQLNCi+WsgaVnRV
M5cUOK9L1d75wIeJTvlzqQ0vrbdOglen53LYmSnK1gD5nGrIBwn1NLkDZrNrisX41x/rD3fB/0Cm
HIQvoqYJ2YPftuWjMyPFwLx8aLclBJySxTRurJa6EaDucvvAhyp6zu7nx9aryi6ctNUSiosjZBwW
4Pkki0SC1vuy04H+IXzaLCetbHoMuKoqYDUjFwgzHvvTetYPMZuALpKNwWk21RHJydL+gbujezCG
yVTFzKzdtM3LOaVGwo0UGFMcopZombi2AIgP9H+6RXRgrXhq2OERzlUeSTxnWxJDsCUSB0Mg2A4u
NIPot69XLepiTvwDtznWMvnuRdl4nVOY81+RN+3aDJ3/yTL6CQjqyR9fNJ1OIU1xBq9hy79fD2wE
5j2Hi0rkUn0bxD/LZIC4cIpBv7G0OuCZ3blT3TP27dYqmm0bUZP1/oZMY4mYzyuTwjv3VPG2Ikju
8VvA5iH2RX1k1ACK+TLTJpu9gs2kmqyFvyNeYqDDYOfqQMls+dQ9+rur6Hm2czxThjEw33h91lCv
Crm4NEhDShXxwsQl3fGk+t0UUoevytkCwceNzcY4DcXTZaAaBqy9uRSM1qRqIrn1g3WSPhmdVbwH
bzvXDqnQWqdB2n53vplcSdaX3vY/80gsrurvX6D2o2P9fNmlLseDKRmPq9tcYbn3tx218Tb/XJE/
7DWvu1zWogouzA6coBTcuqZ27CzZStePrEySjZ1siZTLSFFDKoAZgioFxlWs/xJDI6IEMFsSPkln
O+t5thvyEivt5PbhPldaArF9L+ndCz9dXQblnlmyGgMT/dWHVcze8jj5HAT/efWZIlEsofEBZwn8
rma14+5rVRfH0+e/VbSUl2+JgeywXvi5B4UOocD+49cf/zumRYch150JqCfRxgEgqYVXLtofp0xG
4TCODqOrCSfgVGyd6/Nux9MARn+EHP4duOrjv3DPkm8LC1YG0uqK+dab+dLhCzSe/HoDG19S6QYw
LZJXVg3HTyv9UFFOIyxG6UIy6Nfoh4HEriacTsBD1CsO6NeYToeDL0MbJgu4mI0m321ZkcqOPemU
i7E32DvEEurlcbm7Z+4mcb8YMgUjas/DFA5U9NmSTePIKLzfO/WjJ1sigczj7O/kxx9PfX30FsVO
7wN7kCoPRd01Ndo17kz5YvlzIxwhcqppHdzCE5hXX0ki/7Av4WbDdonfqOYqfzevl4GMN041zUce
lOtP5JM73cvjJlWzID2ucxB0qRaFf8wKvX/zUGwCFeRH765bh0ChKJORjo6u6tXxXkZeJ/B6YRt1
oICdg2oztO7PSmnbAUPDrqSoCd4l6AZzQPLQSTIauUkYQMeUt2AZes8NPOsiNDLwDyT6YHt2D1Rq
iGI2WptXub1lMD2F59osZInV8gtHvn1h05mUoC6tifyp+UH7ViZuby1+Bwaps3dSmmOCbk+RhOgi
NtALuN+k4AeUReAZ61YR/FqVYMn3VgQSrnRiD1+ooIoINCm2mF2uUG5c25Via0OOm2KTFtlnnmcT
7QtojQR/bjZ9MtBD+Bsm0PIKTjKGgxgfGQ5ceMAPdEyrzU2bQUx1AoPCZYXfbmVU5DtrP9jrok2g
71sfVKdw+7y7UJ9dwSplUcUN7AOTUUDYx6w2b8fe6n8mtk1Wd88xLCH8PBbo1Y1FzhoyCK7BtFF3
kyXyQPXygBWDogFMtaqrIzKYytczaReQZCPQby6UcfP7HNdOJ7542xbPqBKSdO+O+V5dX/XywrPu
lCUcw2TeReV6Fnis1unj11QiNic3AVbpWdSIC4ws4yKexB6TqagOeX4E+T1SBZAwPkxCtD6/t38X
Ic/y+dKlrk+0lF8iJv7Ymhidqz6z/VIC449fMDnllUT4wTW8lVCftRW9RJAUHdnIlF/5MwzYtFMt
azZAAQjhsnfzqwPQPTA5w6BQUidWLkRhPiqwufr1bhl2R/dcmEOAI6nhf8QIWs+waRrVU/T4qDzQ
yU3mXTitkGKl+1UYXSrSipptq6sPlZfmmTzMRoLvT/u6B+t9nwSZ+nwWoEF1IZ84aqdNQHb4OAQv
nCpELfdfoEjPpgqp6jbUPdFf1zEXidsLjOgD9CszdOdTFl1o2dxOwJ7tG+w49C8vSjLugOTPvDcV
bBMJGqVy+U0+DLfohMOlC1Q8E0ry3tQruCQgaOVTFb2gL/6Dpv1hYgs5oIJ/iWm0+Jjw6FfcoWkS
iOlMzVkxLAqtmOUKEqKK3bI8C/I501IG+qQZ6Hj7l7ZOWjA5xEm0+iHtt0jmNyzVNPQHuNiMTqdV
eG/kk6V64XlthayjIq9Rq1+FuQ9BUyFVnvyOA1kdgUPiTZBUNuDlqbD4ukXPK9DFkRbnyVdmHihz
37QQPsQgV1o2M+m3tcMP8hDG5EoTKhFaglhzUsPzQ4vsvdeSL4ypr724w/lszmJmGpiaO8gta7XK
6Ohqa8M9DPqXvUjEBIkdYUonuJKKPVZY42505R6/kBdPudFmJd9qedRqwNk3Op/Dpd8DDWW3y0zV
OKE8aCcWUdHgvPi2W7M/ljui3BJJnz7FSrClphTDM+a+V1a4KSBLEGsdbNgBmwLAIEMReNgxd0n9
pO8Ja0+Q7/sMb2tWz6XlIete09HJV/fzhV+M4hbdbYn+kq8XuBGFStp55E4TmpHvSp92er5vynS8
kX1U+IwlmgN/kvFNObjpFy1R2sAM8DnFSRI2KtO433f8lOzV25PcxszLI2WdSqO1JFlES1vQ4NuG
GlG6v8l34eGsSZ0jor21QCC4sxW+hfwrd7nUfFODCM1EUa3YWbBruoE8fJl8yx1ZgMpNCEele4Bo
WH5MLxwvd4L7cQt4mg+bTez/DGWWks37oGL25Mfwxkl+fillfdJOi9m20A5inLDQY0UtHarsg+4Y
MhfgPAfxOFI0GVnkAKkiVvyFmgqwrcCrDbe77arWazm6JobFDbBaNC0EaqW7KC1pb7Q7iLvmvYbd
xHu1/bM5bXgLrTtf9wSREiGtA0h9+XvMmt9UWmyHTiZ0EXscy9d4+z5XYaiyOpTqNIOkMR71/d5V
1qXEsFYPP9DgMWnQgL5kdRpots5eKC3DJ9mGTPWKamF8duRl2H0sDPLhG2WSVZse6H5+D9hPwn1U
Tkk95HrO8XIoCQOfpPfxw4zyLv1El93TJDlKDsfjsId6rqjuqJ8ih7mZZhI//rgslHB6ll5QpvXI
dbiE1we56yxClMEzhB09GsXhjzQbjpV7mh0NAx57FaIYHkSqfaIQgWtbHuiMpB/UQaZaqBjAv7/r
1FlvfRaVe0skoSutz+kwzQPjIrUYjybgYRBdzwkQtWSqR5sf0rF/y6X97VxXkUnJBRjFodKHoC3i
3e3n+cAOlyRbImmNg0LXGJmUaOtrarmvSz2EF0PS2yWP7vRmnt7caI7TkjPrHd9JlUKdaJEJPLmI
h2nTZGYZU43w0zUmYvXMo9mUyvT+PrrNZCv8z4k838Ii1okuptc6fx0ByTVy80/y1JxgiE3otnkf
0HvS93EXOYE1D4hhdq9sz/t6kDJULlz1WKLUdg2YrLwiXOzfqmanskaCAMyLIbSlRYf35Z0Hnh7O
pTdIb7BVfADjFc2qNIfRgvlYkD8zoC5GSad3Juu7mkz5dR7FmN4D12Q2JD9TKd6RavwqQ1BkveC5
VUoOtdNBrdQSV1DG+pnmglpvbZTrzVdEIyYO0a91d7vLGeyfD67xmMueYmm3PJbq9cnbKvXAzFlO
fL8A12uAHFijmVw7+3XbjkMxqt2oOhPWMbOQdVfwsFO8HgZQSwDOCRdqlUrnLamKaBVuPPsLfU9k
UTurvgGmNW/DlX3Fsr5EWUjnmZx+jgfIK4JcmhYZeonS/erMFnc7mTvPzHcJqNd53MGq8Z9i/9NC
p1ku3Qsyo163ildFWI7vGx+6LzrXy0F3nOU10JZXzMhc6su1Wwgn5Jzr3u6a1kWgtbZBymi9sA3U
qjAZTNq/oY/os5UXpE7MOn743vF+KZTfGx3hT9G/FexDZuYLvGNJzxDv6ZcHuoHhOc/GYm+v8vRZ
U3NWRc//1iwh+LeoQk3rqdppCdUNJmo+UJNg3Hi0ewzyn9rmUfa0BvRRdmWUpi/Aiz9ek4iCSS8N
WN9sf3qpWBU3UE2JMLjvnP5OdwyDK2jad0ceyHZy6ULEc6Rrs7PycAlvg8ZAhTgR1d3pm/6tvg3Q
EjkdCWnw7T7tIQcx3vLbHeNTv5rb6xDsB1obX/LiYRgE3HUDe+0KhY9HYN02oWmSCp3SpgCGwjAe
yiAd7JgE2UxMnIQq7QCroTfQ8xxgnd4FIl7cvmKo91TidcaRvYDL/TYN/VeWkGKaTlPWi/moY4mT
AEx0hXM9BjV+ibhzsNvL6Ol0izTeFjyc3cf4LObdbgQfCv2M/EJHJRmFfuoGstSEI9JGLSy4otxs
fHeawWUCw2azZMa5lXhW7fH9j8WNyCWbmZyRVJ0U6E0N55+mLJTD5YAt6Y47YMoEXVux+5Wv2PYx
hhiDY0Pg9dST9B6q+FgRQv02UTrpw42sXBtFAGaA4DLTDFsrb+M0S+LFTbVmY0ixEQyY14Q0KP0N
DkhE2i06MGFSAgJC//8RpiiMyhooyvC9z8q/Iivyz0czBAszIl6/iW3iN4ysBeS7tIE8AK6L2wOp
FyrSBNd0NP656RtYEXZZwHsEjapBpe5IQmdwVjbqkCS7F6YRrGXEyeH84lXY6xJDMyBPwPHbUEXb
eDZgfkD9hscc/i1X/WMnwHFlZVhNAqeuFuNH6Jx8Stg8UdrDgIHpBtQ043BMODDIlD+v26+M5u+7
LUtaP3jzfREIQukgen/tZ6SXjCIMruNlq+lErgIo22TPhyJDxPg3ZQtTY54jMNbRxfRJajrPKK32
kdq+P47Sq2AFNhdlpm5sC1EScc3dkHKxo0PBBt5f/APMES/0YMQqdrPdMhAnhzTTrscGOyj4sKJT
3+vpIQm56XuWGFFypuZAm0KuxuG80V+li1ybKyj1cAibPsAYKAPus86fS34T4bqrFrF7lbREprNu
LH4RFEkEi+XSTdOcgT62UjYZerEI75bTYHcCKs+MgVjCkdGhzeD7dlAxKv55g+mxIQk0jRiJhj9f
1y6H/WQ6EBtAzl/sEp1zgewYkxLKuBoJu98pRSvOPBXNYzRXLWPwEw3B9bSoUIzZzIze7nrHSpsW
2xD87p12/y3FMM1+PMyFJgkgmFIwLMaquS8MBW6VmTef9hSTlsKaKdr+eoPa/Nox3ZcHvdf8JsCX
Qa9G+pxY3K/roSoLfDPd63SV32TyV3j02vaf2BZl4GLjTyR9oZuNGoQKlWYQBFRojkMn+bZvTN+d
g2X01bl5MR7AO8fHiRNG1KRjKZ24gPIB0L8RxxkJRPCfGC+0XQ4WQsC7mpu3z6+mj5/MrfQYC+SO
kELjsdK1mg4V/026QUx3sOes+qYEmwMiXjeu0YoezAu+fjDZDefLJpa3Dvf6wM4AEDmlnwX63kwF
OD9pacQ/+cgjX6nkzMwlWfGTrpqbzKJNdHpOCcbS68GAmR2gNtxKW3X71A3aW7LKNQb8gd9VNtSN
/A0lsyI6AdN4TL87MUTgulDthTeqrYjXp8IiQwCqGqOt+l7Ip7f7zpbKv55m0ofqo07dTFuZ20M9
2+NDAEeI7sLF10VaBMD1fnbEBPgPW7k9aKcErbYobAKlNi+rwXUf413k//c3r9UmoY26HW/cKkbU
8Kch8sGYx0s5ZtQHQhSgKCHf39zl9OrkeHRAVTiqLHx/GPVrbUpmtHhF+oqf7bmZfnrCQeZTQx8M
KJOckRLBEqGR1lFEL6cWySj/6+QDU1w1CAGYkfGYOmcjPV11zeDQlrjyFpf0UR+Ci9VciufarVUz
y1P0xVMsFZankoj4mtsWo5C46JUlqC6KDL5HtDIFoGJYNtoec1wCHoecW7tOwhyVCKKQzOru7rWc
IMaElzvj6vM3mk1tjbAk0jyxR4427P9WZI2Ok+O8lyGK6f+al19VCvek2RniIQlaRu/0OtzVY9G1
tQX1bqnSvEbtoADymLTNH5o3xyEPtjiZH35FVntC6SEpaoEYhCVvqbcKAepODq9Vu38Ib5KUqoxY
Spomy7naoNub6jK8YYyP0mTCgkgc7bhspPyJCoprmXJ/1gRpFRHVL68iL1ISam5DrxwVl22ZOPDT
eevLvzSG84NjF7BwwxSXeqxb4Dh47vxAkxLlrpkPsT2l/op/ZriDkHiKZdNlU6q46XgDQVJI65B7
IE5gXNAsg60CgHzSUQD5Y2l5e8g3DR90lViFqj9wOBMuUdi1jNAjpuMryzuCcXDhYclBofFUVHea
aPWXoTeaVKU50zWhPpHiDKH5osPuGDrIftOp4736JNyzxddIqqHNHbEUCkrcipt0klBMW8AHp4Oy
//5GLV5Gxkm5RPQ5M2ewARWwH5QTwOgZQaVNgfpBAbplEv6ua1grmCJD8Y/cUlZ6F30CY1Gj4CNb
1NrEcOraCPUWJ+oFSsRjXh3jMEeS2Uv0rURICL9m7Xw4eGKBQ3+Z3gtewRzDeX2qgbmyOemHmx7H
DQzhJVRyi1GWt9y+fYc+nuBOegt4MSQaSh3vm7Wj9g3xLA0CocSugXHF4+BKLeaG6GyNCzADD3TQ
JqCEm4fDKZNf961bu+6/FXEt7Y9UbLcefyrpkeCBR5UeuHlalyoFk/u3uwm1GRp2D1rpSXF87ghz
bn6SpTFAxO5anTKzWsuymR9Pd6tsdo3cxJXwIVsytBPbuTAyotHloZC2XYnb/4KSVuRu/g83Iy5f
f8QkMnkT/SdKYxdmk8uGICoN+X27jBIaU42OUlt4yIXpthchvDIfn22sfE0V9Gek0izsedqE2Y9n
j9HFDn0gmBCn1Ghf3W5JMoJkDkz8cjazx4dbXCiKhEBMBgDSjykWZsc319FDE0aDr3CEPT9u7RBu
HoTHjJzjQNoc+48T4XSmU2QO79agZfiikrftARQ5wifgaMtHn0Ozz/0h5uCP8LD3YfX0MQjWz5C+
3LEZn+sgYXO6daOjAyoZ472+mMVRcICoXJSiA6j3oGrGxLxnD3XdDNiqiei0GHRw8jEcrLepKMSc
pxrw62nLhIQDX2+fAc7PC9X+xpok2CitGXMB2NCn6UKYoFed9uxB1u7nMCRzlNDlsSjmWflWYdse
gzPGfSz9XisBoD6Xz9BILZywjZ0q7ssJUY4T2O6ih5Sp1ID1J+dJy7RnnRXE9yH1o/YODXpkJZwX
Sr79kTSb9xCslJcCx2uRRQwO20hTgjBqK8X1E69nU5DbeG1wIcyf976ldbHBgchk+B2oZA15nAbt
GaZgu7YYvISHuwPOPfr4M3WrN4UU+SzvSqAHho7RnNZvZqMshGpLDL8wqi31iKvvIzWh9zUbBcLU
cIOGZVG2z2JYBOW6g8FcLcOof5tqnx2RCqr4x/1QV9rGUluVeTKRQR21dqHUnIptMonES4qwFpc2
rguNWnqXKz31OSjNzbg6V08s4f+8AWvO8ncd6l9knwbUTLAFnzn4ZiiapcOP0995nj8XZ2hXo4gv
zjOcbtaaLG1+Gmi9QGt/RqIb2XKKsxgIz3fuUEt6hm4KKoMNgjL7TGy8M7zBoZypTf71SS70XVID
FEvtXi03cKwrV9wqLkUvtbTBMWtWvegipZQ68O939ikTvDRJdIOo8LCE47WPZv6WPv5RbKG+5rYO
Sjc9FYHzPdcRijRKMWBIIE7i2nHKLWozGE7wYoGi2hozANIuy6D2Pix8aC9NtWz3S6+D3Gkc8bIb
rfH5yEB3AzEMLxcVTR/3Q22Kj4ccNoyDpvqcYAkWK6i1cN+CuY5B0q4lX6j0HR2aBWamZITpK/SE
GhSjrp/U7VeYf3VA3XROo6b+lBNdGCYGR+/ScSo+cpCvYiaosj9pr9jkA4n2UCG5E4xZAYEdLjix
sMdeL2r6qbDT6n4sUA1IWnf0qFrkEGKkh3+ZWa9fYakDTnEHBsB9mlprD2qCBYSSfZRPX5gcKhEe
smlvfuCucQ51UYpfnBCEETIiRBvTcn3CRMKS/2ZZiyjn56MVFor5Z1tfdvasy1KBSOqAlm3bS9K3
nPRTMfimJ7mPhX9OpHc9HhlGMkeT+GgZDaNscGC/tztxqlm/y0nQ4T4fB1p/oHTGKyP3BEHxPcFG
wnqKa1lFnpzUJ1ho+71E6kOaxoC+IW7toVwdHUE+mzQimimGQDjxYJRxMm9vPd+CuUvn/Ik3L4HX
OQoBCdp9XklAlDUd5g4/+Vgkqr8KdCHryqX9xT7PnvpcaA1XeBpRBlf0LpF7+hguoy5cLcGfJApz
Xo9NnC1iqw4f8vtp/TkWrOx6R/xmMHKSop1vQfAUgx5KXH+eSKN07bxiK+c8Geseqe0i9eCHlPTT
0yJB1JDS6iZ9vONGSiM/7ytd3+E/Sg0vk+Rpqy8s4/51NGuamErMvfPulZElYER6ZDmmIPbEMNO/
x1c2QnTIu+iYokWyItT09XCX4bYOQPhIXWNPL1rpfGvvsuRq6ffYExx572bAQcfiN13td0dt4F1r
m9EwTcDk5rM91DR50/7bbTLcHFdgv7S4IFLJ98dbAHSGQhkh4if1O8/UOS8l9ew1+9omgaD7g+AL
9gGQf4rMwT9fe8s+n1V22MMVJuxjNiPO+VOw6iA7ZnPR+TRC6k8eHKYXa1CMndVTZAHl7o3WcFSY
Jpz0tTO9GoWWEIrQEU23IVhWxgGMxHn7c3NqxUlT/VWZ6yhHrivyxnAi2gjTiiPpMbfd/QOc5Tz2
zWe6i5EnLjvsKUoVJsv/qRRolFdbPhWwzAz095aY1GmaKg9JPwCveXuE0NMble8V0mt8J1Uzu6hB
j95bTcgQimyeEE+l+tgy2PR+kg+E2w2yv0fFKN4Ksh+i7Dv3hBSeHt5rwb9eFN3+80LLq7hZEBes
cWQ6/Eywcj4P+A86MckR/Ej6ytzK4WjAquFjvBusQ/jyEu8OjCfhcCT2xRzNYuDjCtkRxElQKD3h
09YxJEaCMxndybvVgkTlCTDWjcHuEw5kesRyRFOFkUBXJ9LqQhPciKDPJfKrwTWMoEEAN/v9sFZi
EeVzOfOR1XruQ4v5T8801fm4Jo9qh8NBkLOHh8zBhX2fuGwDh8RNAe9sBPpf3alm7aqnvK8lb9rz
xXqm1ETZ/pJwUdizEGUw/gQnKIo+mduyEKgGD52eIPKhi4OX9vmAGNOH87ah7+gYTYlyjJciNoVR
sEJwu7phemZQyRDmZIIvJMX8gUUOoi+54/xecu8Ts3BPL47M9XuGTsyal46UuTnYnnF8TxF1EtmM
soPHINdrjnjMiUpn1fNx/HF8tag4rEWRdn4GM1ZoZOfWBJiN7fDNOMlnNDvI6lSP1ouleh0nGXXd
gNrCeUeAuAPBNSw1QdadhsbvufidBi/uX/x8wXwQtsiKlZTmt1wzODX2+O6DvLoJWwAZ8mFvC0rR
OtPdwK8Z4sqouT+WxImE0pc7lvlkFx0ZYIyZWtSFLszGflWven+9kj0rz9y9WzbyAF3jNZZoFa60
bdFnwWla80MvTW9caeayjV3pMd7DyPEA9oi7uyl7QbE4dVvKlxcSvDZdlVxV9M1J0srZpu/+0Xl7
uPLNnbVkCD9aX1vzz3hlcQz8EcV4/LkGiU+PczQ5DqsPPkAE1qfp+8wtLtv4FAYlHrpOeK+Hb2/u
RPVUjesgDw6Q9b6i0u1iIppOKD0q4ERsbmvpjbigtyiNXdWDa5F8alX2IYevkgo04DJ5xOFm2yHl
AsH9ZN7NczON+LDtEQZKXYmshYENpZsV6/o/a4jyfmB+3Vdki49F4t2o7a0Oy5ZgMCuaiHbdlVnH
TQjNspe7FOHC611sK8v3tAA/S86Yg8RuqW3NZL1NKXnerf7UmoQE79Bo25DjCK7MlLPhC4Se0n3f
FQQjfh1Moht+UQg5n69kurGYF3D1fSb8STE2kIXmD+8WSYJvVMgkoHxNn/ZDih2UNgsS2ceg4VNG
E3uWCn9nRcEfs+cnnOmIU0/vhnOAkopKX3qwaPeOXDH9sFDCXQ+zwX2FHPuUdCNgrCYYYYnxfr1g
IZ2nndBoUNLIx5jUoUyqICZtOLVGRgBjq7zsu3g2qt/0KWypbT/NZePXDVCxhZ71Aq8ISLx1heu/
klXEZNHTDfWCL+KWUoghGsvPoHMwTzyQrEghjDZalCCEYWDuwdQ55dv9uQs97GUzKOIGPUsF/Kdi
JqsUds8Jrmv3MTHhu8Tx6yjZ/g9bXjbkpfeHqh8hur+jcJpdY2r6Hvev7WQyneIArB090/KfG6JU
RcIvyf8VtKNdl3ClYW9CKbUwnfYnjco3bjvzt4RM6BPFHh/03fl/ZKfK8iQIzn5nkr1zJqrBGlkh
VU5zr4JO4REaVZSbIa7CM6afVKvnSVbF7u0Im6ZAHkjl31d795EIvV+iO4ntIZ5WjwpoXablQOHF
miuDwK5VL9kK2zvt6BfHLKCYhPdrnyRsINGmbI7AvESlWS+qLAz8H2gftSz5aAc9ssZe0l/+ouV8
ImSqG2W0hhvYr3v+WlnBWK2Q8C4AQTqYP+MZgyfdGoGR4qCf3FI77mjDcytbXR3TRTPOn3T2vyOv
CkZKiA6TV5hOWC/wJlR7/Yor64dipD47OBLtwkTbAVHmvqYz9DBNPL5QWZBxkxHPlUv8TPbRQsMb
CSfrU16we+XUhKn80++6k5cfTM1r2vzaNhu7ouZEEVovUD0o9fukEWUMiMcQe765aPus4oB4O4/J
0D7jFBYSZT/MSnGneZCwRJgOPnTYNAkBOVOxqvy8cVetMraTjgoEz59XatMOXqwNwB6GyRKOG9EZ
biQCI9/eXF8lkCknmNao7qQDLUyNo1iwjM6cr2/brrG0GeXJ2lv2TbJHwcLuKdG9r3gZh+M5N4+R
V4LtLqthb5RtfHmTgsg0/s85heDI8mR+BRagaNBiMgh2+E0+EJS0UUodn7r1W12cJV99/jROs8nd
ZJfuEX35EHB3OlH5r9hyNWcuDiwBibuAdDxH0B1PhKj0ZfENwZbK/TAIkMoaV0+0DzA3070Du5JI
fSFHP+DJJdAfg6iit0yrS16TM5AJvfrZ2lE4nQA71jd2JooPPVh3xCeXM7mniAneY/riAB/T9UG+
iNWp7Dtkuo52PY3jcmMs7k8oqt0ckNg8QknN0H2Ax7lcDjOtNbd5PvGihMhHpjQxp1G1WjON8Ckw
XfmpU6HSfnViYiCSz9ch/iNDE2TIKDUPUveNic7CM48idHAeRI15HMp9tRpZGkdn2dgeQvD6LJcw
/7INe5r7s0gPw9UNx/VnfBZRFl5E0613GY18npHWGX+iTD2jO7C18DQ0ASHoSEMMNxMZrt3R7zfZ
pxbNgAlkb+AsTehM8X9NrfkpLCoYbpT7wIkM6jvzZrryK6IQR3VZhDX4+fTBCk/f+RDEcjzggtU4
w15hn9oFFz3MpkImeer/Q13AeIeVsxwdoYs1AmoX6GynN9jPKxx2iROG/o6BT3gKwBzpfgHFP7nX
21n8EvHEYiwgBT6eWCiCvgghz/AAXTsZYl9dxGhAvwnsRxmmOPFrQJnkrjctUjoIQWs8QqwjIkYP
tRegxAhljBHiwNhtAWU+fSzmJQBr5ovrL1HnFGMp0VApXo2p9S3FV2irARPv2YAKVR44BP0LPI41
DDti44spOlHLv2Po8BDmnAPixaAO66IsSbaQKGullTit55090E8saHVyiDMSSmLJliGIB5synmyO
5afURPOppdS1d3yesefzbekaVDwdL/xSR6e6vlkgFanjRGwOU9USjFOLcs65KBODUJ4XpLhLylSW
aIYDGe3lQNlDYlsMd79sqQ1D6Jy95s6a0YA1c6c5bOb4p8PKIFIYWCNZykEMQ5B+dH/CDI4f5fE6
aCV6cvHif2ViJeTTY3Xm41T21oeVKo/WNkW3w6E98z7rvrsvBVV9+lpgRyTwbEyHN5vyMkCzYBy9
5vca+2iIpQ/AGstel3bnS8W602x5Ecn9ODzpF6ot/XijZRp1L69QfCipyhhU9L17uQCuSBHHx+h5
Xlrui9OssOxTX+oyHyvDmH2pCTd5J89ujoBLjepYTQZTZAAVS8ViwzavXFoEelYgC4PKtNdjU0ji
laco6leX64OmuLbPpER+tdXfaBBIvlvs1O3R1occlHb/sr0L4g4dXn/P1SMtDt/GouNPAFWzaXX0
z96Adi8isVZW8WQtpSCZHwt/cidsiBZ8+WaX+H4rWukEnI2ps8RbrcmU6v4KJz/7RCzvEmb5x2ec
mPJ6TzfHTInIEW/Pe0IXDldhY6TbbfsiL3Fn8a1svwJpyWyzGzQuwTi/IyzU7xuEG9jyaDE9dinS
7GdEx/+kaLjpnuKBNTywCHfOL5zBk7Yoo4vI3FefAc8kAl1rdAcGJKUVMMw6FwsXY4oPtm6bvJ+f
cv0U5f4got7Jirl1pJlNpaMosXzLvWexGObBl58Egp5ZyKByZh5e7l02hE0+s6/wRIJIf38Pe3oU
39FRFed8nbjaDYyVVLxeehTHpQlx5pPNT7YPcJUqzFxrCx7VeYJYYZzL6YSQjsgBMzCBIVrSmmxI
clQZ8jn/ecs1SfK3zLj8/uNxMBYvvwfoAbYLwiTxeshAVA/0ZK1RhDnOVUPjwVYZ/aXpgm8MFmwq
3B55xD7Y1t+ftn9cFWKm3ZFv+YoNDYIWfPwxVZKzbnbSeNaQVhgax2V9iJeyiaxjZmcCYIyTyKSj
lpYBxsOIig9ZLN2LvRLC2a8HQs/JqhsRRP2jDz9KbvLunSRdx4aB0wv/C2EcKDMdI6tu+jzzl4H1
5sh8Swm80EcxlI/f5Ea4ugK/PX4/fKMZAz7BQXWCF5SHrlgCk/62aUxCY1LtWediZlrLqQ8OorAp
7D+LdSsgp9GqqUtNibcQJZgt0qWetI3+bTam6YmFuyaZ4zphXFOXAkhzQUYQDo6W/8RpnUo7EM+L
0MK2h0rq/Lid2VcuuIwwDK5HZ1v0VEQAMPSe8anL1FG2NPWFTf46Xx3VcsKoA5jPBQp8EXXk2WFP
dTGRDJoDWepDLpuMuMaS0ikEBexahEsesV2hxE61jPn6QjYlrTV902CP7PO5Tg1bq8gNRAOpvm2c
ryUqeN4CD3xYAHEiMsV5vZRUycTPjWbJSPuw/xfh4LK+FE/Iln9A24FZJG6NIPZ/C+/lJpclLsIr
UwHJnhIT+ryCYSxuO5m2vub9wQgAI4npc0FAr+AQl5tt2ZHfGURc/UoYoeQjyCxbrUyMsUDj/umr
K+vtDFltdxgOQKGjZY1sJbh89xDka0kklcK3yyM4V+e4XZ3stmQ3N0/4NbCmj9nX6KNPbsB2p5Pr
jGBZgyg8N8t3bXvmMW+zYOlcROCltj5yKVZ8sXEgcjETst6C4SSZSvLgnYFXmSdp3fUOMt+4K0By
2JrMEKYl/zoPkUK1dAKcJh7hvG0diCDV9rv/F+OwngVyxDIxin7QaYUtIanas3ztvEjbs9btJBke
WV8GcBSv5D0fx8j7e7+5ld5H+RPX1oVTBA1xUOeRWgc/FQQJmO7JzwMeGoGrMCDFxxz/14osytHN
etEjHISZlRt95A+VHmjHXSAh28WCX/UYltNC1sxZLTPsNVJaScej3ewiEYnZ7MyWDod6k6BXq9xk
kN0BEN/LpJQI3GjUT8ZSSVRC3F9ILzHK3nzlSl77eEIW21s2PVr7pdb/9GtYC0MFwnvY03d8X6Zb
a/J1goT372tmKLzJ4R4E1e9Y3EFh8gg+H89vRH6ydkzfnu8Uaa+NgRdkhLBUa5bIqZpFeyv+Nh8E
SPpB8t8Xr4DgIrOVywqaNojDGhW7HcDMkCSiTR3sojlWbmtqlP6ntNPOtGMLl5Ayqcfzz/fqyTIT
AF/uhMy67kEMlp1PJqUXBLXXjssnweS2ByWRn75B7A0BAAdhW0RN9SdhNoPIlNidCbQR+0xSGNOK
o2G0tP7TM3HxW3V1AS65WNsaXkveSdwV3KoTTbZcxWE03itEuePg/2hRQrCjSrnf6vg42QMFP7na
FyO1r8gmZ7GdwyW8FH3ngbqa5I4O5VDMhbJiFyRxSzX1XjE0lXBnIAqXe8HgOq9qYx7nhr7WXObp
B9W/47QwfaU4v5d7Tn2WOv3QivMzbHYGkGqix8ik6voSQTP9WaPxfo9nSIdkgJMP8EPsh5wiQ8LW
qO+UsgBUU3sKBK0yASdN7jMzFNirsvU1g8E22RMdC7rJ2mDR8IEv1RvOjhE+DVMK355zTz3Qw8r/
xqQAnJK4P7Y/96AXKhnrpgd5TUS+p3Trh+i78ssF8yv53U/1Lm1ThpWwFus+ue2svQ+goFvroXL0
UlYmDHyG3k10duSfHSR5PAERemrxeKtcTxey2JaTH5SxLI9E2eYLEO0zgyKs26mwJF7VCDW8bbN0
YtNbqWCABBHIDkgUHpbWQbaHaHIxrj6Luj9x1daUx7ys9xYHT7sVPQlsYsjxnXt0k+B4B0a0+bmZ
Qk4pezNh7lz7lefVjGFNKIolhlPXq//r/1DSTgKKcH7iBK8Z7es6uO/MqGoqf6155V0BWX73eyMc
Ru3iKXvK8BFYWPZMmhtluWy7MQ/KVKv2zeGmSGTbSH/AWwQrhYs8CJy13HIKJPflSFymWCvZTz0w
ibzZxNqQRba/dzXYAoIl7Mm7drojQHF8x3fEf7tMnkdirCRPQj/0WrMUF8SiKXkjv+H8zs//YjzX
0+/ucp1YnykkdCMv/+0ycoxuJkOeXWpmCgy5AgfNTofmuMGSOTH/cV1kU3549Fc95BtJqsFIsIUg
geES4yhDzasQmZJFMKBbjUJJhENcw5AdzSwvsaqbPMQ94WNfKlj6C1l0q0bJJZpniQ2rCqEb+X+r
jIdJsgtdOj60HznB+uhTk8iHa48teulg713uJnO4Xx1etBmwwWZBZA58fVjWY2e4xDfk27eSrG8x
K012wWXOV675ZyVino24FbjVtnQ9VTongvW0EI1HoHT6IK0+Kff5wuDx5L+uoaf7ilN04UO/jZOb
M/Vw5Mx3jOci+cdQPshaEYt84cy25RoPeUGZG4Yd748dNwCHM2oVVwf00oiKBwu7uY5iPWgdAMnr
GjcSaYXQry6u4vtkg0pe4uxH5tQz3RqjUxuglZgK/RZhAjTHAW9IRjeoydXFXXQj9H+9buJkcGe+
HNpgqFU2f6NsSsMt2oQ9gC3nUvEC+eolc55BLkc2yRpxTpXqTlPMwZPA4wJD6wcTC44n764rKZcJ
ufU1uHy/6i5nmmCQ2mUxfl9JZ3TNbXbUJqJeFAqixe/B7gpfgFOJEE3xMqaU7YQ/UDrT1fXAYH0j
J61ox9wUZ5GVcyS0fKnf61/gyE0+7AA+u7WDCAa6o3HStjL3wQBKsBcvu0yU2V/PUvpb9A3S7Z2b
pQjDARNLhZstCgYmF8ft7Z+8MkKqI7BpoYZfkj+T7kiNNmmZ8imB7a86fW2QznFJ0k31dHlIoeRe
enHCrzx1oKG4HY2UmWmraI73i2B1npklVdy02bo8QcQHc8NiQi5HO9zmuO+rvsa3jORYYhnnsMgz
zmsmhiuZ7+BrMa9KPXX5GwfNCgNjaw+/v3fGV8i/xTEJzdgN9l06/XsHIwdIOcW/7XPYJZLAEcW9
vgKZC04eesj+DrdywsW+hm9FZybZJbcWSEITrpr/SxbHmGmkN51aWINoVhAOcx9ThZ2T1DsgjjwD
k5qXKEDZ2BxCbAYbKIjhz0Mck9bFYKUvVPsVOYjlaBpA0gIsg4Bd7+giD9wk8WNiyqgtravO/kMb
F4uEZZ8l4nCgGupMLwF2yJuMDR+4e/sbIPAPkt0oCyl3PhRknb7HzQzuBIIQaM4HXrY7y0Gmq7cN
WQ30TSphldIYWyqMRqVQEM41PTpzLCyTkmVgNONV3oqjo7AnrgiAkh8aWjqqrgAIrvWL7sb2uYpr
WHMBbpzKRwutm7OO/JghYIuVOg0+qfjo5irzfmcPTON6tkO75yk28fSOYuyxGTHX5Ia9YIOe/HAz
tnTdr10n3RfYKRT73J/dTnN6eKja2RXGqD57O/uFHfl3waP9/nNmZTIWsnYQ/FX1xsMp/Uzhrxm0
iNN/XtpXb9GR6060+w5i414wkrZru2H4NF87vt9YUzG2A9hfdQUO/Jawu0WzVhg/dn4uSYCvzWPc
Ap3NyfmMOcKC+p0sdCB3VdtT6f+EuBgyJ/jpvuSraZlsV7LtNgDM6Vx4G4ZVubfRTmE1KPjhTe5d
aFZ/e7wpNJAFXcmxTg8McGaiXpx6oxFAYD1xVaCUIZZWUz2AtRtyjjzXOQnU2QXDW0OLvA53xe65
J8dBGDXFV5V1E4La1IOfw97YuHkDv6aNWzIs+ORKMlsiP5NoCWOmtbZmx+DKXr2h7tXs7CBWkIEv
s+nblmoDX1971XkgiCAhzbZXc9q7Gl5tML2Vf060lk/0J3WsJW6toNuaOCwsJBYHE1ss9xx43Gct
3fPPdGicBkCDOjcSkZlyk5bXen7FRvUW8lMa9VkBf2h9v2K2j/qpoOZ6yqyqJA3POcxnSG5nPgDQ
PSIylFslwMh+B/yKkkH2XQYHiy6yN4RZCqLa/b+GgGE/8/0Yfyo7Y4LAxwmHTgpcW3Co7UzovADr
7MOIUBRwjJttQoz78acnZda8d3/cZqS6eGYHWfORlUWGYHMbcOjpXrVfIxgLHhLhM7N2TAxcrZLo
y7tq0hqM6DQ+lb6peRTgHF3hq+GLQQLKmHEqK5Ga7GCE+b7iR53nbP1txHgx4CoTR1enDd2+FQSn
XExt19s9YpD3ju331h+HUZYsouKpzH89glKPwXtqOaDjRXtNfE7qOfkYeO4EOPgPZnGKqzwOJEIa
ni7zN/8Qa8kUCE1//bmMRIHUbsPtI8xl8BCg8qA8cWVJgpZiwbJvy79JD1V/klKgEhWLFWA396Bc
RUQweGhiEvUC3i/jHIC1WJ7kYJY/WQlijIjcKZ/a2bI9F/17Htiz19afdaQQzUsKZvUSzdcFAwkR
4i1H2h362raQtOpLDxDFhwiAoa+6BHRJCwbaPA7sFQCjJXj2xZBIBHlevSWvnJUczdN9b1EvlhOS
d8+hU5iTMZHg54rJxs8eG6klK4Q3/dQqXJfFYzlN6piEix47ra8mwSuoYhot/EXxCNMh5canOk12
qHHY9aTu98nNBTpxLKGtADL9fWeLKSLOplsrTfw5z+EtPgtLnl4MUJvWJJ0+1lKxanw5jh5w6Yi+
gxOHzrk9SYmhFAWckLYi9xTIftDP4WPXJQAJuRqimlj00Yq+g1jd56jPaVWfslYGmb9nhZyEPDHL
R3G8njOgQSyzEdUxcB6pv2r875mYqb+TlIPvQUwP/cPpcVF+M63nBdx2wj/WFgxl2jClzcKdYeAE
ekp2P7wtEW4GMxPfjjTqlQo5kM1wuOCrBWFkpXsARPBF2LzGhQ/sQHXTioZZoohvHjt0qdULLRby
UyU6ucDDU5pLRuZTBiattCFrWle2fdB4wGVz1Lzd9370NHc7QSspHzTEZ0iev3OsivFVZZ3BeAXI
RkaqD64p1JsigFUHIba58nz+knyimwr16cROVxx5yo8sJmF+R1+Gua0N80PT5rk93Ym8clhY0tJG
aF+Z5g/H3AfHzkPPXd8UerdljiPRKmvFgbP972kgNS/ZFgh16/h7rnUdWG6Tt5ZICfJPQZAB0YGb
UxPicQNSoz8c6weNLBAtHSH357Yz0YN3YsUqak6Se3kIZofI0hWJCRlBfkRaJBMGPlJKlMCtoJku
wCYVZTM6m6uzovJIp6TE39ssxSSQnFr1yP1U6dhI9AQiIkpoco9+NsbrjiAyXsKfqGyEw6yr1oqp
h+fujPPcZ+Zk/ey3P5LlmQVKBTNGFnnOX10fXPnLvF+intCDlofbRGIALwlQF6BVk5C15PuugV7N
x1M95Yr8BWoLR4vHbkUa4LeExuzH6sv0EzkLu+KcbJGd9DHPoYZGVbN+maSw0l6dnq0zFYx4u7DS
R+zD0RGJZ05phIamPdXnrxxRSizzwM/J2mkxkLI6XNMsxFyahngTRGnVrp9t2mbYKWHxkXWAUviQ
P+IVTOOQXZEvqhxSkF9i3sTdDCBmA+yU/NS8jwJUgagWPBZwrE/iVwOEs/pV/fc+NCF3wQMHcn33
OGotmNPQ7DClf3pvce/W2/1HC7TmBUApY2VabUYviigtdT5OyxHaoaiwsKpZxbRPndG1q335Bb4h
4ChE7YxgcJjswFQHYezI+WlZuODqKv5T7Hz+GKehMFWb3BKisXMUP/N2OSZAUSt9JLvf5RWgYh+T
E39cRueqUZBFQ76+iWmJax0mbQ5OSEmPPDHmUt76gt3wjYgWWJPblQ5Mh1R4qyvR9cFZ1Xhk/1s5
qIuwTLkwYGA2KQKDMCmuwbA9LtBAp9WJ+ePqTq4iCzHXA/oXASHpfkY9Ker8Id/v9PTDfjKrQJMk
RRDi/S/cT1W4WSU8Ud/ep7Dh8Xo4zuNDTLq7vVrWNL5DS2MgQJfD4cnCxQdGJynCY2ibUIGxb40j
oDhvodNs6a/Fs4Y/6Fbv3y5A3bmCjc2q0UoAFfz0Vv4qLELC6uapnjP7m9sVuD3aClAcMboNq08m
95vPuKruYe1zFE7u1U4s3fkc0BAN4lPx/6WL8dNCb9RKGjP0G4AUR7mKo52WeXHuyyMnx4549ssh
K6ZUv/LqZGIjs4GIKLAc1pwWBMNqOiIYKT/LOCHUHJT5BRbk2sClPnQVZiiXle1ZpqvAVOHxKMD7
bhwten4xr/KUVnbIkLf/j3WcXRqMUbLwLWqxeblspeYqT8AzOSfAgXYSAQiQGrtoo9oVsvUYTSpi
waFRvOVkhbfF5KccP6ZUvjJs6TX9E+kL0KTLURuF8aY1g8tB1vR/jxXYosEYBcprPlmRoNZv5Kur
kT4suOga4MtKQdAROhAQrTc/aDXS+xweOiFgnj/8F7i3QSDadd/3ChzggoAoiH83A7+AqrwVdSIq
lM2+fc+pfAtNwrfZe+rKFg/RN0eIxS1Qoc819dknrBceqA9QiMj0SVACcH6idkSM5m8Bfx798h3c
EDUb6vblgzSGzRHxWuWBNgTOQJ3YJraguwogog+LbTPxxyE+S3D9WAm5GunPy0yECIzsLLlyEVkJ
OLJoY6ykw1WeU28pA1Fsl1XdvLGJgEZ1k8mbRId6rUW5h+KQsOdto9Rm0znorbU1y0KGM00x2f19
ehSKo7EPNqfJxdaxTM9zeHlBQbtYAzaPYLfzq/zvqFmddRoNYoClVHULXHD62zW0B2iHGbMpwSIl
2VHM9WkTcXZ9iBmTTrx8TdOtEyYGg1IGvbFQhxBoVTbmyhcxTN/x8Hk/FEN49l9cOIcpsxOJHlsp
uuEi6VQBnNNgHD+IfvpbfjV2fFAytO8Mp2fIa4OFEXqmpVc4tevvNIgVjV1sZczLxfiGX4tsL4PU
PZHLOEl2lOwsbjpm525FEU81jRBmSAC8y1xUAzqMZESaH7dxXGWGXwn2Gmw0C36XbMKGm82JBLZ7
p8YznGfKYWZrA3rmEMwbcHczMjPNorAW/46dZRd5eohYAsEI/yCkPjdgmW7TWqLa4ZHYGDDlFaNx
64f9iGUxIcCmcZ8S+66ae9jddHzAOHz7692NntBDdd1FnDwTqXF58jcUCUq6Mo3d1nTqy3gNJxg6
1K/A/8Jz2c6IQOc8sR0QXyTPcZi6i06zV0V60E2fjGJYBVMUMvejNACw5PbxonfcSiPjhHD0IAVC
mNPed+GHYEmi6/tsrNSfmZfRcKggLSQf7dCrClHeAEBYyZ1hOeRcz0echQLL4LDQwdv8Qk1HuIXX
RwpTCvd1TP+5YKsFXCX00dNQqCLctbFGetHMsZ7IPdoqsxxlU3TeVJYAW8SApqVDC1tgLjq1PJKg
98lVV0Am9c/SXGoRzfw0sBucJzbcbArMi7OlMEB1yZ4jNVx4vLE/+X444PhYiXh7en0TYwL2FaSD
BCwOMpUb3wtamN9kg6IWqXa/we5zQBaIRFDvCoKpuCQORsor/glw5mK+zwiUPsm0jIJFMZB4MbQX
6dAcB2Y89K/EpHmnH3bALYCZkn7V1PlRPosUzma2RpK9v6hMRykvGj9+MHFToVXVp3dzkck19SLj
7gmEsKCI2qrMG8Q2FGtthq6GRav1NuEC5i67HaLpEbnXCCLhMD3OdVY6Q6Qkefc2/ME8Xm2mF+Vs
WvsRzBdhd/EzSXl/fxzOM5VTZuWvs4T0ri2eHxz5tovn3EqMGuplUqbqh5oUj1LBHjsJbU444qtR
T/uloREZkiZBjSBnjpqxm8pmXlsgmOy68ranq6psRW+hEsWX+E9zYX374jXCBNCN0Sj2syA6exVA
+HCDmdvHr3ztLAZCo7ISZO/i4PeGgq+DmVHYnnnHHX4IPEMZ3OXck3Eg6o4W+CSYr87yeM+iaOlo
zRX0dGhKMj6UpuCZXTTV73kBfaBJBh3ZsZ7r1xC5NUcIBXBmFu7rP5nB+kJW1QsrobxJ0U7UhphB
yti621uIjaPCKOTYLWWDN7C9OryxnywVq7bKE2ArigG/s4fjRzcT0CcvLvxa7L3CHCNdhMhGtR1M
NnRVUpiBwWIDbSUncpsp3cgos5OZzLxBnbNSlrY2d6C2wEI6mVyZTwcPYUW095NL6SqQ3epcs1ct
IQDxc36JL1oJL0g6sxpQ5DGvWeDQGsNtADZmV1bcXcrpAmAJnJ8iDl4AueTq4cKUkf99zYpq5X3A
s0EcY7Q7bNLqbQxBHN8DBthWobflQTClNK8TW4AvRd3gu5DqnA3GQ7Fyh+GVTCxoLwqlbSp4P/eT
dtfnR+r1GEcxqNm6vHDRbl/kMc3HX/r/EvGyoVAkH30vsEYASoVUV8uTVcQEAQAKCVLgB9Oc7c9A
xW001BGSUixno5gjiwKuus1bxzWiYhzRzUFkoRvYnHh2XQcXnuHpAUxm+WDp5i4SU61N4/YkwV/S
SDS0B5k+yCPrcezcGkDxt6haqrY5N7J5Ec+ec/521yYSBZ+a3oc+2aBjHUNJ3PLhK8wQ7IDGUlun
iMo0CuDT3mXknrogb0P29DLZ29fsWbZR2E/jqy5qe0e6SfYwZiNEYp7QIuWSeRjQvgW6GnBBx1xk
eGLdvdSLwUbcKHJRJuCnpAINNJ9DalXFNhoLl3zW8yDVXWu+MUO5bTu5xRH3NzPgJTC/X/fAqyv+
m7lWVygXW8xaaIJgZ3UZPIhmkggmW20CWxNIGkJn0yBeY3SwB+NktLazl8Ol3y2wfGMOgeOjeXNm
dmljxAIBRPhlfSjiLT7Vmamqvcr4OK5vX4u9tcT0MEA+iaxQlzIUELSjcZ0Gf8/HPcsX/kPYOevB
iTgm9LS71tlFnx0E8BrK6Xm2tYwIuslXbc9N8+3KS0R8YcvUTcznpVEhTX5fgSiKt2rZ3J/FwDYW
ETwzzW0SPhwvsgvmQnI+6cjqD74vOOeu9m8/Tfm1LUepCT7Qhadvvdo8wdeN8QwkVg+A0EsQr0Hg
Cgh1airIpwO3aKGSk9Uh7gWwR78evHVXNpXZdcu8lqWQVPukhejW4yoS6oE5OoIVMtFlJQrxEEUC
tXI/jwgXex0nlTm4d0r9zahsK3nc/FhmIpkcsWlFI8CJKr1nmHR2cXAalj3+jYpyJIGHgkTgY9T+
XcVNbCHjd8/dk7JVeGYHVSUw0K7uBlMsr1OSsVi9+R0jrfVOKbtfK8RsHS4DYMSO9InrufxdC00I
y7tdfEkgigHVfm/ypMJ5fP4FqJuHJHc2iHQtU91xjT/BVjhKqP21jIXOZh2085zkn3r6BgfDfUaK
TYfMNkL3n0ggf82jseA7kZ1f5ihBciBXKVLjryjr/guxvDiBwMoq9Kt8blF+AbhTZQ3wC7i7nl/a
NXlUoRdQrJ4BVRZ1t/fc7v1jIL+juW8cqPzCyodKvnjIuS/xhxwhiTscQirjNUaEcbUvo6zu/IxD
JlexcGaK9nJ3Q+qCGshfGhH5klUhwQy52layvorBXvLpYuRYZuf9s2a56Kuc7BzaAfxngsCwOuWG
nlqA2tZNm4CLVJ0tikFOTS1pcK8Z+48oniAgFgiaMkLyse8iJJNQwlV89vD0Q0Ve7/z9FwG2waCY
lC+8vQ9pfwJeuIetxcb9xlrhrb4nitGKr5nio8t2prtR3uGerFyCJKNgT3A8vmUBdULU16bHbiz5
oyszudKYFgft3W7tzavfciZO7qRoghhP0lKLcoDASUrcGPLj9tJvG9X4T/BK1DjSptt52XmV4h93
Rs7W8BBkUbO/5hsj8RY6VFr06HiZeRy7NergzR61KIQiPy4HHxSKDwVpBvRdKeBhsjnhxE0AE7qn
mIQLRAOqNhF6XydqTpKTl1kdBsxfgscnom35RJ+c9jfoToLCtWU7ZcLEsBnT8MLv/A8TU9LNaDEw
KOm27lkm63mlB+zOrzRBQ/SqKHkpwK0jHmB/csM5QnEXGjBThNCnEuxIvhpgmWG74xmnQRFMLAFw
Py2FGqOGxS7Orklm0DiBAkRJ5Rax7LAMCdKMYFcG/BeeJGKX3HnAnh75EgGrFtnXKD7aqBDJnKan
q99mGDBYe/LJomNbz5WueWxq0AIJYNqMV3iKGBzcI7UKNlUu6Ql3Ah7cwbdogO04vYf+L/5bU3B8
RPnTqV65m/FSZ8ugsA8Ps4mTc+S0doOhFCFq0kZLRM66/FKmyWziak3IszxKIMW0G5g/tikgGio1
8X0EWmTdzEDv3sRqtUy3VBfdfzVvr76k4P+t2LAb+UQ9LkpoeCEqbqyLXe9Oulu1C6qqhGO/bSj7
KXy1Y+l1U79gUma90kQ2hajQyNInNLImCFMsw7MabNQUNoWpnDA6m7gyHU4LclW2/xiVYQKQrejd
gHzqC845957VV62+d7tMVOFe39tL2PArKNSEb5GRxtZSX8WlZDyEQxqq76yRNRlpq6gOKGMLZCpb
+m2fN47+JJ4wNvbSDyTr1FxWs+CTBdjyE5mC3Xu0wYT6xf2gEfhMZg8Z2u3jkPftR3gh82M6r1Ov
bUbPtXhxVNI1CMb5ONHF8+GIcSrDFPPiYJqiF7h6vVAyOatTEfkmVJIW6fEyucLlBetFUJ/pqsas
lKQtVwo8Vi4rWfLwMFpcDsV6D2M7ZrDoniLzXhqS412RHgXWJQKMRl2qzEurWDwixu65BrflGKhv
oCNC+YfAeqlWJyi4g83DIfvMTpQxdIj/7+Xskql7WRGneLMh1sPtG8f0mOw4VPObDsb31ecRx/vQ
vOsgdpMW6h5bd+6td4B8mDtsxD49+nLAtVDNPBn7lPlS2BTwHSOk6P+1xOrYkpTcHysELaOUO+Bo
YLIq2oPXDcrgn3m24yqDMcBp2SkT/hsE38X7LLBaCEFqNHJhcfVXFnuPMFHSpXJcPtF15tyco8e/
eLbnISSYPrycwZlYqkJjuq6gt3QfEIh0jSpxLQpAW1gJOuBjW5NHpAv5KYEyRrT/lA8U99qX8BeU
Tg3crwRnrZcgdG7sGSxkwW6RtYVhkohp3t/0/opE9JMgG+XMQVp6Em8QFfI0vHz7RJ6GmMxfqaOm
6zhauHr6LwZJ9ejvoKHQler2fUy8HUwTMfhPEz9jZbzagt9bhXKu8KHDRqJ6O3refZ8+Cv50Fi/3
UCt5LgdPySbQZYyE0AFQlq+ZYknxRTlJtBshf50Xacu5yu0D0yu1TMCoQmnqmhACpi1qI63x1a3F
mtE3gJxzkxykhUcMy/08hrvaCuPx4YcaaQJTIX2KvhAiwAByzkaedWnXxd62cp9Yk6+VtQP4c/JU
g7kPJN4ob9JpoEUukpEwGVIEkWEGsP6R4sLvmldxEGXVV3u9IpeQILExrury7pRUgGJkYo2saVVq
/+zsRkDLqUHnbjhiqRnYJTr4pqaEwnlKEJxgtzO6eCS0bGnmRtZhFfxnl53FF6fab65UvTfBj5AV
yfmi+6GZY7w3oiP1HUmnB9Kq8pzBQpNLBUZS2Td3G5zLIc8+TrZxZ3Jy8M55LAUp+bSVk/n6wg6j
g/BO6d1niwpXyhlRVJ7VpkOUhH7ASS4bncwNVLJ6SuS9GucRYtpdH7ZMcxDDQbpizoZgwl2noV9B
BSg2s51CFAvee5ZWIx7guKSnbSxesp1m7Vp8wp6ZLzMnVAAmf719FtOICfc2LQrkZL6k9AJtAYvP
hjwjMP3wcibA3eYzcL42nrkC78szGs+sGq1UEmU91BKzTsOiTf3U7vt2uxTiZnzQRiMoOuj8sJH6
mQu0ygz68rl75nak/pmux0mDJ3E8/HDzP/SwMMR3inMvLC2A3G+OZoUSzT90oljt8WMryDFd+SrV
dEHHusvd8OUWNoputwt0WcHS7jXbNSvkkwuwXiYWAF5AuO/snEPDlhoZrGxH0/gWriCLDLMxq37v
94lC9z7Lz8Z65wpC8Y2902N7JqOOFDuCPFhdEvLpskQmoP3cPYjxRkYmytxYRPFszXgKBsJ41gTm
SnTrb2WfyG+BXXqbuO+02am50QbHDKLGOQxbMm4D0fFv2C8tBvVYzlQo1F3hguyr578OXb/5JHGL
PIvNvCh2MRSaojoFEshQlo1KVJcPEiM9qCVL6oeciafCKEJ/Gc4Q4TmhlUC36iXhxeGoXClpaSIb
jVjy878ULrS3apyn0r8mNOHPJHX7TLn0k5l2+pJwz3v18VKMUiti2ZKLfJNJ6BNnFJ2o1IqdELJN
FWrEsFH8tkNszkPjSQncTt3BFPlTQ+QiRVn4YsuzGEHe4zpt0Kq/GwZxJswJpkZZfRYhv8+Zn5C3
wFDY6kgFAcggwPrFuEf0hhsZ8hZ50bLT538Wl1nyUCbjZcgROXPyhMfTGl75Q/Hih7tbgjuJitmy
O5FX7eHuM1d6haZ9/ralved+J5zAEXUMcfLjTSzGsVJcBo+21WNlsD1YcfGd09S/nzyVsT/tJYrK
SPffHJiGSwl/vUz9Qnq8QuCoJppEmNj+dChceeDzivfv+7kC6B+MHuFwKFWeUGCEOU/qcVY4vIW3
YDnb2lvmbv8HyHfdObfT/SZbsb9CUDVgN3CrAKSqhv5sW+I7Ndj9uSMdDLbIAat+naAzNmBdxW1z
sSNm+75z8FVSsHr5gVqxroIm36G84htAtUmFLBkqi/rC9+YoST+otUOpCWK5uvmUnOLr5dfyoquO
O+wrjyOMApC1suFXZpyN8x62vCVbgOK4g9uk79RjYtEUgzkDx3XhPsZvkvQ0hYkoIyjgxO24KArM
n7zvWNrlNuBW8GkUlZ1ufOTjx2gGwZP41EtVjPI6F0HNDTs38Co8/rEJ4ycJudS1rNvssAUsom4k
Kz7uyS2p+aQtEcoHdSYK3mkagd4+obceP8OG8exLTxElf5CfjTn8bSaT1TclE82U3I84OyYcMgpZ
ESlgXa8GFbnjm/bC4tFGsRBMMRM543swtsCnMzW5s+gfSUvaJvoXXIjtJXv2NMjVlZhb9XNTIuif
vJ+DwbQQfJ4rt4HU0VdoyQEpNMo6OCue3mhwvGxqDbleg3kYUaFKp4NIbtIFaCn/4dFC+bA/dPM4
2oLM4VA874mEn1piIiMjVqmjQ4g3Okjd26fWgmgm8LxjIgpOif97g3+LqPbM1SorHQNQNy7IqJJk
30G5pEJGSShmlmuKdGlv0Zr97OoLU8R/aNdTvQB5dceVN9ID2Cr7OLOI347op1CDyysfY9HGWFeZ
5nS/3soS90dVI4riFS5e2FYMFUYC8QzDGsIgTLKL/UM88WWMI7DtFlZkvfQZDkXWkjnQMhFKpedL
14QQvPUJbcb+kw659cnchzYqL6kl9sdPlpnebJ2UWwkDKvf0aplYlHyYnNHh9moo8FSuYQVjvpbw
dlBKHCchsOvXPn2XNuMRlncaS4NHwVxJ29RVGVhx/xwyN4+n6oOJNEPRyEKD6t8fFB95uG8NufPH
Pq4i1ieAp2BfbUNZ8swNYRqpm4cKqTjcxdYV3g0H9kYbvRpVL2b/j7jr+g/SJw4aJhY11SNMWVMm
Zz+9ohUKwlu5qn0jbeh9uy1Q4C3H/jbmTeKFrP/QsPp8+mMKFx7Fp0e9wRaXDL0Bh09TIAECpYNM
5MoX2muz7ILY7ET6NEYmQ65g9CUyZBakD4zQm7SAu9zrJQsSh0cndOjLzfUKFhphy4LTT0O1XtP6
C7YrFfdF1BTfWeEOem2mhxnXDAaiqJIy7F9lUBERdmRON0RdRP4CygFE8LBF771uY/K6MSQ8Ufj+
M14k0WK+61IrBs0dWP3iUaiVR2VeoMAKrs/C+ikDXD/HWvFSyI30gn8sLjlCT3MEZDIF5u63HYvE
yX7BAG02scgwY7X7YP0RWX/orM/0Q9Btf+of1v/omXazy04o2XU9J3SK3UTXYbVIhfGCOwM1L0u8
mSlW7+/lL0dke452JtdHATP0KLK+U7oI41DAYGsqAyc4pSjTTfku+xttGsCuF8oeQmgZ7Xp60z0c
f+Bh3a8srCNGJE9VH7+UpmAcx9gh3eQTO5wop5J5+N3mE85hHRRq5Vxq1lfKUwxQHfp221BXTalw
WBanNSxW24Hi97IRre9ZhsPddZtJEqs+H5RogrcyqGyQpnF/Gu9AlMvhnRGaQermot5jQEIZikIa
/QsNyIGoc5Yr3z3B2RcQFv4NWLNeU5OUG91MiKYWa9P97JYiijAp304qO5VpONVNnVkstToyZbGr
v/JisIayeAbhEO78vRDJfvqI0Gz/Nh9DCSFCRuwyvS0Pho/zt9x3FETGmdT3z7lCwATnScvi018S
wmRf3X1HGkyEMj92b5/k+Tz50R2+h3khbv7/t1gOXW9bvcgW1J2pzFX2bbBvoVxbasL+lPP7+Xtw
DBCKtMNHCsC8kSwgAqNZO1OJU/8al5Q1Kbs8svmT8w3n4Ks4KYfh7X0E0dhlwOpu0XZTLVHN/m3Y
WJPRZS5DvGOnDOBYzIDu9kZ7e/KnMDrb4v2YyYDwFEmzimgv0OgW+OrbZ+9Fzdir76sLK9XQTZvn
Gq1/gB9BZgy+qqkH6/G2E6kpW31ByMbh8fGOWdmJ3hEbEtlDD4vfDZPFpJJ7ha86uk4PmL4b1Q0Y
IA2imBSKd9+1H11qiFKtKIdLHySCbX5kBryauRSVyf4adDt6ng+bEuD11ZOHFndi79HRWWr+fD4s
90FFeXfZw440/YQzJbjdOy4lpdYqiS9DYrK/iIHsvVh4EC62Zv3SoZKo0/84OiYm1+8IBQA6KM/f
j3+1opCjWp+YuvVnsj4/d327Bjeko+GEQ/8xzYNpXgroWQfupIhMraF1jOyw5ylaj+HyUmyswVPc
9raOa3iW9g7SQMMQfJv4tWGtm64v6DaJCPCyaf84gVsIvMdSXd67/sDBp75mGZsJ0gT4P/pSQ8AG
O3v0SiYOqQYu3SzBIPC+xuSei2g1qa7fGqYnxYQ7bNFPOrhjozSYeRFpTdZsbQvy+9MANHp8XSei
BRziFxqxd1+f+R9CJ9fqtfWuFcwSHw5//M+zGb9gbddAU0K+P1SrQl3Mr5es0rpiu2/sWG0iL7k8
0Nhgx8DQwHy+30GO2u/obJmoCze7/9fRTwgu7xunOKm8Xd7jBoLhfvVC6fz/lqHC4SEhwUpWo9O2
3NEOdpjVhGR4YaF9ypedCHiF8V2sWLDqfqBTN3RR+J5hjNRY1kLbT0Q6cJUy702jKUPXi0ayQWzz
cVMV8p/pQBLyaiDb3GWk/ME8twoapqKxnMczHTMSCxeQcv46E1ZQigtmt+q7YpY0/jNBTDzbSC3U
dhUKIGowfsKDiRgAok6+CitzDrFNfXox4zSNNBSBYpionvImPg7gfS9jQpPDN1TvCbgBTfxoq81g
QEewLdqmpBoXM90CmFp/sU8ac8QhJkKu/pfuBjFo3T9knFG1T7Cl9zPbuh1fQqboMHuAbobtJQu/
+YhggwxKpZuFnxHq/vPMQp3s++eWT5ni8kk7NL/4XMxZApS/pgjISHg4wSiO0Lsvomje+tqeeKN0
E/3LxBqLPYflLmghL7+iS213P1dIAt0/Id2xc1XRcWxDrYQU0WFZKwS8Q51z0YhlBX2/YF/psagk
w/x/hxlrxFCF1YKHMtKkoWK1lnMp6AcF4Fv0Z3lifTihG5AH5sItDBM7EWZaHT4tD1NP3Bh/QsLp
wWjdEfNKU5tPP7wK6FpLWEtyX39hwCLPAT2qsO7JOj6w/utJCAvkRYOjc1D3Dfe6P/75BEZUCEDW
QmpJycCXOklvCFGlN2UJpkq9UMvnn2aJulZdhWUSICRTBmZqJMlSj/msUuIfOu/8aU7fhCLBTps1
H4OO2ofunMWLtR+s2t0Eo+M9QIGmZ86L3sC9vLVN9cwVrgVGlG6xmFTk+BwxaiGsdLF40PlqLjgu
PxaFnkSY9DpjNxZduyLCXDGLo2swT1SvD9YRYzqvvApnYpP6RoM6v10OSV4rdguDoU60Yn26c08S
fsaAFDIh9uYdnopeCIuwtGRIlcT8/bgN8ly8UdPu2RUnN2dXfWx+ZnOKK6iaGxzYsMh+qo7HWXkA
XWnG11wIK8HyG0MLHlYjuZXE60xDz3P/KSCcY4McAFidAR9jtZ7YdIMcx6HxV84/OOx3Fadw9IAM
WqT42AkfRd1rAr4SDqWKMn3GC1MYk05jsoC/Cn374Z1GL3JM1/X6PphAEFF6gcyDBgmIakAjWS45
KZa0qMki9hmc3+DQ09lq70fZCgdp2SDWBgljXZJ2rkIA6fR5yDOIK9CgP3V+E6NilpmA6SEdKD0o
9xndwCEHSRxrDyfv/GsQx6H6MuYZfe/N0d9K/k3ObfFomKXxFxwj4nJaN1Xy5CZzRLxAtJKBcxEW
EMmzeFGveXov8hZCzT5cOm0JGMFLZFCZe/gyHXH1ywUo2k9ZlGkWpe204l1FuHn6GdKjXT5Ven8o
Wr5OHH/gGOmJmDeFDMBr27zSswQsM2Tuo+6OruyHfQ8uYl9mWtQtYFYF19iz1/3bnV3863Vhm88K
Ytor2rSRvUya749yOOum6iUH5dbR99GIgGg/k6RpKqXNUz+q1zhU6wnk0Vbfd5Ju2WdfHfu/Ft/K
0HXWb1gp1k7gAoK/OKX9lL1pN8Bo2tVzXOIayrJRWp1IAgXIkQbDSZDW2C2Gm4XqKfdpqrJfZ5rx
yFWoszt4Tn8X0A9bNb6GCgC1YD7mRZCsoy4hGzVaBEu52MVXwy0bi3B/MKcorG5DDCaFZoK9Uty3
NQ2YloQKo0HU+5u4lwjZj24sealFa+jOZH6NlzCUYN5NUPBxxtbI+lpMdqVP7WhIeMl/SrMb82oS
dS2U7vVJf8lHxnzy/4N+SAMBs53UhwL/a7iVp30/OHe3iEmZZTheUMSMk5Tx2mzU+1dTaxApZfQ+
5jCsHNxVA93qKBv24D6ZFQr3xbIVdTw85CWf6CiDpZ6mA6R8GNgOmUctbiWkqw88u1Ul52F5UTdN
0cn5lHxfjmGAvcsC670KcH0s3HTZVi4ST5iGL5Fa1DE0naruMhsl5N+4Bwd/OzrPPwKJ7B6pOGoj
oEoiWRM5sX8bWlYkHp7BYt4qqvw4vYCKc6roLW7KAPPpW3j/JfB7v0LBjVOytKvTHs3BU4EgzUBt
vD4NoHyEsxdkaPCKk9go0y27Xddf7S5STISL+uOxKFm2yxxUev3mkY1PEWM2a/D1MER9qE7SmYaS
VmNjrXbn/0g6L62+NXW2I1WhV/Pp9Irv7pH/HGDJlg/MCax2GROqwgTJi+hn86XgV7kkbzNYiNpZ
tV5/pSHZjxdnT7EzHFo+KYkMkJKJN1ykidsE85ABIV1tHHKcP/C5KsCcrn/BXdfC2Uc11iYfupFi
9+muFFqcXPDg0HC8CUssHI9N72vYlwSMZun9Wq2HLQ6CjzIbg9j9u7wUm567QTbRSzK3KDmY67kF
3OqhKnPMolqKVA0IPhqIroJVSzmFdmL1ahzXtuzF7Bheo2ctmsjUCuLRLUzi2wCNZVTtkRwbMZwV
iv+ovGqt02+nA7HR01Xu028977Ayd15UoT5L/NoUx6RrZc9X8G/TOEKdLcRrIuNMQiEBIGCbSAtT
OI+YP97BvR5SsEto0cP70UVKzbqReUsk/eo4fg5hvYducZ8qzQVJZci2tOG51MUGCZpjwbQCi7dl
7UULeQslAbXJ3i1D4koB6/nQ9tZEZTcE8o0Ie+m2gGumUokWRPE2nT+TdxPFdFX/WJzFEAT8MXeM
/fTLYarQSiMLKRecCNkOtgXCQZfHpb/X5kSJjSuXBevk/b3kRpzbzMhDjq2eTD8EJ1b9r6i0hpM7
59W/7oCX+5xBfaq9NR94qxfTRMjoFQhUSW0t698MR44NGZyeMeCD2DjFxeooDWj0q7iNp2gwDU19
1TgdbIpGyKX6sRf8GvZeWA88O5kxsSHGARqCXH6tGP4Tobu5GtRouwYXJsKzp0b94ZtaQW/2JliA
XwILlEV2P/WUEBXeulbpR6tA8U6GUqO17qvfiR8AHYjPWUqxAkHr52OsAyPf1442ZLIX0Ti98RJk
Pv/XNDNOlWrRqwEjNoZkruX2vkDnxYni69d0mPDNFhxAS+qKre1hcI1hRRxpo9HrAtPnCu+nB3z6
//1dU+670GrCQUXOFEI6j67TQEgK9BLrQKuFDEZYHKMJZiLHXK6+fPzRkE+9zWdoy4DpFkF+FqCS
12kO/K21F3lijSF4VkTZiaOVH5bXadD+gA4gUc3mGQo6BN3hNIGVzLJuxC+vyLGYApAXqM0KXZuz
YE/YFJYsJDNd4kor+xCP9DX8SlX8+mMREi1Bg50AjrtH5DA7GH7BN80idrQjdqzRW8itTrDqvamx
dg/07iomQv6XfSpjwA5CFQwASSfGqFtMX0KMgGX4xi/VqgCOep1pb6e66fYMl0fJfwnAhKOsVn33
L1FqcJqKgpTiTe6kEQRQuVjsI2AKQxTjWkyW0OEZvk+Sw6OmTJ25yEyMe6cWodK65JpB+WzUnQIi
sAhWL8DmCcVX9Bfcd5lKVqfH7J7T6QSLbhJLScYg6Zj71hhZnup1Cu58S7yL+y6fxLoOJFiZqx0k
9+HDCu+7jxTS2qmSa0yO23JcGCetEY8huQ2tYhXmRAvhshG1p70ivBBQ1EIFRCnjGsQ5QcfqvR4p
zLhHp2B8B3Sn/A+C7mrjnUeLCp0BkKa6rHIwZL+PhbXR6zFtfPdluouwu1YGXkW+4Z+AMAKBa0So
C4R/7cQTC+y8j/SEdzZ2+9Qw2AqkR30ROoMLpv9U+bfO3FsM1OQghLomlsMuKm7spa/OZocY8vMH
SAH/POKK9KhE/3AriKTmyOn/9lGYJmSc5u4XCPRZ3gGE0yzJNrwNAd6FkbYkbPjY/Y7eBzOhaowU
b4HPZynfWH/5ztxE3EyQNAS50USmOo0OcJgUhLenHPwqKQotmqp69mY13FGGUVtb1bc6GQOO4TQf
mKJwyUNdZZsF397Jp/zptmNEsDHaKpQhw31Ng9H5QFXUjcckm+TIcuYkd87VV5pTpSTMrL4bz7jA
JCPqIBdhTkBxdtawotu5w2wGIF9KKuvHWZCdt5jEeJFuCEClcz93PIVe+VqrtIE5io1vPaRRJ+d3
JtusSv1ZfBs/3+6hG+Dq71RCooUR6olZ6wa8/To3+f5kPapGTwcexODxF2aGg6lSXGaBckLNPJs0
0QcR5lSGIGqXzPHgC3SSiq30nlPtJ73PKDwqjNIIIQOpbYA3jGCaItusqMGcGTVv6MJRbkC1mf+i
qZkrOYrmwHso+PJBOuhAbj2Vxl7ZQ2q/Z995XVnGsW1mgQ/W0p/S2BCie6vYrYLUY/96DAZwAc9d
+TBb1Z6LM45Wr/wxFbOtJ9uFsGIchcqTp9i7vvCQ6MAqEG+PljL5bLFvd8lpZjZtSTZuPG+s6ptm
QKIYhS2B2ly2GVHuP7rgp1KoUQ19sp5oBvt9Kc+M14fN+zm7NkCMf8+wrM/xLOR75S1fHCJSdCeq
KHNmkcD4gq9ulx5QW03IauoGi7wxZB/c1MZb5cCWBc+1XrOAVor7xmk/469bRg8LRgpXxL5jvT9b
H7wO4qG/7ezLr5RMu/A49gAyWjQTFtZ5uuoMNJOUXbJfWMIgitqU2AtdZzWwEDjlvVGm4i50Qo5P
WQYc5p65oKCkY1XkVs5fFLfUpfuHGj3qBkK8KvzplPHJ9MHGfF+/6fUFwfQL4SnofQtobvNG7uSQ
dOVsPMy0rZxoD9gGMkNNeBTGC4+bzO2v62cOVKuLJSC3Urv23zCCyz7UNHIqTy5anKFLtgVZkOs/
z95IoJd5UWstRP3Mzn3R+1jSl+2fknCXNInLX5KMwiy+mnMvfO9CarRbxLEH/U8gZcMochOya28/
axyW0x7TNjDJG31acBgS0IFYyhItLs4k0A4ixLC46/TO1TKFHXzcQWuEQB9a6axbVRxMxgb7knzy
yLiEkxd7Y93fBbDwoFANrab6ElUfb1iD1n9n7xeDWhqgeds1jUaEZz0piOKRpk3BjSJDaOhlwv+j
RPY9M5bz6OQWjgGohMjIFtVpxjfH4X7MxnRp7yxWl2kMLsz7GGZSN0Qlpdgr1NIVY9YZY3qiHFrL
sV7XulHUg1PiTDa+dN8s4r+9QJdmXD7LoXOB1bp+1NEWvra8hRir6rVu4Qd5xx/6Nt6GK7XV785k
nU3SaryilK7zGagqvPwJGn57EqacZha4YzednhleLkpix2OXNckGd7CaroFWUSrDC5mTYDnT9+LC
kMQRGxBwJosAx2u3qcNW45yLSP4lDczZWWy2fXLFmkwzHTMG+Al5sK4QpyhIzjJB6VtUIHQNV9XF
On5IAEH91LpzrSFx/UQS5sDATqJKTb7hwniUYFA83DnWBnIvQQdT42TBLo6TgsIR24phFS4MUeyD
4UpOlsD55cSCk5GEshi7R8WpLZ2wyDzxZbSIn4zxNe17xExXCKDKvO+Y0vsm3IqYT+RBrIgjDLe3
Rak4+WdiYw8Khyr7lJJzSn9mGJNiFcVic05MtNrQ3+PQxQ421HvZItyY+0W8gq/OcJwzJBMHggZ8
yoNE7Iwi568O0hZg2GXw8VjJMsJDOeeMV1gqHf6H25lmRPDotjeuQi7zxOyoNmO9+3N0INyNlbOk
t0rLZeHI//lUpgslQ44NHILnLM/Q1Ez5AiqFQEIkD+DbWEKT++sNGKwrulDh1ZEbw8tcIZcY0tEJ
qaC0sP3kfbQfi4o+xA7VEj5X+NcvuB1W0HuBtXpHe4tugYn72HH9GvDn4WNyaMQ7Nd+yPmGJD6Xs
zwEPnQTS1We/i8pcVlG5AfUOuSQQYv2tf9hFKmQRWxoVDjHt/y+oHUZf9jKms/+0/PFxshDWM15L
CfM6OgHVa4gNObzjg6Vycr7qZ/RlcjoiViML/A0Q38ywxxvVPREJSXBAkOxhx1t3tOSzEAnkEVFQ
ezcCSPUdbZoXzUUEgavPJvri5JP8m1XBgDN/nNeTf9euv5ngeZTFU5FDX/SQYNmNm1t547wRxPoP
oXXTmVdwRgrjC4SAWh+p0fa5pmNQAe0eAr8ApeTLb5h7J2qu1mgHXgRVOEICygfxM4AV4oP+uf0C
QF1TPoyOoS0SM9LB7kWJM/0sZtCf/jEi4eQ7jUH780oilKFLXTckW8q/2NKxpr8epheCMqWB9RdJ
b1CuQo5fLgAk/JpBgxBIy4p8z8lzI4Bwg4LnL0SX73kHxSnF8uN8h+LA/gzbHTLR/kI68vOh/PEv
+q5HLWnEDDdD5KTqIVcYYSHWL3T1p5xr1DlvCB7vC01fTTg5nZat3j3iSrmYq4fRNYYSQXzitpfM
uehe98qIoQzQY18errAO2uA7CmhJrbMEkJjGrF1CN4uPHqSxhoZ+uBOTu5vmLdUnInQFado/SPei
rx25TbXltU0eDXDOEuP1JX+H/U5ECwFVrlzez49ECFa0vMlfAtHwHBsAcJRrmeNp1RL84OVYMlgp
8ZrQkwAaemNliBDiSi4Gxb881ONJSSvKkIrFLs7skGg+FwmFjEiWHB3A3Bosr2HcrE1LINPhVn91
QRy+1RjkThufeEPzFWsTeyC2mCMDF3y8Vv7qE9HVkRUJ0XY/qtUj7Y9DvCA0LPv/++H5sc+/9Yfo
CKjTpDX9S7vDdPhxoyVeb3tOdxy/KBcw9yI+GnlddzyraUzsyLAkQ0qd2SppDS/S8XYhG+KNoYUS
JhYW9ijf3k6tWxsFStnhrGM2CvUFKV2e9NKVfwlygTUKxUppT83jsS/oociaNE5MDKJ7boP7M3NY
LXv1hx5DAuXSwOsnsPtuEDR4tELhYoGahgtANr/e/xxtV6jFkP3ibT+zF0WzMxzoeERVdTNGbdZC
RO++ebFQkryub+H5XC80vGokGPDRZ21pTX7vi7sjve8qAAQgTEL5F0pTnkEpsQ3L6hVlVVb9nRNz
j349ZrNXj+UHL/Rm6DkOSEYqnvYaGGnw3dbTIXiP+UKNMBQowDgipmF3lxsSfr3krfp1rshW8NjB
lsGH2v41sJkRDP4uQJQRvGkT2+J8f3NV5QxE/BN7oHszp+2YCYi3oeUzKZ+C0Eg5lqqCMkWB90BA
uVoLD5/TysQ4tGygiSUbxFzDqP58gK7T7SVfiG1Ivz6WkuJ3Bw2BGsmyBXhnCfCJFW3vhKN2DWrB
qZqo2gJXX4uqLANmZnlLhLGtoYjgDenWKbRjAbSy+TUXrlQ+Bovxfyrja3fd+/MyN1qMLb4Cjy45
ktnZObh1I0UrBtGByL+t6Uy+UXRqN0VCyMidrkji6a7fJ1TeN5+/ahUs17FLlB2pP4makw3MuYm0
mtpKvaK6Qh4Xgi28+0dIBLyzChBmFlZTVNCnI2URdxYnflg+eW6oOfuPxccChnC5saeWEcfkQPq0
UYUHBWiTpnfBTHStdmH3KCAo7Mleu6zmKnx+7MBkN3zom0LRF7paX/0H5g4j5P1P6ox4jOL8vBl/
38E+adgNEBOEdfX0Dlnm9ZL80vkf3afkjFLPuCfqXvEpThuqU4hI5cwUPNV6nS5aHBEwDXKwGDL3
+sK/gRyWtQvvaL5Bvc6w5lhzl++jMPBZmsPPr6I4Caz63aDdjdGN4uPP4TI07xxH1eiIf3Xjf/a+
TleUtd8U3EamTFSPz0wyqPrVtuiamz+HNuggKmZUDllduk18fAgsw5EQMYXckJTBKrkjwk2M47Fv
NLgWNcoqscu9ZX4ThpWolDY2WoDWZ5csFQYegWUddj/dzccVitfI7bkvxCaPU6NmIJo6njNXtFg0
2U4cO4fJlJ1VT1u6NMU+/gPNk2D0rp3XceNt49cPVpvBeP8/sPFKCqjcN0qdLRE1WS8SG89/N/8D
T1E/tsCTTc8tTf7q/hwA1Nqp5gq26ypxh6tyrnWbFmdb7/cimBT6055MZpvINRy6b2i5Pwu5gv8q
uk0sKSo0pSYwayMJpIRslXiG85pTRe+vxZcVvCtzzsr99PGbX/5suBDQSQRiLMBciOZoHGfz0tF9
UzWMhP0yq7IWcJkgz5s8GyPl/ojZswDfQ/XO66eldzLXyu+RzRqlWQFlO++BF2tGM8bQ+x9PWRSK
aAnarhdKbnlTLdb56XFcn4cC75zVsxxz8JHq32GE4r2xRMr/k5LvaYgRGHgxAygj//ojER/5TxrB
p6t0p/0nQ8SMy3EYGeZX2XgVAGs5UYC6BMmiG4WnAdqPcgrTP8JiB4RHh0BAvpopqMdLP5CNUeZz
kQGDtUFVH6OTJfHoTmBqA40TAU9uoiIWbshmDAaSs2+a+uDLawkFsVsHN76vWNNs716LoDaODqQq
bUUiwMWvHLL4L4Hb+U4Jk6EiLAxCNuSWOf7UBl5B5h385DIgbU/1x2EUMyOJvKpvLUyOzLA7Duff
brGzd/LbhxKbwyNI6Y+hp6kxFgLd2Y+8XpKhgDXpiFckc7voctXbXUNb7iixYm81cK4DIb8vHfYS
bzZkG7qlAj6SJ46ht7tCoKPAikG+k1X1v1pRqV253x+jwn5GFxVRt4W5ZQ5sOtX4z6nK1lv1TESh
lkh74J4n7FcxojuGDpJWSdm9pf9ie74jy8HVYeiEuhrBLemjw6Dq9HX9ytQZXabH4SMDvebMSM1q
6emu1Kzhh0hzJVVPO3vfwjlasQKswq4YVGxNzz9b7lslwTUItf9MQqJypQmCbXXaA65975IWz0EH
xIk+/JuzCyjLLx3hpuq+my1ukV9rG1ZLt86kx0jNkrOYdHvQdP0YOM9/eX2HSjAMmQeLYSGdVqxU
Fzr7IOiwTKLCqggl/lx8U3meDUp3DCng0KPd+6zbPV+JDToUwQ9nCKhsnk/w4mL9YRV749u/4fvF
qDt42TkcEghi90XSJfloQ+qjr6/Ktozp4mSjX3T2SXnoRlj1gWZNze0TcdUe2wue/H+dpCdBGyXe
92rrrCfa69mzhVXm47ESn6sH2Rn/W5SVh3taFR8ZwO4PKUN/IgLf8UQIvD0esXlTn9rOElg7sIxB
WpCv6d3hzqJxYEtE7Juohf3mQ/RS6x2lP/+2V/t+e0dZeYrFRguSQl5LaRq0WIj0GKSy6xWnGW/j
wFLsr+QzQxSN6IW2wrj3VMJKAHAcbNDzk6HuU+f2cU3ob8ayudCmVvexR89AiEGOm8bzBcaM98PG
8841x8vUAX8uaqM9zYbzQmFuAr4K9V4vb7rrNAO7NMpWsoAqItUMk0Vz+EPw7URsgedGj6kIwI8W
talrw+HhcsmIR53epWtIQdhcCEHXg+mOcS82eEtmPxV7EbLA7HTliMmlU9ciBNoKh22JY4E8zQT9
PPMp8KG00xrCwB/Huxb9ies7wyswG/bBUzgHvQLpR2MGYZkvI4w3TAax0KksDYSR3I57VEMIYVya
XY4cx+7ijjZmZRu8q3haexBEe3aKpl9k3iDvzpQtURvSdJT7vwsBUxeFE965ovgoFvqCWO5oVOOf
P1VGjjn0vJxn6NzYEB6dj8rP2TmYcw0T9VUZv58sTSEWP89aYZ+svK7/RYaYbLS7qhgJwNdi+w5H
0Pv9dwcxN8UoJmvCJtQh01LDUhJGPaw2BgK+uzuHGkUYvxgDw96RBlo7VHTvqR5Ryb+jxZ+qt4WF
yUbPlsH1MH4izE9cgE13aOmONWuVsrbZLmQwbKLRmAuOtSdtnAie2dFAhTRCLVdn/FfpDsbeI7QR
nWgXsL6b8o/EvtyxwboznOK1DWXxYTeDKypH/slvPQmslFW+teUVKlBFmDhqKrx0frJeklhh054j
n8dk1AZDcrOOBeJ198erGBqDw2ryKR8o7XZcXK0U3n6JihEce/XizY0GqmnGFUNSCcgvNblF4a1r
Lyj9l9JA0dGSxuhb1B8zeYkM8D+IcTjs4gBwbMH3N6jQwj6gg3pgqFBgS5Bi3kdtw2cxb//ilSZT
DkBB22nwUPw3Q0EyWNVEZjizc+ckEfMUe6IQr/Vbr1TfCssxEQgIPKaPn464+HjSFId8JpI2rGi4
qOQPdHLEoVVWmDp4lCOAfhDk0stYWOHaqS5sAiPtS2Jttngm7N2kmlfGR/KqsVsCbUM8ZjyWCT3n
+ZsgRI4E89+mpm9vXVjHwQIqW2/smLGtMUvyhUxkkV7FGmiOyqqjHYTCR05XpOmX24UJHUEvpFBC
tgBsiJU23I63dgw5PtNLfcj2BlhsqPdVJL402JnTpGkSgeRa7roLH9XSY8JNqC+oi1MCcNild0Vv
U0WMUiaoe2Nd1Amo5L8wMhKF9Itno6webDqCYAPQS2IzTiiDyX9sWwexSdYv8LnOQGEivYZVnAOj
vnDx43blOONNFYP0dc0TFUXN17RPG6nMombx7EIoneUJxd5nGB9gwSt+/9y7CD7Fil6VdeI9JELR
nLiXJj5c0MRenRxmbQEHXDi8eDYb9tF+6U/5xxZIuuntw1KETV4lOuXowFfl9GnXQ2QQwUk77COp
p32mphgWrEXRH3xhjHZcQ/TK7ThnWCT8JP7RjeA/WBkf4TieNHLRnVlvW4i9yHkv9Vp+X+wekwpQ
qdt1eAznpDIXhp+YYvGxcLxumqXKX6UWyjjbUvaITWsBK1h2FAyUlr5EB05fce/Kzl+OKn5ld6o5
N/q7TGGs8hCfKnbwWjrbJzD14qfkHu4oNY29kLAOy7XSR7AvRkqObpMTIpVhqypQwlJyfQDA75DR
U5SlMMEs12bVTiTOvT6rgXrsmJYLnE+DOhkozo68AQ+5hhqAFjrVlD2k8gICvS5m6W56jfhsOuDR
WglOwWWTwCMlEpjLO7qyw6OaLLMszjm7iuKTlKkCPDnrE8wEt0mrHiqP0woMTCk8IJlmWAwXhUvB
P/tpXy+mRU7p9d3LLnESytYoiW1Y5jaReszjP4yeZ//1Wa83y70kPSrdvp/JmsoFIW+UJDBPlUkg
t0CoGG9XgH3K3yIZ+bIzRmDh7Fru/CaGebWiSMB43rwyG5gQkj1Yz+NvJVmvxV8AaI4YVdsh9tSK
/LAbS5MB8ArTe/sMrk18PLzEQdv1EgTspYnRKTDP4omzgvxxybiXqQYbs6Rex6h6gobJxSho6fYX
nQGHL+9oF7/3QPS6hwObu9fw7IkIFbQ24BtYBwa7Rv8TShRJSdQtQ6Qantxc1X5f/rV9fdYUpDll
76gqOKvRKmkKmLK4YJCAIp5UeyY9Ms6q8rsIftAH1re+SQRbmZYU5hr9DSKhpWat/3QwVR8E8D9v
dr9RB9g+VE2pe4b7iy2yZaM6o1noh6pvWM+P1Id72Y7Pj+j+hUmXs5PHtT72L5qpCB3ye/CkHbjq
5y32IOUpcrmzEyMMnwR66ieVL0iQ1IJQc7fND/SUnZPMaeoxlEwEgOUD9Z8b5+wHZbhKV9koWphI
zCz6QpUwniCV3e9tFB2vpKAUIe9P2WN7OlK/tMTBdVPU+berf2rOfvWo2tu5VYK0MAWLJbaMjI9P
kMASrIyUvq+4mC9fBxMDwJ/5mbo969L9uWQaxAO30zuK8omGd8nkjY2E+/kij35fSs9FJfKRJE/n
zBzU7/9rVagIIqOEjnomLKVW8Weorv/yYyuaF0HGfJm2vwIN4mXm5PLQXSPfH+Q6Ll6n895GkkE2
mPM8CtPWV48tOLeTHdzCyqruR4neKdywAVh0sGgmH6KSN3I3CFCFVGPIGHbvLf0bdQf0mv/g1ML0
PH/Rr9nllLpMyqkz/FWt7n7VmCp5em2tw5Vtk0DG5HybJ31A5xCyr5FAt7jz435QYqqH37XAmxwB
pn9i9rcrYl5OUIWiO7VElsSztrF4NcGgMr20WNanlzsD9GivtTjVLXVyyNzBRigDQhoohZ7OG5qd
lfpTVkxQcHoPXTYDJlI/lCkQOjPEnLkhoFyDz8YjFUeWm1z8D6MY3DvuiSf8hLXmxI9cin96xCas
hlVmyUabqDvS1c5eE1ur0oiKt6oRFIKvNtOz6P0l5hghXbS0xCbQ7SvtB8inDrilA1HVbRGxX8Ro
O7W5bhY0yIHUwDnYkuGEDy4w04Eb0I9EfbzwfspojdNI32Dfh92phasC5eEpEzl4WmLr2y7S+Edh
Ly/rKW9hs8CjNrL2mi6O2whJNUOzknhUF+sjLa7wqX0fu5k/vS7yJVief75Uw+LtoAeUSJQqTcha
rwq/dhEhxXCqXYxE+7M0owpbkjn9ilbJubqGHALsMI9B91kWpxH1UotEjForC7WS/fppuB++wlNg
36hz1Xc+k4JO8A6y/QgxqOYX8yMx0IP3IG83jWFYOu7/KuA6bJLOLlGcxAj1LDbDuppmnRsnB5Wd
XM7yV04stVsLRsQEHk5ArABxOFNeyAueDSLy3wWsvdS/ORpNWs+3h3RaMtSR6RfEPsc8d++yyxx6
wdwccDStwjVhxhmlsQaAcvD/2/Sn030fUYKTYPKIh9T7rLeVznGk/w0NBNXJDzXkUYPrH/tn+j0G
0vvIHulz9njImE4Xjb/KtzADBwrSKMrzbz4hff+E5/Ujyyp/aQe3FmmLbT3yckl/lq57yJxkGdZA
1z0CKVeajMfT5g1Pt2QLUV/gLxMGD4WHVBs2jn3/ZGy8SBsIoSXgnhAKWy7MLoXO1fYTuKDBGsEc
aZ8TeVJIm8O/lXmUP20VDn5jzS2VAGPlyC7ggAdgfOLnUwstdqjhRjbEEDpach6dnBwpvDTQa5g6
4JFfpMMkTu4Q+ozqKNdfYugwQ9xi82nAih1DS/um7DO0Wckw2EKeCuGlhfA6Apu+ZxTVaQg5pt5h
xMDXVlwtEGCGDUhYTbBnnqMk7y+b+sjoCP/TGuuNwKwITACygCWw0HJ9X8n5c6pAZ249Ukr0ZrN8
eW/RO1cuOQ7L5J4Y2VnWGC/rIFQBnzTmgNKjY/PeF+9ErEW2tpNq8eYJiGZuY+n8VEXDcw91BbIK
FucdfKGclg9jOr0x20X78/i8+FiG0N4sEt0RZFyTxrFKYDWYnMpVCxNn62tWVMvXO+8ApQYps2bh
w9urX0gUanq4a75+jsNfr2AJs2KoexU7IS7T/1oQ32AXIRfPBaEdyeimcRasgcwWeUjHBAmN1hLw
1/+VjsB+nJzsiaIuwWuaIfufzTvOWRCoPsCQklj/NKk4ZDuL1ufSCMfTjf4IyaKp5IgAsoMuoXfD
ckCYABy4GZiSYCrRyvCliKdNmzvgox+Od7oAApXV/7THIaQkafsWXAPmDpz0IM4QxPR6xezU3+Dy
ItF/9LadV8nTHQ02xDhKs1BQOpDISMWj3ACi2MyDKlgUErvim6w9ry9oQp1oQLGIEDKi3fWDF3Xh
YdAp82/6NLBIOybfV8wFuh3Yf59BQEHlYsuqA1euAAKiXMJ2xmc0EYKvcelGEfblGq4BMWh89U1a
q+8LE+F6uXYejE70UAdbC/edYZDiqEALXiGZc2UD3ilbCWFPxFyaQxtEPiXuD1fWroqUyVardzdv
gDYz8jRbtiyRmPSV4zL+K5TcQy47qXlq1o7cC7Jc9zP6mo08uomM6YZFU2RRgS5CR08FoxsXjap5
sYZfNvNDQVpjndYtCUgwLvPJr99YjG3JgByPr+Ws61x+z7VyIwDo3IdD10VN5aacZ0PtmB7G7nAv
9Szfquk9fFsXi1lx0GJre/0Cpuy/GdHjp45epmwBnj0XhvilawP/K7jGVjwQO4dF0fshrbHTeu0y
pIoGnag+uWfS3aRFyoayO+4RyR7Ig12DdYITfR5fFCZnZxPBWII1c6oOSNrAAqrKFLmqJlZhpO3y
6ZCsviUsPY6y39ljHfjrohJzQbsHccSBoJDvA95KrnlcOW7ypQf5KGA2RIs7N+ewZGCH2qZUcGoP
hqSbFg8GWAEyg8lA2ObuL2u2ZVpWCCs3T13fbjcNallB/5IFt0LizEBvHnWAFIsifPO+s2GognEz
52OPfuGHJdDimL89L/G1Ptyx/vB9Us+2MD9+h/bQTs8abc5xb9bjNfdHIcOd9rc6s8eVNg19k5z2
2Uu0vBdnLAisQgJMG9zI1OwhVGvlgPmH3jOK8sw0e2lzUn7maLLNhn41jZ9C5UHqxZzhxnCEeDVD
J1h4hewh6DvO3b8VFpr2xhiEvhx0EBArTOhoDraA1H5JKEgVSfrU7+xNn3U7qABu8mQ4h2su1NnG
L1CMOYteyW4vsiWWdL+WcZg246ovzyCyKBSfCaLtB02lMev0nVbYrNJTTCXUOdlyogAnimRpzH3W
+MVPEOFAKTech6vC4phd7tp4PwkDfGiq3LKJS1T07cbmNjuBM+NFQ8TeQlEFV/Mwkc3MfCdUkSXQ
XmAgQBLXeKwM3QCXzsCqbAihLDH68qLShZzgLrQLY+hMsLOLfv9rP+czau9PAGCxrOiI54priLqr
RCufLjTwuQUgUcpOE0Hx4jwCQ1fRm5Pqw7GnHLeQKML73heV1SXbOvOrxpipEsZOt33CmkRhhU6i
bLfqpUdHtPeuxwiheWmXynUr7+tY4bTLU06sTbzVp3aGvjwg3jnKXerT1wSMPukRC82LNamBbQcJ
+beTZKDzslnoy5gSGnc1nRzwZ8f4rwpNT8eAmT0RqMdypRELUxvm4rWRK+CVCSca7D64lpjzytAq
J439Z5HYDYuy51dt7ASv0doAHDQVm8Mz3KIHQ75Dh2JXDAHZoOQrEUUZrEP3BmYxk3501AYKOJou
VIQz0+D5mH/dtjomNLXD4aVXlVjTpZ+kwAg0zmqiqVpXuPnPzST3tpiaxGTDwDY1zSI1ccEJ52X/
jWeQQgBUidbp6R5UMBOdAThLMU3+Lqwji7+T8OoGsdBUmQjkwXy/Sp1RQwNVJSlT6s4CW1J3kre5
2tLDpjpwg46hrsG9Z+n+/afmnGE728wCmFovfJ0NCrRKXmwhogNX8UORTYgoDcOiZfFA8ovE4VHo
gyiAxAfxBGdjAkhKgpcefnTlg1I8+RLCxhPLOHzeVLrTxvXxvk2ahqRmsMOjJiEBU2KODgGrhaPp
AFa3AUB2RS+YrYBxNUa3DCwvXt35xvkrODObdiz9f1ayaBOTVHmCc+OBafXfuPQCyGwlnCEu9ba9
WuLNcD/zn9XwStnlJ0nBlebnZKM/1dTLTLu5g1xQo7jwWW9j8+9XD46m4j/2GItUnAI/k3g8sxX7
aGKw2CFlIqKOSBDaatD/7BFR2oa7nRw1d+GzOmGOFBkP9SGx75oyPBLCn2YB9PO1/xshsWd4LAzx
c2lnZlOGvGrrKYPeiVBWFe9yXmBolfGRjw61lLeUlwZIbysPucwtEOHkYchKR9BUQLuzbpJuzAe6
uVaUmttMAKGLSvCVUGJRbPq7GfM0j2kx+1OmX4eZubMzkgQxwNfoscOViJIUjtIXuu5hBw5Ht7tL
TwTUWnIbGj9e9gY/jCsjnNrJBGgxhtC8AOyMVy9GKoHU4eJvZVuKeJ2hzYJqp6+0JBPTzswYU64o
PNcvY6WzgGkWDMHUWAv5nGejhUSsQUtZYJSv4WjFK4s1wnJ0HoO+4X90onhW7OXOTiH8+J8Ghv7Z
6dSJ725LqctMKSmAXH+aePzIIsGn4UTpx+WbAyKk6qbToC/ucryY18cG7hreAZTBq5O6kQmuGy+o
yQKE4cNII48vjDl8yxCZw3yGoiIXY/Nxp+lHf444Mx74p5cROlVRCJszhGSnlpYxwdM/vcHs9v9N
dKFETkufQABTK2d8ESmfdHd1J68kWE4vOaFSwYKjC3FidmaPfAnhJRTCBliDezmOPeIGInDV4SJp
5RNrH3QpuS34SogTcrDZBgMp54Nw+1vYLt/8giI363fvtNL2xB3OFOaQ+Mse0U9gG0fUQtf4RK7Z
VmeeE1r3fv2AUU0j+Bvy2abVG+TTYzpV4Gq7Zkid4jdOedL5ZRlsvayu3yGymVrfAIbEvLU9PtI6
NVKXTWZTdg0BML6WPmajUaNaKFTjGRmMYleN4zpN+cnEquMAxkGAP3imbPlc886GZHyyO/evvG8C
1LNExR0zZCh57VP7V/aESmBjEilD2hNM+spAnJTvJ0gqih1y7jI5TTOd7fOF0KCZo+qG8WGu02/e
5pDjfbkGYIG7h5UiIoFoZO+7X/pxNa4Cr97IQ2W+FoyhuKmiglVHMsrFo+SAuRCFXcgbY0/2UsTo
qJ+ncLzNKTYOpXKB9iVKVMiWr+3YfJLesc188hdtSSfTS5NVHdWXkuSuGNNDHiL4PO2dIAag7T0m
z4awMhDpF4ByEn1rEDUWweE2132igADWj4FNL/F6SuESCeC3REnpy0MUJ2SITh8rT4S9jR5V5IXf
sM4W5KPrSeZBepauDEqaMzyXrTTqN00+oLtkt6KG3jlYOE/fYrUIjy/HgyH/mxfxYuD4aXtz51Sa
CR9XZnJ6c5bj9zyGoNhqnPfqW2XPj3EaAei3KXxOaXx3CJo89VxpbOBRD/PSRlNkMU9Hix6V4Bdp
hICnx3pJ15Q0bHvhBzsJ742QpyewCra8VQOb2hXC19tzgLWE1ranM36cFQ4vKjraNejrVTqCFQT5
5B00xeG2QxJXufHqYxUZUoTWrAO/Uf8wSdYsQY480T2znv80QH4KbbW9yah6SGHryHaba19JFPA0
Vf5vRvQ0L+9kzEM7iA38KveGNYbNXSttFqRJ6drzY4aop64yKu1yQvOxdx3wFBQYOLppuJxJ2ULF
REcxbS+s45LGMeINKlb/EoPG0WUsDZVIRaPIp9rHk2vLfkMieQXYok1RfaUZjkY4m77mOx/I7I79
lE92aQRTGMsEFBpZ+yQw+9HQ0l4spyNF0nk2/PB00jNYKraBFfDokpp15g/qfYTXgGxZ1fnOD5fy
EKiEK6D6seC4R7oZmD1kfHkPkezmFe8DxCU+0yTkt6Gn3EkuCzD9L4PaT0/Kcf2CsgpUaUdOSdxM
0QcAcAb6NfcqPP3qSvhAEtvMpiloqu5a5ousw/TvWsMLv2M719oTOsw2x0Q8nWb86f88RZhwIh59
KVCyICtVt5jvUkYNh9EQyJkgdFsW+XEE/Z+yq6QdAmMRW9jRCENGE5fJ/wmclDuwM8LSlGqTK2yH
9pcBScj2pqARWxdNXNgG6NrNOnb2KwVQKjiQOL8Nlq7W4BFjnUmgtDHjx15yddP2qL7vOzgm/kpp
Fc1lri9OJswVa1x+SU3xCAl7mctvvoXzhgkW0UjKgf+Y5b+5fwZMingzS9x8VCG21x5aA9/D5MNe
p458yryQ3g0nJer8y+JwEPQgOrSBEUENvprVUp/Gy04WNgry2QZ52/D0Omr3AKRqf2EPOyovIHBB
mN0z9gMw4ag6nU7jWp19nKC+Hd+0nRNL2m5sF0TNI1r1Xr/WK2n7ygIep9oE3sUQiVA2FgrCT38M
enD2kmz7fB3revL4Dzos3Nm2+9xFSaNCq84n+VZDM0XUgHSsZMFzlHHeU4JEtc0o6wBKbjeYJq0k
iRPZ8csga15OJzfAJLSj4TX0tLpqdmwN2G3xGcjrrxwz8cAQS8iEqhjpCB3NWz4oOgUg5sBdcif2
dyEZxgcLsih2U27BhP0A9pGUdH9Q+msFbVqj6bclni5lnu/RVGX2dTWjYZpHEA8EykAYUMVkUuKM
3bkIzERcFVc2iYBml8bg/aPDhSA30h2CjDO2YEVVHW0Rb64jiPdx6coFt2ymqFFoWReLzlo2Uidt
Mqzlj2C6Ft8lODMo6KnM6OMxxYvko/R2KncXYxksHu+7JJ8gUBzY62vheMvNFFC5V/yFnZaMVc2E
NyeHIe3i15aof7LzOc1ZBTBTBrWPHGJOHlylt9oqficKs+WfyENtIzwTloERRkS8MkpPTuBRzNA/
88s61q4nup4HRY1I24hmt+TEBwmCXEI1Hu4szqu09NmPlqoikFgPUR6Ct7bqO/5++DgWAowFtbuw
U53++pErR2XgWyp51AieYRX5vaAoDkQz+oALuN9lsQRW43Pa6/a42++KnPpT0eWOrDtIq7j1FZ51
gZqI4dGhfHfttVIIfQSXNDCv4Zxn08dwxQratLna68JZO6VZ9aFs8eoybBkGOITucJOYROYat42/
kqd2iugw067tWhNQo8M1xhyQH5fmyeZipKj1/n1juAU8kTqvQJMRuJ7/Wpf84qkXiGF1CitU+5tx
SvGQb7BHTIJ3RxXB34kxzdWb/wAmBkazE9GJ/2OL6AavO48x+POVeZwQ9nsQqQIqYOt9v+1Qh0vv
HTqeyXyTDnDw363hX66Ukf2pILekMj31hkjTY2ViKqbN7ni/OeZupRe1qwu1GskVXHoR4OTZULL3
c2eqPIdE+dMbTm+zXoMyy1Ebo02+xt6a0YUlrNNm28HjwclxIItGXpRIGKsyrxncvZFZO2gfyr5k
EBXnq0KsF68H0RltnGCMGkHLfLP4/JTcUv9GytoJzjIOzsBQHAaE9+y1imOyJFSkQw92uuP6Mp5I
ter+1bdpkzID96820vyomGZwTgMiTUO1qcd1pz0l4RbtA6DEFd7MJHQsfWAQfg2u7sY+AnFcwmt0
jC5r5aWlY9pJVNM3Tj2bH6F+HcYxykfKmBfu1aY56PtFUSyPrU0uwqvnF29NOdXvZGtwKn+ZjNmc
SRMPuhTqK2inzGYrAqg2GZBlRo4B6ieIwY/Zg5r/CYefKS6yq2YdVwxAHw9JSuV1KSM8zgjjjTgh
EKpA6se+dEjzJ2pyvfNwkGlnsdJKOFqLlu+Tkyl83tN3D/lPDY2xUH9p1V7kUiQi8ijfNZEjGtof
GzGf453B2wT69M5hK9XHfR7mFdTHtC5WFL51u0OhJPf7exHAmbbfVdrdsXio2qxRIfBMPk86fQ6i
+J7cbjg5Vi2VQvazi9yOl6QY3roBIPgxsl/Y5O3s8Kh7erwip6wvTnJZrnB+uO9er8bext1w4bti
oOuSQjfe1w9C3fIqs/I4Jacy5e9nWYHbE/5JFYu2LWIaYfFaFQZabfwV3CPUxgTTRReIH5Z6p6Sa
6Fo0KtcQtS9TPGBCHJUQaM/Fe+7YphJU3rBbiVub8g6eKERM8KTEdmIdzXcWJOX8ygHIHb2iosIJ
Im8zhrNTHp+tTx2Spp0wY1JZjSSteJ+AcYtyH87d8TARyaA1X8eHaEb6qDNDy4AAGY0xVtyjkx85
FgLirkJhOUm/3kpDnDjJEiqjgKsPsPYsToH4LH8nKH000Juj2vBtMHq06Ut/S5VS8o0kMUXwz3B2
mFTDspEk81KKxCBIEky/VnF09Id8OmGoandxniXPH6+kggh50ngBOvUOeE2ZUchPUJfH0SCiiiaj
ZxBtAwaztIfDIhFExzjdKUfK/W0k+d66VMZ6lymmvlmoDWi8BXru9yGgHPb576mmpuaXs/Nnv4E3
bAYBXRhA+y3hG/42VA+LR7q4anV5wYJTNqq1dd7RIJHFLOs4aiKoVkVdW18RZynpDw749p5fSuIb
qF0NIiwz5ubXQhqLRE6cWHlsj3XuMQ+dIkyO86MhXmoCuAXa9k1xiD9873k1gsubIfd48GEIapW2
Xb0/NM5mxKqnDgVmRR+zTNJWlQFX135+4h7RCtzDz+t7XIwWIB3VF3CcFK/80EgEk/qQhjgLrp3a
tLxHruiCPpBkPS/XrQTXcvCN/wi4M2EfLd0+iDb+16Ox8yw/svMlEijtm/6daJFNlDU2Kygx7ZQC
AMEZdnwkrF9RlmOBATn0gor0cvRyLLnDGs3RZ64vmzqqMEFUGlvZTIohF3va7/JrVGd+lRQQeRgz
FKFcbhyPX/JLiNXyKIX0ERVewy0ttAYjfyEfttNMNYZ0kP9EVjTLcTMxZzqFsSRGXYpzDNfJuOws
5TWBkFPu8ZDfCJ5LH/BEcCM+rMsqHJVqJi92v0flu4j5p6lHG7NgQAHCnxilk+eGLOPXR1eEM8w+
NMzRdueZw9x6qYu8kzD+6jdLXqgNdLxAKuHmSR8CX9s7txlW7q2OacK71QRE20QAzFmAyEMC323r
jGJBiqpj49HzgmsN7Ezl4K/Na++cdChj0c0uBI8X9Kcp64XvSheRY9SaMjSAAGQZJB2St9K2P5Ye
eiyLFBVx5B6yoOioNz5enVY+gjEtuDrue0MBjEZw05Rq++CW4eFzyuLIo0FPq8GT6Fpw+bcYSJNW
ypzg6iB2vU3jlWJSqpEZu7u9EjSmT+NGGShVd+KqJQTp9+3KN+dNOOtZnL3x6EcLg3dWZ0+zXiAS
XDDHiJFc9CX80zTDsJq2qVEq3/ku2S6fgtDRYRk3DATY+VSFxC9E0i9nvQGBzVE16lZFyv35z0QZ
K36ARLRSKLzginmzLUGL7W7Z911q3iMpLtHq4IDDin8UsgWUM02KIaHIrdGN9Arj9l0gpMmhIY8E
WLWM8do6BeQj8xBEt5KGhwf+37HwZfOKq0yXSNABWiw+3e4aUsqBBpTHdQgQ9MNY75BN6PDtCzt8
wpY+AmYenHfcf1WhUHzRmhBOCzW2Yv1BTXF98HW39GWEtfQA27m1BO1RqfOMdaXEpK4Dsock94qH
+zeaHUiBGcKbPxJAtWAOGrxoKOFpi/51COYSXNEI3P88YIhvH6nfKLeFQlWIk2jRBKsqwP/jn/TP
oEXP1h6heeDZSA7DQb6qjRjpzGRLPlepHVh/9/PyCC6p2UJ91g0WtYwdaKaAYDE3KCpW7Yr3We4+
3aJXq0aN86U7UwDjHGk0CNbzkQ5zrE0fBGRZsKbAM6JSCiSCMhAjaD0X+pL4OMZVcDKIBDZOkU7x
eRs6j5evDP2NThLiOLod/Q7pWwQuCMMYopGOHf9HIJalzen4BS+eReMbbxZySFDp1uWgdvzHM1/9
oTIkzkm86frJMoyK7r3gZLeeXxdD0pBljMBpALgIx5N1SaxyT23n1RRIsgslGoJS9fwbBds0zDxQ
hT4Ok8ZM9MEUxSXb/I/1mxGYaQbAncOJ++EloaM5uprzmMJnnlAPEXGZhiOaSEhAOLFOk3AmNyKq
271iFsypZmI/vFjAxDdbw/yK9tJ0dWLfdTTJazY5Ni5+apf3JgWiyymoKnBsKu+u4NXQtWLSpbA7
VL2D+LK2xjI/xIuoADByONTPbDYEVuKSqrURtDcGO4aXiWejUJAUkKa3ESf17jmRtiBF/DgRq+u8
LrxyJH+5lWJ+6NSMPMjueo6gX57+Hb0AvQjBzCWNF/kt1fTomudcgJwtvxLnQ63MjdVLdnTbUpw5
thEusfXmf3nm3S2J4JMfen/NpixOuZB/CfSKiA6SSg9lqYWuOopi9w6VC0/bjixvIcFMhtv3c7AI
Q4QqAWhZX/KVUmP6feDWYPCTTZ0VM5CqFFIgOV024zrBcUtwm4f3/mdIcg8e1BgLKARUTnmFsOeu
060Or4cJQC02TmIszF2OheURXSsO7xjJXo4hFOo4lYd+FklgviJ256qCTt6Iw53XBvNA7EP0D+rE
XMk8TptXGyLwbwSDqnJYpamGDL/w6DddDgOemgpwgBFUE9Hgsd6s8xD8zFSwk8fi4kId2ifAkpb/
KXlfHWIki4DvTtOemsu0y/B86b9TmCtLutn3ruVdgKjodLReBpbwfAXRCf4yevLuz7O0ZYyCw/kj
P3v6olKglv3fVdv19y67WS7klE3r0vqilPhoiQDJ+XtVg3KKKbrknT+DLln4j5kZjHD5yJqIExK6
1WktgjEOTr1gL1oV56mKVkhfKfSre07iWT656/BxG1A5cuh/FB4DrE07VaB6spgVWWXngjnRL1pb
HFFC94NlpZclh1FhSvn1D+ca4mjVYxQHZB7gEetm+KfVb4HhYwgqyjcjoCOJX1MpUOZT8a0ULCXQ
XRWkxC+n7Svv7Bb/q9OAk3MPt0VaEZuK0wbZxzc/JZm4XiOAfS2jKugntzKT6k8tgMPROsuTZKFB
BZhkXg1B6JKdiurUdAjhPOeSCmNp7NEFWWG5NbWNa334rmC++ZIjRw4+3oFtUrQGQeWhjRYARfRM
cM2sKltC9yMBazbuMwmwhonjmGLNik6vjkGpEPNO/A5AS07m7gtUb+8BqnF0ODFSE5agiM+hZgWO
l2FQa+dywArOhkpFIV0JZ8PKj1/Qf0V/n1mAhwfNSqoEvbswycUoD5AVf6VHdGP1J8H73+P6mWum
RC8zN+sJ8wjvSvAPd51wl5s1n9di+ac6ubVi2g+H8oh78pkbRvZR7rCHEW9pLzx+b2OiiiFhJJp6
4PVhTPqxpq1ITUKhEy/OpyoYgD5wQVr5S8omzZeQJrjz8jQjpmBkhAwHNad7ysXDJEAQTUfXqkm8
2pv3smUFWdC0MmRqS88Uw/Tx0bhNKMuS2/rXxpHniT9qFdtoWWZ8WR0swJszygUbQ7ipMu3/X12U
akZUzrBscGCM0w8mtijkTfIalHPUgRKcH2a9788Nvd5PLB2zb1pBoCJ05xE44D5vaTix7mPcmVyX
IAafR9LktWycNiJMBocs97Sw6KvlZ0PYeFzEfx885nRge/M1k8xlxkOpW1LMmnyxvF+NR5fCuh6z
m+YVnsN+4lYwCiY8ccpHGsH4sb2Zg59SmRKaV5id5SpKODDAypSSHYjlmxOXytP3SO037N5l8OFS
VKat7TCaAHPYsdeW3/9iQi5pN6ID3W4JLxP/dCotkZPwlBONHVM9q2zjK45LxNFZu3UjN/306xZW
w5856geAtW323EwzHORfZUluE0jmEVwjd+sStRgwGKJjNIpRyi/3FX3O5wQCU5rbMPJqzNEMvRDZ
PSrh5W8CPsYCeAMB32B7YiU1JLZKNxuQJHBVhyAwRsFSPOGC2CXK+FM9/8p0HxvbI/pIIi0Bhwrs
Ni4vi/eGkUecfIwESqt8xMJhjzYqmasCP01biMbPrphMEQkvAZVFe8ILyQjJiJzlPSgHjXu+yTJ+
bwCSLIrXa7zCmQ78GG8z54EVIW7IAfcaH5+xTopwA8OIPNbcITfeYk2teTI0w9GuoaYC/ORHL0Rm
jyxYXPMElbD3PdtVn6yNWjwRBe47t6nFkopzv63375OqXmnrWduG6OzkXOBs0U9F3lWukCX0OG9L
5cIH0FtISZ5iQnP1fI/O6qmIBqYSIetAeBlazgv5DsNSyc4cN/KrwXuova5Eg2eahkN7P00Z61M3
11kYC1IDdLH2yWwLVqTRFjFMN1x1NgynBahoke6DWqhQf/kNZXC99DyvqVnIPuw03qOqez4uS8g2
qFz64C/mAO8TfEanyI3oUCnI2b+O8zhzuCi+UOC1o5W83GVX3o0byMlUxVZxrA3TdFXWivhO5Lw7
no3MuDFYgWYrr4LasHBJgahrfGraGALsA75bFhU2LBY9n/lNk/66afiU3FkqB5aaq1fTA/wQ8nIP
E2NPm4MoH27uC0ykdsmLkrVHw+LvyjOAylcNmRkHhCXm3BoedF+pm/e1BNePrS8XDJMX+ywimAvm
syzWEqQP8/V5bZlcowAn/HgYpTukrvHi+NgDUGN3e818WZemd5wKgXeAsotr4sEAgDREA+L1O2z2
TIadfJz9Ya4wcBYpGtLUSefLl8C3bHZcV8MR5vdzlXIyiGuzFq4zIP0LybeS1HqudFHiCn5MlfMb
mupc4HJE7xJj1dDhk+SFCvJ4cX1x0aE3mYYgwa/UMIUZE6R5gex/57/KL449aYo2xEeYuFSgTD7Y
9zjL3V0TMW7gNjKvn1pDrzQ4HQAqIE84UTOkes//mEsTDJ4V2LQk1H/WLFP41vMczhdnOOqnSXJS
XZZlN9VLvrzSvTTLN3hF0i4Yfmp9pjn3QsqoPQsUI9t336bQUCl4Uy2jhtDYuGLYDcdfaqsquogM
fh/XIiXQxvlbHed4tINtzbd5ggL5d3Ve99NUgKVupVIYPvoXLto+i2/6ppkTMgYtPuvfEWIsK05F
UWkEveiWLz0opNKZFG/YswIjPmBfgyecSD5oy3agrTlXWYf8xyObZ1KmAGPejVXpCvXv/gMiXFfx
/CRCCQ5+LJirNKq8Py/eIpKIIV097yYOzAypaavo71smfREz05q9lS8KnxF3ZTdTenFORDrjCJSS
oRw6RcUKgMUi8aNK2HXcxBXwYSTQJUVX8dhtoXAf3vwzfBRhL19hUcQSkAJo6XMUMctoOpyMNtKQ
XrkKTrDaZG1Hm1RJnYATyFFVutNrd0pYPVWiRpT+MsYaKUQggL+HN5BVSWDzoUXtnD8X1lmHyGHt
8+Z5s9lZln9v6gciNO/l1xA6brTH1HKCrO05ExTxMArHsdeKMuU7w0qYgbbxv2KuKUtveQuZ2rUs
Chh0UsAwAmqnFw+eYKtKczQzwN0EDCa5kr17Fle4MAf/4BK3bsTTi4IckW6sT2I1AkoWjkFt2QMN
A2lDWaT78YIcCSPsJC/NbhfJs/5JmU7NcPc93YmzlPUEfTJebNGvfzV9BB6G95Y6nzjQPEm+M4uO
1BEk8iyUT7GRQVSt60T2kZBN0qRedyG1N4DO8EuOepQQcflbJ5CCAvlBrzOKiBYUZFLx+YyU40xh
OI48wUI2NmvwlbY7nXUZ/9FKbgUs1F5T/6Lk3buDUg9vwJwF+KBCIRRKEMMAMZLS6tr3zvQtWEVI
4xcJyNABfifdVyKKfIG9+HfOmPO7/QObMa0JvLf+TTYShDXqM3l+0WrMV1M0xL9sQooYwMOBosI/
su0cCdg9nUV52NfkhQdYRM5BmGYa1cPfXHkHKh8wRFm3OWLba6qhC+5bktbjFX6ocNcnZZhUqxbO
oVIFKbC3xqbRuWpCqgjyczGignY6dy4hzANQGFqROe6rlHSMqRIYQRbBgmB928L7x12x9Uel0GL+
p8xwWaKjaLRgHS3cL83d9vfuLK4ry2hyROnB1WGLaDlnaE+VpVGOXxJtOi8UTOpmMMwL+cCSHwHY
flKzz5tBTr2ARp8olPOhzFUsdnJR4w2sqLz5nDnriclWVASwMRHzxBalXUQoEecMFA9w3Zr6osvP
3n0nbGNV90Bpg9A6BMkkBZTNWwbfcwZ+WMcFkabwL7NCdD4R8LOFKL1lCFuEQNFdAseRfw/Bapk5
xlXcYD+OIik8qRmFnC1IbRkLeUSZthBeS9/LAhqDjgBPgfFa8MvIhXvk4sajKn39tV9IAjXfEEfj
vLYkhr2mf8cgMeIGYk/ZK52o4U7gHCNcnZ1gD6rWRI7I2YPd9R/12dsQYXBgi0fNSvARgXxACR0g
DSOtHqR5+h6GKjE+ZnbN8gkAQyvxf5wpqpcCgo0gCSO7Pvuoyvw7syOSJ++80S4I7mwY1EFq8yAc
qDtysKVerQnplM+cLccgtz3RC+/vK0MM9uSQsEf5qaidqPGOk9hKBCDJ2U4ueQr+vYJxhHpVzhhp
hIrqJGJP+okMjyy2sduYE35aO+xfh87Bk7FREZ9BA9ROwc9KEYeMFiLhrL24JGMwcgF8ihNlh4bM
byhIBThkiCkhWN7Qcr4hKwL+kB/zJDkCgr6+nlFqgKWRB+SkCwEibdYNkiKJOwLHwh1NBiIefycI
szXXCn0OE4fNDcQsFl8pbNQ6T0YSXUzAa/TOOsff3H8ohVgKMUEwXZ2Pe29bcP0A1yiYHj0wV5iP
0zm8qt+l5YFcSsBF5BWF0FDTB36gMb+lLePjTWo8BZtiFUgrkXbgnPMcpMAvTr3vCMi0jjcJvx7h
3b5cgO3VvjHIu2W70+Q220uzqzazQqSFmGSCb6e0PQ3Cna3QIg28Zf/+Sjur87g4JVR6T0pustiz
lz7PRU4YuXEh+HlKVyiiEhRtwcUbvZ2xfpxXlom9xboYoytmRhAG8c5uKPPYjnYE0oM4o+LWPUO4
79jZmMsEsgugnQRG9hIFq9zkBeafESiaKczXk8BoC9AVbWYQJBDXgN9/xtx8empTBmnUZtvz5S0F
7dckUrO2fOWhkZYqLVA5LrtnK4DLHpgQui4S6TqlqPvJ0Fza3eeKKWr9BF/hbjeOhAcZ+WKGjYzE
UxOt0DhXYLbVZ3eNYEDqq+go2A1m79rAiBD6HIo7MVBrfPvITDlJYspBQo4wVhzK5M5BWZiKJiMJ
BZfDMenqjCXca3GVJ2lr57TGOzpOho5XReG8RZxGkTAmipV8r7fCePtYR+PMrQYyiEMLN3rDnGSS
FGywoOaCRVoLrVXAXHVXQcmIZErawJxuvNOQtRctgdj1gK+bHMoyouer2tX8cV2ofW4PpL3oRdwV
4VEUJw3C0AZigqvkx7sgpgloSEUJI/EsCHCs6/ppijffXKcSTjZ1EXRVKHHz5kXEbpfISUxh5Lpz
Gci39QH+Yd5abzBxqT1RQAkFYINdaqFDZQx0iGGl+KwCjNhc4kSajMB/0qOx5kFK8lEdNecj2mog
J6WSlksVP1K7yalfbdkkbZxCeu2F/ZCMD5c6LUDTSxfPIKzhIB+JAavBjVN+OH/BxR4AGTEPGkTp
f3jUYVkVskXCB9dbL5F0bFwG6Csfe4ScSicThlkMa6qV6WT2JcAI1im+fJYP+vw/fPn+xzYISrwS
4zIiE3KzHyLZvGbZOehZQgQLXiQKw8+3j0A+7BeLlZGogEcPYoZBcbDXKwDLnFaAvSpPoMaBXebr
I2n0w+k7wkFEBB4TuLQJr/WRcdrhlY/eK1Lqju7yxRMkxclRRfl7ooLKdj4lYgjtFSszDOat2Vjd
zasaeGOXD5nYJ0N8KpDrVQdm627oeXzrakaO3FU5dgg9NSxIt3FCV/sHmYw7Oh9NmviLk2/y928C
axnMIY4nyNDXINLqqjPOSipbdLhim572LxFYc4fmb7ygTZ4HnwqHi5lCuJ/idcaaByawJR2sXIi9
DnKXdc23wANAgth9Aaz8sdhHQclrN/Z0pV/kxgYsRC5mgpMB0xhY3Ze4T1AL51v7EuqC4HQQzAxB
qwrY3lKY47qznhY3o/71sF2ebVPkccX34l+zoOgm6hD8pB617rJCqerqdGhkUdoeskftYxrpFzZW
dnTMfSPVWU1hgmbiSoAIBrS8UbrjrwocZ8VSHJJcI/P0OXsu1Tbl0AvNezrDhlrOH7rrXfBbuLyk
Q41Umcmk8c1dvKzpmcxFrkgemyjer1+JIGP+3EGQqZpybVl2Z6w4CuwAPqpouPPDkG/4ERsi08Um
Np1zs3D4hzCsmznNTJXu1ANG1bNrmSGdBz/xRapAlz9cbmQWROwYc4vmKpT2pXm71/1xxLR2OhRJ
Zn3DU232Q2z1fCXkOCADybldj61YEVWAWvXIoVV4U16h7cqUXX61jwECHqLK3JFuEILtd2EZ5/9B
VauLrw9+tZ3ItMxAlO1vew5a61j7sxHuuTiyp0WtaEIGPNpVEo5OKsEGzppz1UTqsLc7Vi1OAK/y
v2C/UW48lDIG4ZW+n8JIOXXLmmPxcyNpPLtfpXVd5nvp0dSaiP87Go85+PbEjDPy3f4SLcN0/NNB
+UyAKZHSSfo1krBW6vzCOF3kBYnbUJ+EI7xv0G7ogeBxlonrGp/CLLAPOGuwWUU0gfx7gkpnG7DO
+6wFauXjdOfmRv3C+H+Lk5yks/jBt4m0Vble9UpzDpKkm10/JN1NjaOpOJS7Lf5zArn+RsYSjpU+
Mu+auKXPWpEj1whVgktm6Gjkofg9nYXqsl4yXpJfl5wJwMeo2ZPn0iVoo3+67wWvKSTzgSrvf720
ehL7YTRXcas/PJuy2DDFXbr+T94gxqwcfBUnL/KerCSLcz/dDiNdOjZpwp+NFzPWuoFdBzB18I9P
bE/BLS3U38Kf7fK4R7mPueMVct4w1JSXGf+Lq1n7EuM8iZDEcRVzw4aQgscnZsw24L4wBKxnFEeM
nYI9AIZHZeGWQzZVOtg8Nl1siE532qe8d6EVumoPSU2B/cPTGEMYh9s2DT3teQpSPh0LBPxxUQ2r
qQo2MKhwbpwE71EbM3ulnCwWMrLNPop7BGF3c9z4Foo2PVqe8Ht0BmuZw82KEIlNn7EXBJvdpzXV
EWCs+sqxEW8ZNTZcJNkUXx4Q3Hav3Tm8X90VeSaJbRgcuEKw12iapCvGorolPwrn6WpYQoyBMvrI
YdWLVZp/G7yZy5NMonzw7aC1IhEsgF1cbrONn92imvTs0jBo6ojkk0v/zM/Q90VlXGz4h3mUfoe8
t4YhcJgipzQTbq9T+dfjZb5RxNpipnGgaRW/I7rN1QULkRhjiRcnXGbnSX3mFazKLCC/piIKzrT0
uf4PyyXIFNviqL2yCPyxtWBgOzZte1DLjY0QsHPiBcFzYQ1akBrgc0XLL/+olPKvdQs+JyDreY5f
76v3CJ2UmFC8F3i+KHdaVaXmLqsCFDKNa6lMmmQsSvQoLqh2tZ8587MtZv/xyXGr4uk6PCw6lWav
qD8u7JLs4ghhu6ZCfpndy1YE+9Zl0WRp/wZcTY9ry89SEqlHAbumZrTsLxfrhCfrOOC5I1Wm7NVe
IzSkNMjve90xtphmns1WEjo1EFcFjGX8xJcita+MbDZxKJpG7Kuv7FvKIitIIqauh0UBV0uJ33Gp
u9/wFO3ZjsleyuMJn2TX7fMWB1CnW42W8vYmdvCWZq2Fkb4OqwOXGIvK6F7ggVv5MjuZ6QoelagH
TxF8Ktu0VkPtOO90/jxeJfNDNZWePTM0UV6iBNKdIDPO+df9BBxiWp4jaRheFL5QUZk2Zb7ty2Fu
PKMSZQysy6/nJG5AVQuX7tesYV4tZ69klisFjw02EVdB7sbPr7OakYoJN7NTu9NRl6rTj1cwCGgl
ZCeRuCPta1vItIppAiaAMeEhOwtFTtDT0QLl8F2dzEtBIJ9tdrcxS3FyqF5fnMXUrowehtOrMMCG
9UtrudwM1DW48mqC0hMYnJ7l3TAbOMr7mfcd6C3FlYn8wwKbm5ZjrtgMS1RMHQ/ls7Ztf4vphMgG
ekobbSNXW1VJQe/GuOj3vwpFzWSaPeWmDbfb3jOqCqtp4k8ouZJutaQyD+0oDCyuYvEItJzoCA2e
7bxWLEGHMMwOnQCbCy63jH3g6+HNpjGiC+WBnlYvD5h4rjcdQmkE4ntxnaOTBKtMH/NbetBXPehk
Wh/MsEnrBNHymOJhCFfvxfPI0tldPybygWeT9xn5Z5+us4Tl+X+HsbP07A2WbqqnNvN46oJxc75h
5zHrBZLEz0BacrvC5UbBi5Jc5RrGenyLJbBDAJ9Ie262c1bwQlTDZhRorRpCaV6yVW/WSifInfcd
SglEEBMdCRFcRtXtdwVhbZ7m+e27VAw3j30tb5VAizqWX/HwntIkrHRT3nQVVHN5P68wZlZ7g4/Q
7X/cVBOyja4hh6xGQV6kkoVfKGW7hXq4NVNNBB1Z92b8E0P5l8bKKbxR+7tuCdt5+ug1JA/Ga7oF
zyFlBGgNXAA0/Ot0TWa8ryaBo+QN0xVWEBbhtNxODVuYEFj7NslSOrM9IX0Du2HkOgqWmz5dm1Xb
n6vKOzPPuU98YqRo2nRxTH6Ia0LEysqZd3m2EjOLqTQtutHJEANZ2jjWcD7CkyLkpYeG9S2RB6Bi
rlacgRpH3QaT1UuulItqb8aNEeJ5/jSnBqfzZH4u69TgsOY/fzQov438czNIKE69rap1Gah2VcAm
8IPoYi1t7E/k4mHKrbZaVdrX1mj7/G/0VUT8PO74zKJNJBOPgle5c565PC++fSeMayyxf55EQ/uZ
Tq3i252TNJMgXMdMyTF6uykVwza+URbp4zYX9dn6Tr5FmMRLaaTAyRI615PIdlO26iTHuSCAsgy9
FsBvRZ30Cn0q5s+VHJHOHGHdubEmwQZWxtxVIH9ReIPbuIrBMxxgChHqNny1C2HyM7pPfhH1njEd
cQOqjpzBEzW6WhqYxrDfSHjaMpQl7t87zU5MdVTMiDWm1suM5R9DLi0auGpBYKEXY7XHs2XAkiTD
NBpignPHurxRHEvUU0qw8t0ZnGPTquZyovcKigqpPMf4/BvS0JX7JXw6KAfKovQmo0RqNk9LeLgY
+tb8sQ5u7zAbjFrFMp/aTs3IJ/fYpotX2vkOQ/eFIWoUYoFO/WRhyyeYtAndIHGelCbHPV/MZHNB
GkN670W7Z3303zcelKAa8arIR98d5F+JN7udcTs+zJCnQpiBK/5GU4/+2O/J724Hf1gA+E1qLAoV
byCZ89b10YRmopSxWXw3NSaFLqVJzajHpLkFDdZny09Jmzzkj5WmXeSS1NP1Yd8Y2NCQ/2GjzBJY
vVY+p4nAkRp7ZO0HLeD4XR/+PFiH3hK+joDmU/w5Kw3qL3gVAgvxQ01xP0aqAMYt4i/5HwH1/OHS
wu+CLAY3zOkJLi+ZmiwMaesP7BQb7Od+drCbh9k0zNVcDH1n6D/9E3qZIZ2JxIvg8WLMLfzDBNvn
jzJhDuS4MgM32yWKSm2L4+3RKb9JNCrmXbPLV/Y/hnC9RtOXipS04BjJOP4+8MJjrBkobw4D1zK7
+uh9Etodi5yWyPs9yxj9bAq5o4QJw1r4d/gB/XrvKdeRA6TOElqIbKAKs4bUvHGJxibiOMg0THM9
+KpbCCIf/EJeukh+bNXuCJsLOC//JGW8jHTUQ8wuL+7ZbvllZKxsB65dH3Rq5eRSEl+Nm+iB4/b2
vEmAOrP4WahDfkzlM9h8C1QLaxVN3Fp4lDh2cpWLq/vgzn0kiq8ATrWT8jZg1rG8tZxPJ6gtIplG
6xb8XAjFMq83h8TTI8IxtiKZHWkCn2CBin2z7moPNb9GS25NaMZezL3GhRkdFxBKoYB8mgfbZUBb
4crESl+/SJA0TkusmtLpEiAF3dMC4upCinqYoc1PkmRZS5h4zSjB/qPe8ZCAhmJq8YrNdFhR/sv0
aO8vtsVuvChIiZ7K8ScBrIBEP+oj9Udpg4BBDpMF5N/ExOGxuwEvfbynCGSBjsv/3q/UoVZzPtVR
x1tpysEglNWHhWvGWsjVGFobvICw9NtZXvKDj05pkH+epi/tDYDgdnuheRLD5IeSGb/Ldls/LZ8i
vpsSPztHYkmsuaslpUTGmhIT5R/ikCm0jOXrARNxaXWA2N7oA0zujNb/ZMT8KlWlKCdNgPRbexg1
xWdZok1nL7HxTSiW4Fk9kcuv7cnLDhny4wgA9LuhZmMfSCBdTqYHKnbHHNBVgrjKGH1BDSu8HnLf
kCIVWP4LNqzMstCiAbOzkvTeh7mQleHzM3q9dCyW2XN6sRcTY4uVusxCNIZYYCgt2xsJBW70OZoe
pzZD3ld4hH9U7+Dp2zqeHfzJU/wC5vzjF8VCSY9VAJpUtCMcPQLZR32CPCSUzsWgOa8Q/qTNo9Zq
fGRdVBOJ9tV/Jnba/wLqnRckr2F1hwORXOi125qE2rayz75hmCvZyuaL60JkTfzUltQgQyF1wyzX
KhUMNeVK6RwouA91nrggG/Ns0TQEOpp7uG3GUX4zkYw3Q+hdswl0AhOrtoUS1rYdqcL59U14nfxM
2CX/jptIqXqjBYyylmfNTMN/9uBcrEVYm+tWGBB9l4G/7U8wvb3X0ozayF543kASb/x+ZXWRT24F
NqZia9upVRH5wWpP4y34Gc9Tg697sYh45BwAPS8vLgZwPKpoYT5kqd8LFD8XEeMpOeTyIbpeKO4d
+iojzWSffXECgfSQ4YJExod7FkVsDCwNK0nkzTPrpyTTgwPkxbbDYVchscqTELMLU/nTXBkRjTot
oYPWLX3lw7kjREXYQsWNZefBgyqS7kNSPu/jsRgm0DZwkYyqJ+NVGbjoupkzirXvSx0AucoTQOk6
YaJd6Kw9A2UINrI4SJZ6hc0xpKZOoWGpg8lpAhGQvQdtC1Ab/V5da4tlS9/L7IhQVC4hOIDmnJ99
x60xMtMlcovR8ltJ7vBauXefKrqXVUWerfjUg9N2GG/GF/JhgaYyFwiTXAtz8aCjZsAMjXRkyAsh
fI4yyaMBXaEQi5VADNBo7A9Wc3ph6/kE53sRqiVnyXAaxK7kVvlb10HbC/A6p0SiNh8KDmoPhXm+
18+/3/C/CCS/T5oIkCtqFIkQWXg9OUqXCmPJa5VvxRkwTnttncneTCI7DEvcOan25WElw/jbhnDV
zEYsnSXC4FW1QN0/NPnmUrmNR/rx5lfsr7zwjzeVlRAqUkbqkiyL5nL2keLajVqT5yCbKv4OEaqd
S4YKjbkQmrl55niefjVSP9MEz7j2NdkMLVD58Bi1t0s1J/lPHD4dky6CudeCcSwJ+0gps4yKD6I7
W44C3MTRqUO70SPoSKdlnEPnLRdiFZ1XeMY+8HbCHuojfj80sDFapefefr+pqEr7Q/NoU1C2S4FZ
GtnADkXc23LARrIqw40+y394A331KL9N/WYfwUJNlgBQtYJUPUKL2vAJ42v3Mx18dCMOu3bUigMM
eSvGDWl/u4XKEvoyiFUICPMd1IsRmWHlMIV3muYlGfYR27SMC6fXiJVCK/S3pkDcxjdnxoodALNh
e35C1ijq4umtefzyeEMNEmue0LA+6XFRrniB5AxZYKd6it5WMKBEtiuNxkvE2+mUlOt0G7i8CiDo
V7eU1C7rFY91tKPLcvyAsRcPHWMMB6Esdl2G4VF9dbP/ODIAHqwj4+kwJCKkxRNfVUn1h/3PW4Mu
VWO6EeTy9qYw/vnorZIAtN91JQ34gzhA5gGKG/hWuDA2nnnTq4iQbSpya7jerLsk1nm6OgIeLRW+
OM8OH3pu0KlzN0Mo6MDZ1N2zi0jAiJPoXa6F0hcFWRL6wMgWMOsdkgC0huiJ0t4UnsMcxEvsSsaM
GT5v4QVu4jdUEmDML6nxynLjtXJXu+Nc6Iuk2PtydsWuatjLzUmdQfEjOP98IuHbS+2454gJUcxW
+0b0BPm/GC89CAbdlR1GBnkGC9U2kzxCEVHn5QnOdl9NMzHvMxtW7kH0cV4F/FHb9uAhsQnsgSsd
hJ613ZPIVp+76r1byiaQ1k5P5WRCS3AFkpwUSuFqyihkKegD/2XuTpVyMJUeW4tgGXe6wKxjR9FQ
9mq0FtmsA5jMR0SZ7z71b+NNjrWnytgV6orC8hM0haNhbVQhuy99whhyeq+qBuiTKUNlSHC6GP23
W7wpoqddUO7vDGsZD7eU+uJZ5ynafML6iID6vX0am+6aKJRVH0NiY+QL6u9ejDZihU2acaEpL+2A
J6a9HPF0DBV56wZ4EeKMPiewzrBIp2mTuEmLhsmjC6y0N3OyMmIq4S7W8xY+/IYWD3le90slMZMC
y75DAFOTO7NREBPBWs5nudP/E2aiOWhg9YhBCg1yoYtJNKJGkdpgs+Ub2rQBzj1ooKTMAaZad830
GCgWXINEe5snTUWhUplkqWlF9cT6NSX3F8qkaGIrMaSgG+vmGGucVKnR7fBuaxVE7x4IahooETOr
bisFIR+6NWwz0OsIusob3g+8Y8qTMjSoK54wKOGbF6cFrCMcr29+kbu8s5bBKEtugBGzxyqE8p9f
Wye223oDEhct0Qcv8KGxloojSWVpkh9cZS1bkmdesexZRT8Ue+jSYbB8wKN/f3rT4bB5XuRgLkNq
5JZiuU3WjFBGJBNz7LIPqmYVTFKiFezqXPsoP50RjWqNiBRZ2oq1GXbx6EbUK+/WWJVSELQFN/Kt
27aJauzsl3KgxiYtety46xvxPVsFPo7GNWRVGH+sWrZLsjkv1JUDIXa+/1fo3v2FNpiZs3U0c8FO
fJYzswbetnxvt0Sxo/ysYeG2b6RrIJINGAMIiRNB7cgevShRG9PTFA5scWrfNpt3Q6cvOLcrK0/5
J3fqrkJvyC8hiGQil7ydBb4ObQjE3iwMUAJDTEgX1kOWLowdtjwVabj6D7/BCTVvUaXhX24AbaLs
dVVtOI0KV0qMSqH8sC6EHl835Nbi6zrYd2SSZUq+mC8iW/LoioRsGQBWQk4rXYUUExRXvNlg28uu
3ucmAeVnelfLFB57xyTDTgH/S06k+ljSGMh7UZ2WJKsGeSDFmFhiIgbNHP266Q3hY7xarYYxyfeq
G9wvULu5dgSSKvBg+Msea2Fxis5L4Ut+7KeUemgBlQ0YQfUrDT0gcEm7OUMm+r1NfuSjXk9wHp3D
JOSTy2Mx+UVdEIFi7WzO9HvBgUtO6qw0Y99UFqJkSN8pNKJU3Ne0YA/LbAONvbAg3VulpLBYFeb7
eVFZIFO1TVCKA8/tWFqCO4sZ4Yfx7zWsN/awHtv5lmoAqnAU195dHxVBSg0wVzNsFqIiza1ptLm+
JMYVNmmdpZavxC7Ch5WpmBX7lWXTF6JuAh7gkvptFqapvczaglJJTWiH7eXBbkv65JC5gXXKXQyp
ing1RmfcDvDA9DL0NPsZH0mA8lWvLLTqdfZ3IVsKJzRBWjQA6gBjEhVjEtRBRXjO4qVmmJCSqrK4
drfO1/iEfX+2+Ff0LAT0GE8OPJ/9ImQ6QT/2dv4j0i98FEm1MHIHYQSrXnbrWADqDqegD0XX9yP3
yVYx21L21vxG49ZElHQTt6E3tZuHh2c0n0XR8LEt7pV+OjJQjfa7dHPrgHjyPcKzhEBlp2sLnhHh
8iHvN1aeI/Qx2aHY5+NY++abBUv8TcS0muqEbaeMKNn4ICjRztPJ/EGDmRj/asTYMX/CZj5MgG1O
XbdjYkHnSf+yAwNiIQf+aKqQAOJUCfvtUkePI9uZZXc1tUfwM1w3AcKNDqz6BOy7cKmKvdwKp3KN
EhERDwEHmM4sYCGS7Mc2iMyOhBhJMpHTQ0X4Jf1+TUe+9DLpQlS0XdzgVIEq5WMJnxc1A7LLt3Rb
uXKcloIlFJdpFhAaisODR7xv8WKJ/Lzunve5uVXpvnX7JcfpQcNqxkfTdLxxJLjTXo7nse2Xsyu8
Q1EyXbQroixuFgweT7B6CmtxrPL3oVdQC/Pl+CEQEllZDmRZLECQDRmIMS2tnBy5VxQ0fTescIaI
4r4RiqBrc68NjwNIpYDhc+BUds2LNkYVjcRI8kACo474HPnnIvh1FUsRd0DpP9wC6d7rQ+lD0h6K
TcM6h4HKDCbUYVyHDQnMxQj4XZ3hMlIWOaGu2M9sU8SoZ92xhanIwbDl2REkLbTKWbTJnvxnDBOO
NaBDPNJ5jo07XiAJ0lN3uX/FYhHoloZyHZQ2Ud+84fe8xL0OUKu5eivrmx6VQuPV7wT7xk765qVR
6xMuxpIDhqneVTqJAeoec4ERdpewerPhiHWr5yO7IxqU7gwRsARUN8E4HRZ0zSdls9yaxVp4I2xU
FYIlcoGMQ1xLCkWMR045LhzunqQEo6ac99p3bB5cdIaAB4ZN8zvVZ1rF1/iQ7nvP2ZUE2G8D65t5
G/bf+jLBL3BbKuWrwWKOSo7u4Zv2eiyGxj4WYRfjE1AY++Jv2r4zzdLj/uiB6qSCVQUPndDNrMMx
+GKmfqGVoYCstduIKt2fb3X4wqf1NYcLf3QqBJ8HDhRctjk1G3oYRkk/2m6gNJyYixbNNJwn8BFT
FJVK2VQKPV7cl/SAbR3qNNlQICkyE0MMJvaWGrDpVQ5L9YaD23xnYoFRw8388zk3QtTw1HXEVX24
jOXVYwXk6fctKVPYXitmuGN123/2yLYAznJI1L6V713BEYPPKz5IkeXHVuaIsIqajU1g7/Mjr8Ar
2EPMcXKFfWGWdHB11ntzyM3/YWQ9chlYSVsTcOUIC6iwvP/t4A1rMZMkQ27koqhtXEZEbiCvLetP
G9WV4nPvsuE+EU6TB4albC2clh78YIcs0dcaNde+r24bYAi6CtdGVxwQkDHotRWgJvtNOTZXr4A8
xKGPEGsxGekh9ZIlA9FFOKlTaxNESNaelxcBwQ/rTFWhHZwSb13z8DvzkR8Pr3WMFGTYMm6DvBzl
nn3XF5kxMHi06NVAfySYklcDIA4xEIrx6uZwY5ngC3U0yWoxMSZqtgS3PuthbBRKFHSQXae9og6g
tpbqzMqusHtgt56cvGj5uKToQgFLOuwR2uv399nt1jjVxDHWGadCNeRigk9MjErvgVTwCN4U2AB/
5D4NShTQPK0/MXq6USSnNVTlXD4wDoL0cejISAidLH5i9iw9sFmYBDbxfX4NCeTWSrK+9xPLf6Q/
J3axzeQO41b4ci/S+m7z5FXY4ffV3G0G0RCSgLjk4Wn3FUr29W2eEqkCybEfMTV2IoSxBy0OXDvH
fyi/64RnJjgwfczPwpjOC2J0aS5DXCiRd6x4FUa5w8BJ/QCRtQAj5VCLHFNx6g67oTYdizMPeUV+
ppSQSODyLq4RelxcCKfLxq9nGdRct7XIxkBaebS7Skyg9w9lKs65DuUk0n5mTCMIcSCVEtoqD23o
yn1rsAlKEDuKewpoJ6ZjABvZeW/kvBTD3MLUL4+ucTm3VNJ98g73KjfWXq/lFxsDqXvoXiY4HWUc
hgJqUyJtUdeLEotXK6b5Z7Jh0oalj8xavhojjUDkNzESMq0DDkjFNtJvi33rjJzngQHoTGvY4LxY
eZ9batoDb+jR9m6Qm5OaxBnkuSWPFT7QF5yZgS65zt8mTzZ84GRWjzX581XnafnKJ0O1daGPoLZq
Np/b1nH8KSKeIX6ihEIg7vlookT5SlKbQn4Y2U2XEs4gHwOx0Abr50xzMV19gf3qgLRmp470rN7q
8DHZSGBx/Rq+bMpkzl8nL2Hs23ZXd5WYwHZ8pUMSYaYOs1bEIuFSCGQ50df2bE8DqvOtAfMOEryg
gFBXE5tzPdBblsNb15WQhdRNZiMhhJWvVZwNqWLSjymsX392Sy3H2VODUiDA2bSljRP7EckqEnkD
fL7Nn277FW1CYlWHb5DprJKo4L+gImCvmAcojJwO4uYnXCrFJ4dsSOAJpq6T0q4h6158eg5O+rYp
yWb3j1D3WZ4tTAqKTfZyiV0uTUosFa2f/dSSg971vHEJ3YU2eUSnUnWLJo7Z5dXWRzkDGZfuQB2d
/ICsEF0/GX3eg+bz04ZHFAPc0VhPoiBezctddUJBk1o3zJ1xe+HAUd4W3A66AuCaJtf7Na6xmajG
fbiGx07Kk7pgWu1Kza7aBa/suwOxXe1/J6gRoYUEC+gMgNGKQBfETHb13SPBE5Tsz8M5E0QWVtFc
xqgRICCuePadgIvOrxmVsES92/5VIQaGWWxDWHHthxFGS63nkY7f2cPU9XdP076iKm9ai+jN1CRM
OIKhiRFerVVtRTvk+cqo1pMi1vmvcI+ngBA6jCIe134q64mDKs0GonY/4DYqs8Zk8KBiHhdwxdYF
1ZQcGywZd2+nPnwlcBZ27KHOqnOOPhenAjgGH5aHhBPQU2yPiOsmWysbM9uryYs340BvSRj65Y4W
5D+0FEfO0Qm8AAOQXUBCKVup3+abaitVm6uZ7cl4nFaL5dIvJxcstHtevNanom5TdG6MEBcBV3yN
Jvc//kDxbG/yOytwyR3DNN8RbLcTZltulpjxQdZ7pAuAG3d21VOMifa+2KevJNsCDsRVO05Wj/QV
XF7FwNgVSdiIlQrKXjhZVHj+l4s6wyJjKwpvRMTDp1htypZ6DmqmD+R66E85ni1deZuA0kWBc2eA
QT0Om/nO3wvfxYyqDD4xZCcc5IJDyz0SJ7OADMHYxJLlZO6b5fWn5htH8WgdrK2B2BBmFRKru5ea
/LnuBmn0G5k8N4IoShMGJVpa6bt9TbtskpwBxtfqQZepFoRKShF847q5mcBLo42p1qrkMZcJ5z7z
2qVolZzvq9MZgMFLvZRoFaSoxEXSeYouUuyB+7jaUH65gZJ/yVvV4I7NrlBTz9CSzgIEf9Pdlb7d
UIdViwvJxpcY1nn8PvYMkPtfR4NBK6Md1p6z5LrfcwXN4hef7F81xrSAHaC4YA0CarVSvPEULXQw
vVjkBOUuTCdMdGrBIVQw4pCiL7dEXjdIZ/6yyv43L9xRz2mvCgVrosB4CC+TlejJ1wvWrpnsFrlQ
tiLg0hxlaqCW/q4sq1JrlCM/rDLwu0iVFcYghma9+Bk2GTKhdd9OIKEJUlS7XPpX0pEFzfGETWvB
qVzxjmscM1+omQHOlSdT/DV4jFmkCoSP3THRilIk6l9nbHXF7aA8XEFXIi5Wy5HyujZ5QOyAf0UU
98CUw8mJ7ghf4qVJY1gvtmskYY+8plUMRQFHoWx9ns+do88H0C0xSve26EIJYUGoMWaFjgKDNAN4
Z1cs7zR33VOtyXcNghzZOp7SfSSrUaxNfX/jfDpIsn3fsSi6wAJe6R1LZ5hUcn0RE6FMH2aRh9xV
gtrv7xmy88hvpSQxQQ8hFu6GfvK54k4B6P+4EeAYjOAOmvmJ3uzdBc9Ri62W+c6OyKlyMbmA3bZK
tF4YR/WlpvYeNCrt/jTPqe1/5aX/9qWKk5JRYx/Wa9NwFpRcOO7n2oKhP7C7s9bD8zV9drdDbi3j
RUmxHlWm9fZqJh1hQByEsHfTL3YZiheTttM6CFVVYWnn6l+r4bXddkRTJrLob7w9Ej0TeH8yZuXt
FuV0stbWDY0RJAOGSfXX+jNaOKYDtGgnvC0eDHFVy0hyfbofSmk04dE96wFItnv4xA80x+9ze5XD
ZZ3/GnEX6m1lNGDp3ICrMVX5TVdvTzKVKdeBhcy8wvYgjOR/WcjGHqb6cyu1vB9iLcMqS4rx0Lcg
44UHZbozLotOkdt6FseaaS44i7yp+IcjRbgOXeQUj25PEbg8sNeFywJZOmbcq6MlIgvKKw6ZJrmE
fXPe6H3ajBuoDRVc7Ra6L4cCcG7PTMC+wra8FcKOQ7KBHB1ICC499CRfL4p8/eEA4jB6n6zIDfhi
/szNviKlv+7GmXKLRvmGjUlsJLhHHU1GYvqYg6xViJgQKQTXt9U2EHJgZOSPR0WPgHlhUoZqvlaJ
9UGogdfbyOqXmXdLLswzmA8UOdQSrvd4xWywzU2D6GEak8Y2BH5Jm5FIQP/cnseKbqHW11/pLrm7
JHgvatXuS1rkNpAIRS3wn9I65Q0zBxV3P7fc2QbC0kF7BIPLCOP1QVjpGjecCxN1BeA50oj3RJ3x
N+RRI13qkjhvH10xt3zkbFhwDGDyouNHHDB2jg8+cSg3sBqdz34LZn/2yboLhpLSfoj43vqtVJjE
48OFqVlSz8IHY46oyCNKKwqGEikqxEjoElzPXbgCYuUcip74m6zzxJc3mSgSlwcvZztr2bPfkpOt
xpXl/bZ6NcpaQV+kUamlcMZSK+B4qb4+V8jW2LjDVLoCk5Na4LNAzhhvU5N6iVRVqVCf8sAf2mAx
Gk3uGccG9wjPEcup4ts6i9nDXs75Upzv4+mgpF58fxY0gcl/NKlUP6RutoYcx1x5uRmXf878gESZ
Ex2q5JHcCUg8j91QL3K+SD8F7XhLr67Ff0OGl7cDsOqDcWtMgwE07bvB4XdxBTPr5PBIsGpYSG8B
uF1Yx6s697Hhzuq0mgot1TZv/rK1OXnAbkyY9StCKcDAddQv53P8iMVk/4PndEo6r3eV1mdawXTW
myHaN6oQ/l5ndt9Bepcgjgt875kSTDBtHkSmR8xY0A9klVth8ZIUjV/+YnDN4tuk5wmz08NBKxfY
GkiCuR3C4vjZtLipYMreHFK4s5Bw64POGykSqoXChdBffq50oYXl/2lC1SSvRbvG+RhtznAUIm78
PDzIVqwHzBYP4In0mdiOEbIbOBodithvch8fkSzAWY5Gnn56QEExZwPGaQWXDIe11/ZLtzUdZKRn
I9N8t3xjT17eHXy1VbjrtikFnZxr11qrW64Oo0FS5oJy/IuIEcXVGCSx9c3kGT2mvdMZjThHnGBW
qnvz8li+4OO4gfyEelQzFdBJJbtI6yo5KLvcPUUXWpK4Ycr03zIrdR8l642ZuxhtYaNWvAUYUk+S
IUMAvJ9+X+n/HHe71xV1KoO4+afoCrAvzNU2pxvQHO7iKIe6IIjVcKDGtGmfb7V9qlMsuP0gkPVq
q6Y6JCpkVgT6NdikUG7exmwxCUqsrjQIvCQ4hvw6S++MTHl33F8+5ixL4vM7IwXEhSU9wZFLnBpO
WEWrTqnX5h4e01f18zg5L+EyxjayYM43yCU1UM/VdiwzLgQJxlae1EBbpwNjEpXf9RsLPZJVJ4Lv
q2IuroH2vgtbQBuQ0jdZFny1/Kkavs4hlhZ2Ire1ia1fh8M8dU9ArgIlvdPMDXyArbOzycqbz8IS
fpBc2J4EXQ+4kHkTlbO/WIXqaMq+/lsycNgjAS/7IyOaNmXQ7OrhnFEcIv8OiTsUZHVOvzxkhciI
UcnVtcVUtLPMx2V+iG7i8lmx7KsYsQyGQB6cptQ7iOctAgwP8v939Tw7QWGmFzZ5uzXV6XdU8mNY
lMwaq6T20L9hDqY8xgQ+/aRe3MXTCO9I+ZbPA1K29/tGhksY/wB9qiu0qHo6AB+S/A5ALb2rNUSb
RoaDW3YKOU+SdqKYSJpnzeaJSKZYO/zFEcfWSNKsYgxx395aHSVW6l0JMDis3J7BHf8U+DrVQg7E
dIUhc8hicGLdX7wM8wlfR5rvzn3GiDVkdcbITLGV72guQb3sOnwGYzR20fBOtTdl814HJXDeNiOA
uf3fvKoT+0FJO9z5CNZRQH9+VtsMf/xSyve69r5hGuJ3xJcPUBtRA7Ljb2w5AeHXzlMlzgUvH735
/lfnrpNo8tvdt5r2I2jh1CYr7cnTGc3A44vLcqlu+6b9NM7FOTbUbLUNMpNK1IHD3k16lMaRL+C3
mHKHiSuDECdm0l30zcGmnsNZRo1KEykaPf77vulaJEHEB5XaT4J4BxaEQ+QEKaq+fG25SmRNnIzO
hXPGXJ0y5Oj0wMQDvzM8142cYBzpGPNqUFYMd1fz/dtFUZt85mqeldM0mqWtCvFNjhrGaklgr0kp
YuOI+K5qnFMoT581I0unPFkSc/2GjodZ/qqaJxkXUxd2sF8wr1l0Cwb5fPVTy+vAR2XCNwHKEJI0
JHZRwm8S5OUspH5QjjJB469M3JqjwYDowU+PvhqZ2hd5Yt29OK/iW11jqombiQQEvZ9QmpHheq6a
Tar6798ITH8OQEfOP3vZU5FzYzEeQgpk8quPh2i8krq/XbDYRAcLaK0TCWZ+xLqMLY6m/xwqUqXt
5s/pnB7bpBgbp9gDW/jmSgPLXEZMH6QOchPxn1Ng+ySl7nEnT4YtOIYuw/NmT7n0lNFZexGSpRpw
UOJr6rD1XyxthVwhAJAvAG9XDIi5mtk/2DrJwOvNGYvTYgPGH5KnfJw3bIqs5HH2ixoMt4vlMV2a
fH+zqMQm3Iis/9LobJTnuwh2d0uDyPnPL4Nodf1w5KempZPLJJxRO7R3PsseS6WKx5GTeQ+I65H4
4FCElK35rEYKOA3uULXPIQrcseNgYlE73UFp8/xzW/sr2xUtbl3fnGF/Ww/9ynn/El4lHliq6Xpj
ga5eGZgHI1E2tY1WN0B95tq8I3anEm1gCH2bLZG2NxFzJ8ipg6HHS+YSvRtLGGM0MfM3drDNCD45
nwG92XzV39dd8aeoKQfzpBtuHSbXJbmBGfSoqCKOOWN7TdHcMae0sqyw495KYkccAqpCLuEgEc+K
AQ7VXDzY/o/90R1gJ1bsUSrwkkYvrdHzcZkRQUMKEVDRQit4TLgRBKYqv466712Vw5p5LMT+nWgf
2hB9O7Et2+wrPdyyZtblGNITUoTLx4u+HZzvBYsqDxy4dP3jQt9GHCAPIW0Gt75I2Zv0AgMpa/Z6
4uY+p3HcoXUGI/eJSA9h+qLZ3S9irt9gY+QTdPp382aC0EYDcLPD6vU255k2PZj1DX8c7tEKKiJH
WNdfREJigmIwujD7wqUTWAd1RGLDMxlJF6aYNJCOg/mxQrotI+QboNOsrKr+/L4DVW2kp6swyz3m
6LaBu53+qTkfvQ8t1NhnxVb/bmxDcOUW5qJOKC7J8NIvycgPl6J+Uau4iHQ/NED8Sn5CaX9QbsZj
5tB8qwQskS7+AYG4a1FvgiShBl8H0DOzZIzB6r5dpAZhbL4O0f7tzPG1uSKcSoSzpVWgVYA9Czj1
GOBzeeAwipWmzehptPy6/X7vYKTaJLva0lG5QjF1acvw3zEcwFybrvUfSmKu3mlh1tfYUlYk6eqQ
PSRWVmkbiVuE1JFJYX/4nLQXIy+13ksRFQv5kItHCgGvENrxDPIwk9kReocU1p5WM9dsrtQ2X134
BCDj8hOUpajeIAEga2fwRhJBHIrcUdfE0qDw8IGi0R4Sf+f/kb+0O0iF+9ZBpSL/Onc9MCR71hq3
9sdabXzpBio+bqyqSlbuYwxsZkWaOUug65JP7+nuM9SPWDExZi3jJtla+w/WP654KDsRujbZY3fi
Z/7u9tJl2jgleHELKA3QG5G04o4r7cloDMf8ME2CxrKoAiVowtFQY4Lu+ZEKaUPyqWu6YKVFkWSX
qKRO2Y7gCqZOV7IYKziMSPLK+jDW6p4h2NFRLlXYLHzXFXPjaFkw41Qn95ulPC6OCe5OrqkWG92+
bLMQWrNGm6Rlt/Ph4q4Q8rvYDbB22JorU5j2Z6awyLC94M+qgqZfMe57QV6hkVA9wcDiKDYhxSmR
CFSn0ZUV2dFTAHLrJoewWuKOrwuiQsC5GdlHEOVxrkhMHt7dF1ru22Ntyv4zi+CEFWKeP/F3mw5c
pnzInY1NuiC6P2Ka5oLAtypliFtpvKoWKYLyz/GxcHdO6G6/LGCZaKn0hqxZzk7xD6yuv2EWGPLw
Nf7O2sP98ik7Ly6vQvs6E+48PQfxpy6kE65u14h2lWleASW55QXrY4MOOzgPTSESGQNWyINWH6XR
bZ/xJF539oCBTcb4qVnTCkKTHfeoj5FFhbrsqZRSc4/wvHbPWt+wHjeg2KRi8hGOAlLzBzXmG1K8
Ltiq20j0HVOZOu2lKQ0NQuFrcBZIumFCr5A0la4Dp+o72hurhRQwyS3yIXyTpj8aAx5t9aV+akE7
OvABtrkP0OOlc394ZiirVLAaaGbW4hmYnZXsF/nyopTndHQBHs+nbhfukIkVeusM+KgnhxuOLbW9
npb5ImXmG25uWsIyzVK3xgqJUQIDZt+mBPBMn3GosWeAgBLT7QAL1klFVGaxNvD7Phr89bKErFFv
PUkx76XirNpRm3nFoWNdyYli5BgCYj5s7Y5LsaPcGGoVhO35B7bTjumJ9y7QRiVZJj0YSm6hp8Eo
cs17BwgFoc6aMwEK/VwfL6y03h8ppdqrR6ETdRnM6g7r2qDAf71OIPWxnKbHFc9x640ZLn6FTM3y
IRyBSZrz44J34DcZ6dgbxQtO3VI3xMTTm7aULx5hQnY65nP2TjB9qxURSFOL9lItXEpeKo/upsTh
U3+lxDq4m5BTp1NiIHsC92CyZ79CPaiTil4F+5+jA2QXEHll517hdtvVDC3eBMGzWC2/Rt4EspAL
SVpkrOXeH4UvLogYyKKvwJ7QJZYosisJW6wimHLciCWAkSkmGodLXHCiNmABB2F+txyxgG7PeKia
grbpHqrKJeFMHOMs2EHaJLMneJZ+CBoHtWUGvrQTLWOyMZmq4Nedn4Cm15yq70tafMjgoK0XO4AB
5y8j53ravU58YVCJHCPJKuKfIvMiXSKQW2zV8SaRRHAka9U+n1TpL19d/QyQy8GAuVdT0yWoX0GT
X66t5VdwiJYLhcIaWOkPg1BMnQPUiHu3oav0y/1Qy5OkqeADYfc69En0O83Lsb80IspvoGcSqiFW
/a5Er6brexjxnoJcD7KDI71UIRV1P9QzarZCnk0QVzkz8IDNP9Sw4ZxjO85HVMXEXIRKemlxj+js
n1ZrTfqSOkeGZBNV+6pMmLkSUvRKGnlfoqv0yLjNrDt805vqS3PEWd7XB1O4LKwKVU+COpcsQDrE
a+S6zHF/NtZOVcWsgj5p1GZHKolctnINHfDgeJ5P//h7WDjconhWf/OK6PQLPKBAz6eldsNrnqbO
ec/rRqOLx69mEiW4jEr93keDXgjzb2vyPrDvESOx+5RQBXXFISzffe7NoNN3u8H+UW7z6XE2FhJJ
J9x/R5q+xAKQfHR40ipmZLBj6/LTC8I5Itjsr+OZs/EVKmASC0kxF9GSeOIT2tfHsp4kOm2xADR9
DYH/PAN+mn5Sm7YV/RJrstQJRQ9KmtHeh+xv6ef5VU/ImFGAUj1RjLJGcpHA/jnUWT2kGvALFcXo
BR63Kwtiw+EwaIEEAxhEnDnSpdd8NaLq6zJcntvP8WKM9GLDAlKdUxqvk46iZjOn9PvYbF6j/SKK
FGLzSvFfn2SNus8WUB8VcINLekWPpGDYkjuytCmK4wPBCwXC8pAuYsRIw/G+QRVow+pd3UB+GMSF
MLHpnplCPfhy4CpZdwsT4KjZ9aanFlQkKDGakggqUr27tVlwNgl0pZx5M04VSiRHftxwgCBHp/1K
lkR1IPyEC9N3B9gfy7ujkGf/mig6xVudylMjJiWEbnCgyLEpzM4Kn6mk8RXfzmxH+I/VqGsf2SJP
lUwxf6DkKmjwxaZaPWR4uIco/BBaRe/c5xlfnGa7eW0/Q5EqtHVpgNfhd91wuNSS45QcoqHwMo4P
5dS8sbM/mdzaI4eFTyQ9x+K2KS88rTBMqY9MKGsTbVaxA/q2KsVTPsnp6NjlGSs6Wotr4O0dPsCr
GCfde8NF5KCfGacOcWjXRT26VLiZEGrT9tk6l3hyhGYfoIm60vQxqH02/bq2FLOKCRjzXFaBOcHQ
SyBV07vU5gcYeKbpGUrpLAlh9vaE6RX8W7rqjCzpnNm6AO5+BVDMjSoUWq++1XLobzPUS6DoUGgi
c8aVVUnT1FyyUtAMcJYdOrZAPWHreiCafvzXnyNmlTPIHXHvsGiRGJcSBykMGRDUP8Owe2ed3i+A
7VVPLduhF9ztDFOW771E3hmTB2njpN+PdgI4vOlFF7gaIH4mxlrpWEjADVBckUjaUk3rJPQBkRgt
/gmDEb1Y81BhP2WhXQgNGYYPjCBWH3wldiXSSO/s0+chs63b0pzfzhLs6f+AXnbR4TRzXyWU3lVQ
u0BElDDlqD4YbThtJxwPdMasOxsyk5t/BBhUSkFV2L1i2WUxyxiXen7fWCOSMlVJV9m+UK27EAv2
z7cLLPBR7JWWViFgiBA2pe3CqzLz4PJVgaVIn9iH0WuLhWBC49nOHtbOW7LWujVqdNXrWV4vj0V8
JkC/ahg3HVsNgTCZPmmLF8ek8AEORPkqpQpv8jW+4tb8vKcawZJkm8KETUrHbuh57o5Pkf2oQcwg
1J4VS7ixO6zdl9Hngumpq7OuKd+4Pk+Ra9PEDC3y8aF0uFmOMRUE5E8HbkywLCY5TRSKr6vrvo/+
jPQICHgebV1dKzUujBl72T7tC23ftp15iJTWGWOK4g1aIBDR8ggJtKYBAo6voldzBXJHsAHA17WT
JUwxAJHOOkvZLj0pH5jyPlNcog/qWC1w3eqEC73sM9LLF9I0l31TXGsVNFG2zujVsku8X3zGq05W
xecKjoMgiH4/b9NGUxDOwwRa/AP7KrQUSwjxFWm59n8XtYxAi7sR6eNyi56BZH+S8OmLBYZ0zTGc
IdkDYnUocpv9RZzyMlEEbGGWA35QvB1YJeBwcTLjtTxiAcNnBMoU/Jr5WAnE9jEytiq6IZXBm+w4
ikfhXRlGb9n9bkmktnKKB+mgvWHIdgk5mjIS3g2OuT+qJD2LPv1ejq0tKzMbtrLdqJ4+TZ1na0ut
tDW+snIuORvkGH155zKE2ShBKLYZhM1TrQTvSlTuUy2vvzUpAdqn53meDw5VsAQcPLtwYAmHJ6oz
VtEhTHuB8+EpP0ZF9EDxrl5o8qmgcnS5Eg0qipwRZ9AgXRae4kbDFmBDaxe4N5hw2jaPIaXtWq1w
7HaCyODY3E1qzAgQYrToxa2+WFGnySg62UnfKI5CHJbWjdZ/NuILaesC5hro2PYRIbkl/LYD/E/z
CEci3G/T/9RcYzhuY5WFG34xrHHv2PbPb1/e31BuBq+VcrxZUlwoilr7ytk5CACjwgFy282ExwXy
g3XUIoCe/Sv3XrHB9tfTEy5lHDfSKKXGoQZP2fPm3pE5UevJNTquBqLSw4d/ees/Wl5Sfjnft6ih
W7SgNyPqa9m0C+UNZyzX/BtoMdr4VF7ePwJ1Uuqak0DnSYeN/jywkqhNXm7o+KrfV3V8aPfIM0nK
aMChvE0NH/hPnBrJUsP7puFoaWfd0kuuOfzHzWedwqjrFWTzDcWvXDWWUng0oj8YKqP5/gt5+ucb
WoSh6gN9NMZrHQZ8muycYfdCj1PLgIvzNlLMGDNIhn5FDumQsdhcS8byRxsZsW5L638UIevQKU8T
RG1c0rN4duRVpQXyyti0Zav0yr4Q9xitaLoZEMURyF88wg8FaHNAx7hq9/2VHNnamue2uKDRrEuX
to9glPv8vMKZRmYJxv9oMbK2qAhcVbD04wkZMA212TpwFeh0mOY8TqcXNROSL+kBUVdjWSGBVkWF
QpvIO9/7gqhLIoaIb0N21tqEOFsDeluNCLGFv8YQiqjygNT2M0CNZUbLhZa4KqzVsEuVFSY5UdUt
0evd7BtqziNHSkMeJW/HGOb8/CZOIx3rPz+mt3UtPIJbKXZil5JF5pupFOTpCqA4tCRtRnmO+Ql2
Npb5D9OyeWN2N1lODDPk2UucUcfIcLpRog8hgz78qbwMRVvVRJPd25LUpUeWDFxPYFvZZM3VLpi0
7It1zYrGZhUSDMqXxnzyroDY3/EeGkAhBWy48GF51HM4RVhQzqpeuK609WL2KOVvCciSg1FHEDMP
V/ARPrYu1m1HoBz2VQvw5tvb2SIHw+mCm7FtQ+RcMmHJ/uAKThYecpwvVFsjH/KiUO737q//u0ub
BNMMzQtuF2tIKYvg99q2pScPCJQr/Ccd6bSGocT58bFPnlnuS0jFJp/8y+hp/vHgVxtZOoAEzXAF
/RfKX7r/hvCjJwyshozYAxWjRrpszmxnCr8MD8904lhwhRuI9ArO/PcaoEmJP9pe7mtGuwt9OD4M
Q0yOnvsjdCpru2NJBzKvkkPbBPnl5RdUU6iMw+Idw3zVtyx4e1HrpPCpWV2noaFoFHuIFhHWrPJy
yxWsmVyI2wrw2arkpLuC22UiXpP01p71J3uE393+9rWtmOcGshlDBHQwgXT0SZjJcOYG75/ElfUe
Zi+Muf04VRwqmJ8aRJx7rWrssPJ7y/Dr+JOnpZfgUjZWuA2i8AHl3BiPgctUVK2yKiMqGN0ELq/V
DIES1fHZSpku/W6N68a6uTK2EskK5RTBk4dnqc31moswqL7Sm1szKhPgoT6khaoJfh9bpPnFVaWo
Z7jyrYRNdxKxXKEYsWIMxDV+uypR7L7L+qFzD+PnoHj/53J+QqgrviMtv//8IDUvL6nCGPnsS4Or
34SA746wOoUu95xuRjR0WT5uzXihg08YbjBEV/cGZqKRqBFLBR0iXWNwNzUDf5nPbWDhxyGGlg4I
poHuZPJBix8ivOBTtP5PGKh+QyK16n+448M2S9pQkr46b9aevZVPSF8Urxs72bzZagI7RK0NvO2a
b3RJ6VBdEDPgtyRvtcewBObFvFeDvItn76sNmtNH/RNPUc+0AjZ91h7FTkcMWRKt0d4N0mrzWibr
AW0OlKUYqzBBvo79X2+KHoJ6atkXft3HE8NyAhkoYTUaBQT7VH24LZyPym8l+KOth59tTR1+SPZW
6j0s4ZAtpsHxO+P4SqO+S3iR5j/vCaM+tiPQnGpp0tYbdbXf4LGYwwSgme8ayg/jJdmQt299ZifZ
yVzlu6b1zLv/Js83IHVaqRujUvjSIWEa/wwj9G5FSs1jkCmEvzhozUwHUNtY1c+E6G5H4HVLLBSc
yViVrFEPA7e3ucNIlC1pQ0Rt8xKhyRVxcT0FivmxXwxjdQSsPP0tGz68iEBHrkwcC3TmOp9GvF9D
E4nu4L/f5JkKWq1jopRGeS3lOUrsvEDonoNqinIgMbYTuuUULxFfdoNZQ1GzJVmY7Ooow/rCb4w5
Er0ewsn9uWzV4Fu7umxgMbgm/JUnBnA4RkNcW58zCz1fPfZ+5goZsNtC8WuGDxGgG6Oj2cD5IxgI
JiHILcCspMdLUrU8LRKGoIVW0HTVy9TGJBAb5lsUGaMsKi6GHFQ5Ct6qKNWESjZRXNNCDTuxnmPq
ZP/LV952qetVrlHucCKyuTdfJZgmFPgLcdO0alrI8R3IqYlOAwOWhV+guQThi3Qp6UFapmptEheO
Kvjs2s+PKvkoKMOgK9msRobiseTMUNrdN2mWEJbKWBhqD/DDgEUijaRWzsW2rswrwz/Rp35B1345
oVp+zgTmDeHykSUzc77GgouCeQfgw1B9HZ4UEIwgY+B5YfSjkqgRs1Xe2UdbW4ds21BL1PX2WiDn
ZKcfhdhzJetEww5ysHSqcNkA/FFx8X8h0fx5xSOSlxIaOjwy926mBXauD0ejAcfSb+5R8CNhUZxH
1T7hsWNxJn2jzwQDE2iglVfn71OC8ltLZQmy6OOFNgEo6nrm/17y2lLFHGrnOUiQOh0JW7FBcDi0
nT5v1bD+41XZJXGWKKwT7k92pS9rwk1ohlI8wKcexxgo96boTKgn35/HkyvGUawpM6ARCuCx4Jk7
i/G/Hfd3TpLktu5cuX5TxC+uHf0h75M+FVugLJpScq+7DeEgM7xL9wCcxhDNh/r/2KZfFW9+LS4S
2T+OnFA+1ksQK/rl90C+fhsPYzZQn6vVc8OCszy2wXKJBzucB0SCfbk9LD+qgiyiZkS9hD0psvsP
cGkoBvfnSzJbHGilqxzAVSos/qdQTjXUqeljoOYMon1qVXjoSHSQEymFlVNW5Jt/tHy/ffamwtKW
2SNigqJ7h8PEgMNDHD3d0MRSW7J1T4xg5OjBFSViAyHTMTtp+hkgQ3mc74chH/oZgGtAwUE1hm27
ETo39tcCi8ZOTJ8LHiWKS3KZUQSApR4pVOuFM1K0KOBweMb5rOOCKOtB6FVU2T4OkWv1+ulmW4B+
RVzvTIS+GfIRppXIv4r4yQ8ndBB5Yo7mA8Ssm5CDIB+0nCxhrwLLJIeSBomE5/ulBi53p4tT1g2E
BP//4J+PPG/Ga9HEeNnnS8N9UTTaVVo1Maw2WDZW5TnPwl/R3OjDQOgMHczYitDYcZ5/m632nWhM
7KKaP5K7hozLj0CSeNyNEYA3GiqgITysr2cia3XhY9rRUE+oJScTlpmPSo+b10pixuHcQLnjkYHu
3Z2RxHUYaHEkdzW22QMSUf4K2fMm44WOEkDMlUh00LB+PkJ0qf4pIDZe5O5V3cYFYVwyk6ytrDXe
OIQMqvQMYazg99/L4w9fNu7Gp01uEhkllxDUx+UZf6UBRmNfImGX4FQ7jbXafz9+CgLGX8c3GZWW
tUkkIb0XY87gdrlsnCIv9SF8fF82qXW18WPBSRry6NWqb+gsQ0YTdNKxaqURxhGKOky0MphxRvZT
Nf2ejVN9BI5/i8UVaU3XJ+Z9voOoW57i+g6HULLfKm9dLlGFQkeiD80KIwjmny6dptzDgD29tEni
MXe+58vkGIrM8EtJ6LKRFN90NmX/LbcexYeEL1ILZiCQIb1DXhi2yJil6OvxmQ7GgpdHjGX0TNip
QW7pnNAHJU5ZiwM9sffbmVegJeIMLg2MOE/vL+OwwbDEaarQIzpwQ+ZCOZaPBsyenNXyFsKoB/BO
3LcEEg0qvfwYsvOgDO6bNv16o/uX/KZNIc3+D+d0zVm6QeDhnSbp92ESgth813p6RXJDtL5okqCv
ee540oWvEAXh1ULIbWesBHOcciFaAdwKcq4vcAIduDqmJFnNbwAGAiQp8eCRDOxQ/3yv1zxnemE9
zP020JGThtLxjGwnq0ok/9ZGOr5ptp6d07bbpyp8aJcEeT7dwbStinoVbx/v3DN16DtQyun/3cbD
oUJ4/wRKeffZxTB3vk16GBdoJlkolFaz/drboLXDnIAM4y7bGIq5dUsQ7Hqw/fDdJDxXPAhyiWvh
S7BvFwxVX2KnF7btE2wcv9DPTe9sYLeIXvKV20Jxfcm4+6xK3fht2EyAgQtinFel0HYwxy5cASd6
8u63i2kjTfaFBRlO+bsgLz0sYq+Iod65qFeNRLCp28cpRpND0+PBUuitZ/9XCBfeTtmFovBI62pI
DOOSuVIAHEptMvrtM00ADbYrDRCvSa4seeqTNQyZAkZA2JCTKJBQ34fyaQ9Qm3Yw6gcIADy1m1Nq
kPYVVrqEJbQM5dc8yNY52pCk7eHboWRVpQ5a2Wa/i2ZIBCusHwF9UifWSZUOkQszbzYUhDc58ypC
jt1VRxmykJ8xNfW8mnvB4SEuNYdDmg+pzgyb4+fCNK2HveZp2AVUIuta0bTIEUV+AgfvjOPWDi54
n/j0MYr7LYaZrjucMAHvkv+faWa1Arv1RhhMvcLjx7h2MeSASjE7yJEDK8rR5TjHB9uXyXXxaJm1
XLcJv0noD6UoJVMLiBzDjjyMtHJkyLknPgBKcJq4WquvWLGnzpyQk53KRrhjT9AVut1ynAL9yTc7
ayKXoGEDljxcrpxJ4tQblZwYqROtflXTqFem9j/iOzwjIxbvIr/mT0Y0J+Fqen8IkQ2RQRhdMoEM
3jlFB9mKnvGDH7g2cQPP2lWHiWQwuQimX3HOgp1Y37z6L4ag/LSkTFp4PI0HzXh8o3GPtTSZyFCu
lzXuiU+kOjkU9IwReiWcxvdX1VGMi1XuEPID0clBAfWRgzzhQisNKWjYys8e/XgPIdeIWpGLSpS3
6QIvlPVIYx8kqCfvBrxJc512BEvdAVU7Jba4QoJ1Xv3rIgAFuDR6P0HrLJcUl3/ZrRpkl/eI2MIe
3eaNCWszPled0OYvD+e5uYOUJoVxXxTlMoGFdD5/YYnUIkoyjQocInOFYQU/BhrYtbQgCIcHHPjV
eOqgfvUIyZRvsKHMXPQlKCTx7tPhKomSW5sRawEdLkpdyinHXkXeG5C0qWuis5rqtmCJdA6vcy5C
AzSVsY19SqA4aGfxUUtZdU/4XXzM3OZPXcUptI4ThAUMjeBkbMWZcKywnJBVvEx04ZHoK82OcZXA
GIyDnbhFBoiT5AClgJFZb/SSYkDUk1E5tLJkKcupgFVhCVCiFweQnnYEvlFmtOIo3zogL7wbWYos
kydyrI7aVN7MogGWhfy170JfzYXZoaVkYPk9IFwp1mOIsLSx77kwiA81lAcfKde+psGG72r7Loqg
Kbpkwyo6eSuorBjLf50fQMgvMLAlwLNLxY/eC2ka+j71p0gkW1dn7E+kzn4n7xxzPVcKqdWVpPl/
QCXJCFCdV3zFzr2ALTKrhnw9ojh5sw4Qh0VRt4aGX5oaFJ1EwxWqKHSY2tDgpGxXnwQ/3D2Z5b4h
lAUow257j69yUUJUoEpLJ+U6XnIRyzc9vx8Wb5fVlpEB8ezVfgYhkqIg7tA+tUdd1XC4PiVg7lMC
9Ph/rLi961a7oFQdKs04+eymA3pOfblPLY1V3A/OR8O5J83TX2EHoj3qWPOyULCLCvRfXuBq3cGX
d+nfcCtZUAemqN/yYl1l1JyUVaiH9UaPW6KIf6sF5RudaZ9F2yPykKnXVoVp4GOoRo0Uqf1wC6RL
3qMw7OG5mC21JNliuDt9DacwE9lfBum4YDtIo8lgSOb9iO+wGy0tTRTI5kHVKSgrm0tHJ4gtUr+8
atnbuvTvabk3qi0YtCkZPmOgDGTe0EhmjwZUcGiZ+dMjx78NtckhMZuYUAl2RnpM34gQaOb5Es7I
hy6Mk5vnxomsJEBCIQBnwbKzQSLkUqJ+Y11oLyfyfb879m+TNxc70v/KfjvzPbINRiwsOvCEFddv
9MnXIIkZEUnMWtH0uChrO97Bm1fhpJhkKhmvOfuLFiSc3N8ttenbenn6462UHvoy1v0NK23kzT5D
Ei4HPN07ikqdDENUrYFWLh/GRPyh94zQN9iAyiGlWJch9/mX9C7kCZrXif0kGaULxZtt3WjvUauF
RoipkaZsiK1q1uIyfFi+wwcVQGT77nJ0iq+Ot5pN8BCLuOV971qe4RdKJBfsnniGd9OO/rLosigj
AJe0ypFZkz6hgBT3Xvz7VBsyBLodivprOTyJi4TMBkjooe3S0NWXfkE7rlQONMbOzf5fTBL4tpDL
MQnY6CncCl+E/w4l1bI2rxZICYnX1wOM0pX5QQx42sF8V3O9uuR+MGMkLHNkR/m4+3Wcgud7g7x4
VdC5hyIIZTWG6pKiIZ/GANzSP6ecHc0wUR+yeNtWQGfPowv5/NA/Mpi18MyE1ZUdNtWDCruZ8Vhv
2RyYIUfB+C0dUwPSwhoUSiMbuxyLoqywCtB6hyzVFHnA6K/h8J0rBVtbuNf9AdKJ6tFjZV2sP/+n
UZhwZcEU61VoJARMSvn5gBY9PN6aBEBRYgz3KolyV10aU7hLk1c8wGKVQwvea5sQRFxEvtkwx2A0
H51Id1yH9fnVzFc28RG2w8mQNLA508tvuyjxHkII0lb0fiGYemaH+rLlFKmBrDcUufXfJa1RIMuI
vJ9OCQUXYc+uAkTfFUPhXn6W0ueXC0Pwt3JGxr3gv6TH1kSc4mG3G7xRTbOnwQ8EWdPNCwYKumwj
/QdKo+fK9WjEor1qDSMnYh2Uyu8AdFLrOSGESlyvpKX+bruKLHYOAMWzLBwDHXO65lSZ0oF43uNa
In0WVBOeHZ0eaocGXR7kEsplnD6h2I8FcVn+sz7NgN0KmNcF1/BkzjrxjFO/Ia6/iSUT6pT+19/Y
a13OD4D/N/fTv9yq0WP+8w/TX+57KsleJVgAJZDiQNF/hte9OBfZ3wL2ue6tAvk16JDn7zE9ZtmW
FVIchMBy3k0U7q+rl1HKh5zZevtz/gRLsDnG0N1/00lq/IFN75bYuOOa3JvBwDQAt3qzQI2DVCzT
QQq585juMyJ21oGF4wQ8CF+tGGD2Z1pzk0Kcszg+cDpZ3nyMlQx00TdpzoziRoki01GWxkgAvBan
GMJbupyibbGkZJ5iJLV5+AawfuH2S4vYOgmrOBRJ+fHTAOSh1qzSC6MOR4SINAJlSMXblr/42env
id1LTm5x7agLIdKGhkKX186DEZKAvp7ufsp1rvYci2QmJDT9Rg/Qy9N+o/MDYm75Uvu8WKAd01vt
PIK+fUeTjdxKCQDkQVO6841rGnxO42SgcIIdn616jg55ENfJD1kaynlWFOI0FwtiRkJ5CtXYwDzn
MzxLY8YaLXmpnt+fCe3TsXaxfCVU/Ds+HMUdhzDJg26hXxynpbfuBHAzZrd1/e5Atnf6hI7Z6gkG
yE1wVszlIUkOyN30k8hBwaAchnZyn+sNiUd7gCcMnoasviE+nzZeOmJQeMjjnyQAng6w3L4UDe/U
IgZsCUjt2DsRBUxvYuAWV5Sv+WGhOMNdXdhz8umyqbDjwxKB1gf1r1jknioslmPAIJxETxPTRlY2
HVP8+kaOXkMDR5UVFmEl5GPJcQwXf3t1H6loXx1ujlYVFytbUZv0O7QNu4sXMVva6vvxFoS3V200
O7YwZ/1Lj4tT2pHVBTKRNrSAQhpOPBGWspOMABU+3fQAYarJDU5lbjUU/lkW9F4yQcSxpuud3sVs
2pthUEbZM24nelNTDcaL+g9GRBW7olts0Wqhr1Y+7h/jqYBqanltAv3+u+zjLzmbjEOCIzFdbJ/3
wJRaSakpDp0tvLPhrq3ESAr0eXrz23rUTQB7Zb7aMS43zaFK6AtqX6v/ryRqy5NON9a3U2P+zxF3
aDgrANxjy+YvA0AUTQ99xAsoukUV8poljWUtT6rRkOEMvgNP32KDhrDvumNa5iEwbqKsFUavBc9T
2jP0nYVb+2DyigjMp+d7gmFJNy7S2fdaUldzygMuie0xgnJIm80qLgV5rlmffZYmQP2kR57XzmFn
8tQIldG1sx9LHYjzGB9KaM4ajZopVnCq42OkdBJt2JNLbLuUlsX6QfsNgJiQUtf9h+lEAey5eYiW
lKYlNYb0gpHAgtqLnwHm5oixAI0bj2+/XdcCzVyE2NL5XjsoedyBa8tFy0TTcSmdspixapMnTgPL
GiZSztGNE58/eIAkkQGvAkAmFKbYV5piX+kbjBDqm0NxUn1Uynn1x6J2SJYIvAXtNps+c7e9v9dU
5nCAnR8LfG15hxV5TtDyA5++cU5ZJ9G6p45q57B3D+Pje1H5/KlSr15nvUk7nWXRo5sFOefFWItR
SU1BM62LyHVm6oyYY6anwMY2OTOQxcP+uuW3Xe5hi6XjZibha9sTBMa76Wvm2I/2lgdncCTb9K2U
UenKZzgCQ80RWYibJw09T5DM12crLcJv1lb+KIbREkQgJh/SNru6wDa8RS0GJD4a29PemYA0s67s
h2qHu+qHn8oCrOPHZXpmZLmj8TmoqpFyY+Zuu1zXLd8I73xZm/mG47y03ozzE6sycwuwO2Ilau4A
Iza26Hu5Hyq0ISgsRx+fcUn5JRoQAiEPMWQRe4mvFCzpnyQj1yRW95KKUxBN8S+XuSZp+AonjT4Q
pqSGKBzlyPLi4OAPIDjI2JNKvRZO+7tKjdHvc+nHQVxNSHLwxuwb6iWOBA3bBOe2yKvhXPZdA3KV
hI/lk8YEd8gqvtPCqlkCkauqZIZPVjnil+DyR4qsKhfaBkAsg32AQRnizQHlBCjQ+qhhxB2LDTTd
f1Zg4mgSOQbWuuuZp87zRp8EIY9tPbEckub55E5jRE4BGjDmEEn6+TTh48ba2LlVdouhtA9q5E17
rIzgs07SZho7hzu/Cerd1fT5DPoPUK0Q8N0B7PBJ9oKnHoBqtlSkq9XTHkFWZlRWJAFWEtbPwgW4
z8ODAG2oYXhbG1V0ohjC2c/muCbBk9YfbZznLyup+cITOr3RsZ2H6EkWe6YSkV9b5+wRP2bO0z5l
mTsXZ6ZINvY75iYOfUFM37R3B1g+gGkGryDkbEszNeZipYikVLLcor7ZjFa8RIY7jhYa9aM0s6Pl
TaXtZ9NofVwfxgvZz9oQ4R08u9p+XaohmHKmsLNpc5+WXvsF3Qghsr6Iff1R9OjFNdRLJ9QTmzEG
1biDimC/zgCTVsaMuf5OYCH4KnHZk1OVkkIzUk6VcTZsGyt7DAlExsROQzH4BSgaawH5oDgopuyG
ui3eDxRbe2zNwSgktisyIoMngnR4ZpKHefPvWfU2WDbjQB52XYlgCzeXI4yCIIntK+8wIIUnBK2T
DbXRjlCfqpkSyp5s0B1c8dh9wzQV5dJjrCD1+IVvxC4avmcquOFBxgjAyuDrMhQgRsMd2xZzj5/r
TbKK/4n7APSsMU+OYKxOfE63MWua0WcviGnNokDqPSd53WxazioRLpP7jZeAR250buaGSwK4BzG/
55J5bdk8KEIb1ZJXvxxorlny23nZlvGWSSVCsrsKYydMQuiZ5IipCx5J8FDiF60An61kog9612nE
oO3t9IWEv5ssEoRM1YS9fYuOBxLRHOwYCIrPLbxa2a9yr+GoyLvbIHBZ05di46XvcACooiPzduhH
jWQ2Ee1CafGSNy1FON2ivcKm3r38y0Gs3iYSvr+KPTYbKX7J3SPA91WUpTz1coZfUgT3XFVu8nsL
rIBHMdmq9GOeycetsMXS2G1lGGvK5s1FowCGcLX9bgredjnyAJgYTIIYePQ64rAIk3pDQ56Oxptt
MH6daa8c2Ray4sVBQPe3WXGCBiArVCx7K9O5wJzo+DiHyxO1INWi1XoPJM7rhrBNvoH79kD9X3/i
aulARzo2Hvg+pbh+P/d1LVCGw1oI0TeFFSL5GjRTpiqnpVzVth5h5GAs09KzMPttcjodjuIvr0r3
/IFDjjQu+21To41rEJdW3leMKaHg2lc6mv+BdJFlYXuRj6LC7agMFjHpDxpAa7wM4D4T8bjNa+wK
TxHIxVcrkYkqeyBpxcLPnTONG/OoPF32GfXHUTG1otnxi7eNBm0ZXOA165TFxg4FnwwyvOo7llms
l+kcpoqWZLjhDuIOOsLzEthNhy+8dsk0F4ushE2i0ACWvWPLAVBC0BhO0X2lgXzdeYlJyMC+kcT9
34BD1sYhRG/GGvx/Ma7TfzFkvsdxvl392l167I0yG24lGlDZcUvp+xF1gB+v87xudVfzJUXfWBEL
HWLoe+CBAzEIKzLeMhayxmphTDWoIC+mi70M9I21KRgmruW/eFMK1Xdei1/YNAhN+zX6kzC3j0Ts
lqloOgqS3dhMf5mMXCGTto66l8KWnlni6NIBe1ZLxoml46YqaEohxK8bYZ1HEF2XatbJLi+DUbNE
Ls9vYOdvO310gUtVxtwF3T4IuujCm1GRHK5KZxBJVQFa8yjEQELUzuaJdgkdr/INJgZf1UXm3pvZ
9G7D6X5O0djhCbaey23yCvj/coj/YEOmICUMUBzML58nnvOQF1u7gjpESzA0VfvnNkWAIRmwIxrC
GfrJdjy3lMkrDEYzzl0a8DgpnX3gcuYGPvgZC226fDtmYQnpYAV1TadKpkC80z77gZFITeeTsnjS
QHYcQIDDcYbx/ZlvrQ/chSOrIBxpmBAVPQFRWRuNhRuk4FBVncC/3i+IFrZCCxhWF0OCXrZnhUC3
P60QbdD9LORrIb7YaaFLDkNX4y0s6Nh8rtoy/4Hx3EoFUGA7/O0SBv2rNYN6NFjl0NdW9Iv+w1h8
qk6rrSYBo1ak+I+69w+cXbPJaFf7OdSy0LFyuZn9EqtdD2lasVu8jR9gudCiXEnCJmVCMlD4rzV7
AVal+Qzb4IEqGi2uRVVhRqDXhexapaE5Om6xicQjec27mV74gQGxPY9LA8qRgHDUIYnfBucOTWef
/smNhFhLiMAOYEbXyAS+wjRwntP6crlNS8qT0Wk0sHvwgVtid3s0teUiULR9HiXNyfD7fYBYS5GE
1ceYRghoclHKQQCwrOsKiN29KrDCI7u58xkUZSsaeLuU0cselbhY7ZijpRYnOLe+zgvEq4ORFKA+
8zmbV3M9Dzi69xipcqB/ufyMCIe5EomZgTxQFYNZKczIxPvi3dIuppMUEPGJr8SQskREnsqROIL/
BQL9MIU8Ne4T4v0Ny6Gkn/Qf4sCmiEKws8RI36OG9Ocu8zFRBdeHV0NRUsXZMKPSpKkiTu4lFWJy
iAjtEIublNysxB5kDYagHPcKK1VWxIblkj2QJfEuQVji0isBHTs0+VNkqkPQA80dJ1X3MfryBF0q
By2b3SatfypfE2sOQm8aJfA05w/AcTR9YLx9FXXUF4uo41v5D0yxaQXyLMoLEdsxp5qdiGlRkTls
KLMCZ+vzK9Kvo28w0t/3Rce77kJI4OGAfOe8BXwi6Q2AU4xzhhMHNVYn1c+4ci0OikY66hvSvOpE
/RlzHHg8lkJXlIVYl5koQwkiGKDhGDoBzN2ICjXV/qOy3LGit7NCFG6FSC8I4A7S25i9RrU1xM4Q
zokQ2Lgdmt+jtZoRPrF1ZA+wsVjeQyomgjODwwRLzS/IG1DVxl+UFz8pjv8W7ZCEbcNC7bddggyz
v7Bhh//OKcV2c7nEEiuKDsGCKZe/k1h1UuU6RiN0QCQIGrBfSOBhhBwAE5VGag5Rkw4Ko6McB0EN
awmIEWlgtdDvVJXwg79yXRXd4/QfSb7ouhiRTuydp1W/ssNuxkIhyk1g9+A1i7iKCrFvYeTLyVsb
YEmRxPxFQ7QW8ehxGIhhwV8NDcEmD6Y/B9mbe65obNKrfYDp3sPcXIBYE9AHB06Onasrg5ExbmoR
bJY1e7EqMR6OeB+Pny1Gnb/Fzhs9gRNoa5FwNk2I/BVpSXRtPeo047LBAmFtFCniCvYcsPkzVoMr
Djyaw48TbIsyoQa/XJ5+scD0U3smSY0ht3iKSTWSSFMHQLP9LUK1F9gnutwcxSDBbud7jU2YWrwC
/92/xXgsUaAk6BV5ouG7wONM6mpbyOSoFnA3tVvHVN5LF+IJ1/qu4KVTH1h2K5ccDoKl8R3lCuZt
lbQ1AKs4GyqChtwmfY2h9aPGssBPtU69EyeoB+EH/vFuX55sw1pJFGTJ1BXZipEFFE1NAsTI/Ue3
6ggGlyUOCQtLeNxD7cej6M8noXipgaKXrNK41X3VwRxuAdRj34MRBd0DW+ls6NzNCTrQrNQHoZc2
IewczQ5ThrUSHFSg+dV2dAiGGEgGGEQA+nYG/i4UK3Mt8rI6yv0BJtsgeswluGe76yow73H5qCRL
aLHsCQywT0q4Uxh2/OPvkJnFQHaVk7nZdxk5xn3sigASvfDQtAI7tQwTlyK/iMcuFhFVg8iKIA+f
85U3vlI/C6gIeM/9dtH3kvEDexgMQ2j8pS6ncKjx83rKULi84k/6fdju6ENVU/RShYtTjCmqGUlZ
VjZJAEAEWfSUK/WSkd/evP32Lf5TxqAPAFqh59aWR+g5NJPKRDuG+1PxGt4WHqaMgzDTYOkc0f/l
j6eYYBJc1MRU7RWBsNs+LV2QxbBAi4im5jDre671ziBvU4GrycAZwm7JbwhXJYcucQlPG5Hmm2Pq
df9MUn0KUNs69WBHplJEK+rXtzK1Frbo0UrwVyeLJGlxSxfbmXOVlW4D/ma+wRaXKzeqNLd7rZAu
vWiCgCMID5ibhbyufW2/xpz/+P0tQ5RTK5HZh3a75I3ut5rX0WHthjAKXBT1cIaRwIr9asHr8omJ
bBZQDiHVi5RFRuHZ/dYa1Zg8xvBMrLZc+6PXv6B8cb1/dr9sUQ4Tc6NZPObfN9Fd9mP93Iut0Kg7
gqz33yrKB5o/YXZvZbaVhrMFVSNfGEkL07wV3nOLAa6yddFE6hofdkywZHb13LCrv+4Th0+zdFnh
b0368+UcKnJZmG1dRg2bWZ4qLE3eQtf/VfaL21KUD4a9YAdju2eGDQQDTPw1WBZ5rV5AvhzD4M4X
Y1QIEuZhfe10cD0FJpusXawZgXSB0GFxwZAX/YqOrVU0onFefKkce3QnF9bir65WByto3DbgDDvt
EqaK1JKfAt0kLyzDc8+hC5MXeOaiAgH/TrbJrxsh6+Wy7oFlcIVAdVNsLSEwsi8881qAda3b9Fx/
VyE7mcq7fqIvTyFLrx/cerTU5go3N39a1k9ktGw5g/a0/USl+e8TxGsI3cOgjeNF/HxXq490IoTY
Z4Du/xPzgEFUDsp6aaqAVLPogcT+JtepEdmYV8T7KTpjigr6oi99Aum1egRsPHzvM4gJPkM3O4yn
h4M7p4yTqAhc4Hm9HXCzMxUSjxobcuHVMtk0qT2vtvRI8sm5NoIFApjfyUQc0c06Nk7RmYZgnzlx
1CSZsxqwIwvV1Vs9XjKNARc9z4UrtS3bu19tsS/MXEwAm+PzPf1fPSvWPrgUbWE9fJD80skKKtOS
9lrgGnMVVVw/r/keKCYxrsqTh3e6FBSXkjjRcwDByhLhAsjbZUKb7F+ZuHNLBsCcyHR9P2oBkOEl
bj88gjQvvYiDDdkqEcGvmhVR63A3iCD5Fx7dXerMXTIq7jzEzwgOnHet6qEiuaWHPjbP8SwhxaYp
CZWtkFd8yvzeCCvM3jinCRQ0JFk6vTcVBwNmbD1nxfA3e+Nq7sT16fArfcIH1NJiMUZZC0qBqgMT
JdDSOXYhrnsGEBcqeLZAhM62ArXDe3jFAJrYA3rNgdD2Qe1wnvFgziZiG0Njo6oqVfeG1bnX0NVq
gjg2XezEF76EoDvrB2JOTZ2BhMBFfEE6u2C5P//oLoZIShY8y5C1SiL7C4pv3+WL/s5sf/k3nnwq
MVGRsog9Uj8nfzzEN4BiJCnzQu6Bfr4Ws8Lv9cuthPXeqxxhISvtqls92LocKnM76zZTPkip/TlJ
feAaj6MJnEkMqGUMo+MqWKCLIcV+LaRCiBKD8nPc6+cOlKPNTH4syx8/fa+wu5wTtfHIlcp+8oVm
DpoxSoHOXcXGXdT3PRxCke2Fgr7YOwfPjx1N6JjTqpUG4uUJnvqcXFKpJCFeKm1vYMpV+q8wwrje
OyozYp7n8Me4fIIPBA1CFiXeCWoteUYcjmEFIBEKigmKAAjNZzsaVkmsh19smBIMtsA8JtcW5oaZ
TrrlKqjTUvrPQa5xoU26+B+wm4xUSPQyz80scYzvePepa0IMmPmLRWUmmiVSvYbfpcRrLkEqIbBO
F9LYCM50sb0CIquP885zixWvmahxqHFm9X5Bj2WmulL4BOD6tVU7f/lwpL18qFNPwyl3yxasBsPH
4neAVpAJrniN+siXtE2LYLDxpqE4uHI19lTsB/6B37Hb//H4i7zHh8v2WsALfxTkAEjdvKc9bNov
bJDby0+xNW/VWdKTd7S5BoD5l+hJRyaiMMtJs8NEgMp+D2K4L34lUO6Pyb+J340K/Dfn1mgk+PJX
sT6yWm+JbtO7w83B0uxZxSFMMHo4EXIWN0IRs1adbmabkNkKw8qEvPvDDmViQuJisGBpyfIk0s9S
XcBjULiZxWAhjRq+mCo89pU3BrJuwPik//JzfPvTi1umUXxpdn4QN9q7StccK4ywAhpfHdoNhrNg
RHPCVy0MUmJdRJmjQKZ84S9P0JyJ5Fc5v7L4xwzMUonKmqji0v5STdNu6ZAQohafrGKi5i84F86v
n2A7V6vBZursYj8hGxRPyDQqs+UfZyLiEifmwCFx8SIxLLCBcfQZoU7VdJ3LKVRTUWh4Ae7Yh724
08lj7ejxht1szNTPYXtYN04WV4R//8lM+suwcAxo5vxFXirdcgHnCMInp4P1nmsPWl/2EIyqyKn1
9WIGPsWkNjhsg3OJ0R1SibgPweQY1PmEfb5yhpZAXbzPnCdOLJ+xVj7HjWpwr0hQhqlpzqnH2KFR
thR2ysUQjEqRxJYYxNqfCyJu+wIqswKae4AFNXAbAjym2Jinx6yPoVBxWNpBfbHaoRc3smvyr3x5
kOm+V20pWyoUC0rQUYpdjxhq7ikVxFRoi/XrhHYq+jjzZ/ogDxRPsw7lK4TtHNeNcSzD/SkqwuCV
NwIsZ/ko9O/RyxQ5sgXzvdr7wKzdw9IIZ69cgNYywbQRYHKcnotnhQuiYkbLic0pBN/jYXXiLiJM
5YEAsubPvEkA4CqUTA/s9qMKcHj5FK/BGIDe8I+0slUpZDewbb1WOV0RkIbMV2VI6IhWLfoq4/Vx
YShACxJRrx3d1gQwntfdhRWxfF+Mli0tlDsOt3dXetZWWm4atjjgPY/0JA/8XxvRxKov00cThuxd
LJZPJbrkJeQ8jNwV17f7RjH479iF1UXPjWBynXv7GXIK2MGe/trArhC65COEtw9s5V47NVPssAyd
MYbk2csmf4Q8xId2iwYdA7zJULAUXOgDMUx7S+0LHmLWA4jIC7PpXLilCs1gpGgCavqSK16SaatL
bUxRQMdFlwvD+rD4NCuqqCo0Yb5mBjBhFWuDxPh3ywQITXhiT7x1RBEHvbqJ4hu3wQJx09i16XGz
1MGKoixtyqwXqKA3jgjxmm7NdbHvJlAO1shoFOuXoBjLHDdusLaMx8iWe4zptyICt8Q72D9E1zof
pQEmyHTv8FZjpW5z6nej6Hxn7QhkiV2k1Ehz8BfU+J4iMreBI/sEw/5O+aDYI/HK3W4cLfPHpybk
HhgLbFwtCyQzRDzM+h76J0w7OP9fT6jEe1PPdteaJV+zFk7kyu24E+r/fNmfF4gomH4F8jXtb9w6
ZVvTFYTcKAAt6rQxNKJ17RbUOCo/4DzR1El5D+Joo7YxakWR1t3dSCHtSFEH7aSmYcS15CviCJ0e
rsjsRAoJOzVbJO0kzhfkUiMJ/nMiqOteTxLL6adk8iXo+weNFuJvRLeOtLprcSIg9zkJyTFIeWrx
eMb33ZtmeS77eywiAsivLqI3BizAzNAxpZSpCyL/oq39FyRh6umRrWQmlFY77t+DMlhv7ttZuGNf
K5u4a0FuRpYKL4WgI3Eh43zwjy+5IVcamkM8odQFOq3SeDp+v47P+XzRI7SNIqCYcvPu7NbabWsW
OyScdziW8oL84pJ7NkkGsyKK5RuGrY3MXuBqF3fxidj8+immpRrvBcDNIC6FEWJ9yr7i5dtS4kHb
LRtKs8vDr6oChaO1u4541wJNvhd0VncTk6AucCisMgxXxbXdinMLIf+K1vP8m5pSiVu7RWSR9H7l
uPwuLZfNrOcsRTkMXTilZU0o6f913nEejbYooXPg6Lv4mYvDfjBhaw2AtIRYOJyx3rm8lfUc0+4E
2qee5Niiai5EfUyYOHuo3+Ftj0FGB058g5uqt3UenrW+9LjggvS5CpA813sOo2sR8v9ikOn+xsTu
3Cd9GvcJF4Fe96o0m8f17Lk3XwettmjKBqRy3LrFxkMIAr44SCnuZX7vUMy3X3pLwVMKYqHgDRZp
Btp8iQpKG6RCkDFzcpUodC1uFhbG413DlPAxj5Dp4cB3r6ULdpzPq7BfeVxrmJJsgQ70ULUkjdVV
plQR+oJ50ORiXqcyOEB2D0n85Hf1ClEvB8Q8HMlSxpy57lKP3Xk1NrmMOkYKILFWWn0r2plberr6
KLtwZLGeMfjX9S+iitT8+3uiSS1C4V55aSpjFF3Bvt/pSuzidlQSX67MbWCP2qhY/wGfO/kK2gmf
5WB5byCDvo3JM1bvrqldFHkKDQO3wkjx5ECctK6mqKpmYNkWK3eCNXzjqH2B5wHOcYffnr3hq1IU
EfmepeKSC+/D9H1yfAT+rVw7lNsz/76vb7mWtp8fF7wmSwlLXBClS22prgAwKQdReQhFDGpqUW+u
OXNn+uij2tni8Tz4VJQvtDH7fDTklTWauppXrd8pp+1RZ+j7wNSdvon0qgjFm1AzJinjnHOiL2QM
Q9SRYhyOj26SUHrE+Nxw1f1/dtF0sVygWHH5KEDqorseGoH7Bdc72Dhd0UnLFJzZRrC5uRGz2cF3
qu55XjQSCuT7P0+ID/VdlZ+eTVt+L7PQwff9Kw11PXUSIWKULVSFy0b5S/A6Z0pg9761JnV9+Edx
VIA4vVBjeNmamkTWFBFH8o+Cq6vm5Ur0WWczZdZ3/xy+cAwnyJ7WzsegSWo0sNS9scNZ1K+LWjps
WvwiJcakc3bEZnJgTBi14R9l29/LV8jrXqL6jWmozwGgUAYkREgrHoVawXemR2w7IhehPtnifxgC
yOAPKl+4mtizFb0G1PzS+wxI9NPwH3pA8mWK0AvUS1iO6k7+3a/rYpwW8f+3Ynsbp5eJLOpZsGwh
G+BAQA18CMZ7iGxI/woWVdmOcxJGceEYku83K+NNCJMaQJW5GhDc8v1+EQU+6yC9Wv3RkA1MgYYA
GyOc1e5s5CjpDXPX9bcNT4Ry8NijUy0cZFwA7ksi8DBTGYdxhTSo3lqLHrZnVteVZeLB/t2BdwGg
LmVLfrZVxrSNUUWPABlSs3AkrZUz5Nvh+FI05UKP5eRmCNMXjEO/kl7BhWMk3jyoxOGxgHKlxCIn
Rt8BH0Zpw9G65Ts9wHUdLwwDlMWhXXng3TZ5FFjdD7jZYhbnUYXwI+ldr4z2Q3QYDM5GnP1vOWnS
xTKJhKWP9ThjulC16WAJJTQig6SSnkNV8MMWiRv6nCzXi0Q87EOdo2tW/T9r9OpEF9aVPEu27/PS
aeoxCwMURyXkDoIe3lPe4GavsvLkIdJlBrkWie6VXIzKMXgSVR6olPQZG67LYQGUB36WR1leM5h1
9UM9JOG/VpuHqoWfvZR2VANG+dA0/LWLdgwYEiwmVq35HBoYVilgHN1jM4qfbIe7M4J5Jbe3vga4
LeNZM+C7c9oF4BHdMglcvFyLmJimRO/tFgAtO9J9jEegvIuEqEJzp1PyobYHqVxCxF8J+9odIjcj
cAb2Iq/Ns31CFpoAoa1/CbIWo+3U8KcWjvFsIwr1rsAJHd8FaW5sO1Hl/51vWW82MeDxEH8jv8J6
QG6L192sJa+Jwa9ZRorm+/YKKwSgVrTbixnbsvTQAIaJzq03xVmaIrbEvsRlJq+LOF7ATyLt4fNu
2mnKBVhfLBNtyqXQBvSp3Nu01i/MVtfBftEoJ4olJNAa+G29PTl6flHntDl7DUIYNu8wV0qyfwG0
1UvmfR9T8bLGiM1+3LN6ZYNd4uh+B6E/0L8t+HzL0QWR979nD9pbBGrIdVCiXq08hbw/Aiu8P4b0
+Qic1cj2z8WW0Pgpe4w0iAIbbnj5PSa/CzNdpYmbH0Qh1bXxZQDgOsA5qt/0FxYMpB7hLFPxXm8u
YdXv6bEvqWFhOzIGXr0W+kOOlOBV5EM0L5a2c+P7X028tpsDr9lPUtG35Vg8EwziwhAu3k512w0z
tUCMFFCpoZ1QM/bYnVRHMXN1l1SHMV/pV/D8A2jMs8G8GZ9PmieDIcGoMDYH9TgAz//H1E6LNLZc
QcdozwoloVQrIuKgYopTmTy60BaZofHCroEa3gwYC552H1Nk8JQnM/5Re9Y/cgSMBCiacL4WN+gq
tEZSUwDfMuYP68EDYCzOR8nhclcRqO5i5mrvmsx0W127xff31LlJmc30gXK7aKZt3AexIJnVpkKt
DxilodHl4TjgV+r7Npsjf210a58Qsplz6cSifoxuVLkw7RjgQG/bVuLX03ci/e3+aI9AETpPuQb6
GVxmAs/2hAd3bsEWEWhA/YhLRq9fNUQOAwPr7efM9MOa1323M2CSN3/WW5uxY7A2UouMlb4PaHWX
P3qRZq6boLrBN5inz9vC0xxPyd9wVYEKUD9l5B5jfvzI5/JKhdEvHlfoLFqJrvKKqMtWKRDOY2yX
zYfXZRdoEfpmXpd6sdBklo5oeSNReyeP1qOWxuqvRW364ARo9qoNvbcdfyU6R685Ba9JVsU40I3D
ZsStzrHgZDrvX/tkStGQBOBdwa9rcz+2oDlWYR8x/ePO9nY2jJs3X53d9FIgYPKfKTcEuHYmmXcf
K1msS0O5ejRo0mtJlwXncYfFlnee3ys6bxmh3dgZkY5YKpovk4qnlVo9ZUmHvcZIMaHA0W1JP3rG
DvXK8yWLYnqz9pqP7gY8JMdKIDY3nAjWTz0u6/jD42we/zaivy1+AwVZ92SIDQDdaVLjjjXo7H6G
pTMz3WPwFWrdUAaW0E35b4ywgKN90+HaEZfRb/hheXHYfF5FiG8gZe+29bkTUtpIY9+dVZ3NuAcH
4F/JbS5vJ5J37mssl98KdBKMjpSfsdnTuRTsE2eT4gRYWqv7yExYGKNVBmOtI+m1Bd4rE5cK95ev
Hpl6n3JiMZo3kc58rE4013rucHXBwmMSnt+3GmiEAs50dRtSiQWOL9OF3zuruwVxIJsOkTRSAQoF
4airg4WutocUFKodFDZYoStLI3Cs2kfiatfM0ZOfMLVQCRDpqMwZxGInr6fP84d2lUprPXRE947q
BKyiIZIaFOWxbsCbxES71nfuy+YVuKCPTUZSr52fjY8M1dpZ+3TaXDrq40f+jfijl8KOOQ4nD0FB
Y61ypGz2fm8hJ6vWgcbGyHdWb/ugyLK6J32+BnMReDjkL1BYkvFRPVMdJqUkru+p529ZNRWhB6Z2
krYsvatmK3ApRpiKhA+ctOBiOzUzktvPoSmHpycQa8YRTfByHm6oxgNSukQmCZeTAs/DmbQwwL3I
DlPmnF/yei4nwTGX0dlKZ6zsvC9Odvsnl+ZhIEbdu3ZpQ7+Bx7Heikhn8ADiRcjpgJgEbr1yY1iL
meIZ5CfPHuKJSxe0w71t9otY6l1iWd6K/BD/jlrZal98ZJyRLzuBjxZlPX7Y11hEeirY2JU8xDPi
ZX+705ShUvtw9UL2j6yB42Lbf6DEmuGxpgLxipUvu2ydPKc9+w96L1c6WoEL6ksaCZQj0U5FVi9D
xi5ZSA5H2aPpAexHwGLZZec0HDQ2cnCuigX2n03dVEn4iMpuMYoBmChVsCUIanSU0bQM6nHbBZv0
MUblEJVp4s0UEwsI7f5mhD4k+Ekva/od51EKO2KOLx9jRm51qkgtgBlksNP36lAMk6G/3axN6/eX
ZvP9jnzbUTPPidagX83DU2RnbzBUuNjbJnpzag86Z7HD2gO9Yu6JS4AmWlbejJUngik2sXKS4E5w
iJ5QVvIvaJeiJ09+NrbIK5Hp2gd3QtSdrOCHkK0Slnt3U+T7sdraM38IhoVMLR0weamxX1m40mzH
D6xivgqG0OHJ0ObW3swTAgxzCS+mnRBw34aDV3wyoIUFPBqUCHmYgrRttjodxq7mRFGMjZ6Plcc/
U8GyXlnTYDHPM6gITmiQuraBn/hExsGYA3wx4NEXXjBbY5+162Fg2qG2XPsOJiqnJA0wyn8eXhKh
P7hRmI1Dxdmzoef77yjQ4BhUIPVFY3O7T9HdNCPlE4rr5zoGrqxHU95tsPdUdnDZmYFvsBS1LxIK
swC5w5r3zkk8//kIifF/AfB9TRmcTaiLZrhVvo6yywCyxduO6kfQb5WKKtdkjDB0cwWy4hx8lCZC
rQ8sSP0AAnsmSZc+/62mnZMpdrFeYnRapWZKRiFvVIaSQXP7hnDuuyVJMt/O9p/cw/UgE1AhooKx
0bgcsAFbpW4uFRVk2Ng959A/5BwnP6J0ysaD/cEastL5njMWI1zwcLJ2QJVmTsjpZY+ztSxOqoZ2
UYSOnWVt3QEJVDMKxxACJuvJM8sVg/bxi0MlntyZm39utECJA2O2SSvNqjPkPh5i0U92krb3VsY5
B+JfFTRYhD9WVJv0dvSuAuGesm+ShPG8YLsr9XscKFjfBDULfDtiktyE1r1Crn7fHA857XVPNY3i
RjeWfBKmKr/Uc2p395vgNpRIUQ6mfG2jHXBpYUK3jvabgaq5KhzXUfXxh7zUptvld5MCmotEN20v
a1IEJxhia+E4zKixq7zWn/SN3Uuts0TejHLuVNRgtWM89NS+mIdgPc3lW7FcGX+VGrBQTnqMljI6
5FV5DShjWNn37J4k+9g7Mfdvtlc0LTmAfnoMhaKZxvTsLMZjhUpddS5SruXPphV2mQJwAt7ESAf2
vuyigNU9DdpnLq3HDUbZlph17IBDhDcjmx0r6XToyGnoNUOdY3CyMacaLtZwd2OHrbrjs4M26jsq
hydrf7PIFLHsqq1XDajRmvkmcjaXHXEfPc9qDB9vGFWhdn02v9O37Uoa6WZwy/RJCzssCzC4iK9U
33w8y7gN2geMHz7YxAkepdpcPtkqJNn/N36i7paKG0EA8x8/aKMUQ8oFhKUxh+3DUglMsJB14vrX
LMcrAUO89RFjscO2uOgrTqKCseKiz8chJQAxkElRfOmAaPVhKiFIspkeJ442LWcAB5Qdhdd8P2Wc
3C3qTJMBYDo4wCG8kj63onkVoDIfYhoSDNvMptenNNTXJGo8zVNuH2O8INIryCg6Li+uZireRaPz
EM1V6JQ9ZFL0s9JOkDTwviGdu9u42CteGgNgj0SnSJHkOVDl25YwoU22CdelVI9UcIs/FOOaHdEr
EbbvRkE7ZjXvX9kZdu0qC3plOhqGxJvaD7KSVBadJsGCzXQkmHnbSuEk3sUwUASUhrCK1nkYsEnv
LICDm1ldesrVmsmYjTE04bmHfCuPS65JNrm7MuhEoeVYvROcVojb/ybB0jzTv06QiMuo2TrFxyk9
AJoc+ZhJ1A4hF2hffWpa0OjPPHeaJCKK5kYi+Gvrd4zBU4HsGPjeUenOunfK4TU+eXk1Li9jNdhh
4S3XJCkcD11K1CpzW/viyNG5HrG+0YgvJYXY/fQZUlCD2tj0qfOq1/OL0N0s1jHT0fqK6/DomRDK
Tk7GB2KdEJJGQEIeNxtzXWwrdrHSj69XIrgnQ5jZTk0dMmQr1dvTFFj29kjQO9UTDqBT+/jwf6ET
d0XUkAVTv5WEwk+nzVaPX3dAKpZwaisy2YOWblYJkaTj+9xQyfts0Kx7HYzsRE5aLpNbx+/tkVPA
5TS4yTDZbv261SKZe40Wvr/DynTTw6ipWCsjFfDZSAvbdKTXMGHQ6uZd24VD31+1qxGntcc5FhoJ
v7Kq/RFgxWxPsELsJlXUyHo3cM+O+Mwi111rYA+jVgj10xdkOTQbDu9bEeKJdCdk6FVb73bFNshL
uhZLc6f1pzoUYU4VMNAOaTLJw6KYnMNg/IsqWfNVvEJiILATtBir8wrU3zwro7F4Cn73r3esyZoC
R1Lt+lV5cGNxL9mdxS4kM7gwRjtjsGoLKJgVILUzjI+huWwm/kOEPq+xrZW2xG8cYpmMb3YsghG0
LpTaYMbsDoV/hK7QlOfddqu182wxTNmDd/TDtlqS9rGW7Q2Nnele0QciFmkA4A7G9iVf6S2ImtbN
eGPH0ge/mvNdmQXaU6k60XrZsgFWyVFXoVST+diUQXjrZBYWcaQe2kZR1W9MjJYAQ/1DmgRv/Tcl
JTP7lAM106r+6NOyTeH40bqslb4LCNKO3TmvR8uc+jgU4waHE6fEJYIHxe07pGPGZpLEUJMMj8Qi
IBapXg+qRmobxlUVkQcQZeLn/sQpPtd57zzSdg4gZ4Ij8bJiAgV3WR8cqFPy93yQdPaYBWBVvdr2
Vs2JOW6QChy6gV2WiYI6QyCreaeoVr63QQdr7+D8GB1vS2a26tOUFQUxXzSISkNkiszg/O2PXfli
fMXlGvlS8PRPKvdFOdUipFcUHC19N3TkKcvzHcYlWqvBLMLgDRbix1RKfeOZ5cH+Jc1d57Y9pE/6
uvk+1RLmnrrHuLFkGEQwEXr/Ej3FoUpyL67YkQtBxNoLL+3AAB/7OAZoSVBobf0UgcYSMybS6FOe
NAR9LeWGHL+LvT/FfKskOqXpHHLj+g3AdvmOGAP8tbRhYmpEUB9jsdI6rGBQmmhSLr29kFZSw9h6
alxQniSHm9LiBQ7lQLZXYKySdGZS+gqcPoTH+FRxcPElU8JmJ/Mrcll3N+cBKCbF13z/AZOfpClX
RQpcKusaIuy8dEGQCe33bOa5diKxg1nnfCRoGzrtkN128ItoRZzyMhQHJ8NB1jet+uxCFKVAhh0B
IYyJ+qV9c6gzgCdxpOYsHhwe9ErEV3p9pdsEnEphdp0ElcleVBT3aei8mf/Yl+BqRzKBjtHOXH0a
I6sZ2HQFUx1CduA6NUOHwfRFkgvvzPrl7A7/4Bn+W9qnFF9/G7S702rZ2oRGsSW11bjX7b8oyPuq
iQsnCXbnnJ5F2wsVeA50demYboeE0Vdx4ZBH6jAxrGct6FBegfLclWdCa2TsmNSBoBBGr1B/Stwm
8FSrE/CuoYC3lUrNo035NoqMhquUMm0rmx2KD1xjCDPx8mboTR0NgHWBoHHPeOPCXkpOi3SCmWF+
F4e7by3Nc7VwmIKuniq51K48Mo0rJUfGLAnwyRjwxrFZK8dDtcP2TOPDZoeVM4Ly6qVguP4wEDdz
I6Drz2dnu6Ez8rik4uoCMCBB/GhXydE7jcZ3ERxCCRBW/YHtB+scgqQwuqtlXUsXn0nsVCh2erd4
d1+GXYCClOAmfgpwCmD9DzSqdv+YtM5jtVOhpLanDrCkdI65EW+9+fqtLD8AKR9wUR1a81dKrSUN
EHLWplXdJq+4gVZHxy3HrXPAXjRErg6F3PBTLTyZ3dDgFcjPgVSMj6MXdVR2KRSzExR7yLOOAONP
AoJ6LD1cmrahF9gyXV+9XHEKGAQyTAyd5nhp1GVHF12XNR987IWpYh5yVEnTYnl/0pF2a8bqeUr1
mdT9Zi3V5TT6ng8HV6+00ay3Yb9esMuHUkoGjXnBsxJct2RYn8Lvmfu8h7BhPN9WxTqxlmKOKY38
t0JqTeUICNcPyYjmfVOgrRrIcaCauFwe4SPLA/mOAeovMBWFCbj2HjTcUxC78s8U2KLb7rIiGEbe
rtqKJBFrSRiYdR7/je2zSsEyiaN6Mx9kOTQHe2wmRtxrblITgKO8eOKPZO6zFKH8M2aQsXqwHO62
hcbOTg//OtjRt63n7/zF/hRY9AgUZ07xy0kxwAyNoTHEP432oK1cSfeGO4Lb2806AMq8VAKrTMCJ
KmSsYtWoejJKnhFsUn524XjCtbkGBeceJbCJajdbHOeVoqXP2TdYo2ykYqwYDDVkdgVm/Ez+Cg02
Qo+EBz3AWpoiSTo9Gm9j8fu/Ac8mn9K5L2jqWDRLF7WMTkEHqt7r83wo3sBaexGOLYzv/BEfwV6T
dUg+Dvv6z7zzNNZho7M3luST9QDR0kyyPIEsGa81SE8mGQlPljZcsK+mFQvBdC0XqDJtWHgLQ+UA
+ACB3UKRbq9fklrEahWyM03s13yyigfzibkxuW7c6MAm9HdMQMzXMQZovMixE1Q/3bpEc4kYuQ5x
DyM7YOz1qXu7ydHEHu7XLK93cPs8B+RsB1FSoGRwhYEQA4dgfn2qSXzDwq7MEQhcwjVpJQI0Vw/4
pZEcMuuZhL0azMtrCAP7ZfhPBie49MV3VE5eZqzcTADTOvipD2FcPQimar5Hex6JB+no0NUbs34s
FP/dsq24p+7raKqiQgPe7nhhJYpmfq0+bSQV7vdhkX1rExgIeAbAMnSrkyYmZWYfoGb29lzBHof+
IXMCR2gkJaoylWEqh+p54LKVKw2JgX0VMcovx6PM15+oPJ2l4dJd4VZCW4BBPUN1MLWAlD1NGthB
HcLkb5yjkYQQkEU2RaRDcVqWX1XdIh5H/YsQqrFUdQQyML5evt0KWUuE88AXkTDDBhUltsO1N/vL
eq+JLLxnFNqDfy/zMISHHiDfJoFh6A4k/waSI/TGgBEvGMNtTbPCxk1FRhlWMIwmPdsB2MRDFULN
WVgZij8dzUo5kqq0Xv3c4vYZnubf9fg46CspkbtvY792HOGq9E/Se5/SzLvQOKPoYUUgzmVg20RC
UGwPLu5oTJor99HJtAGMJ+oy1kQQgLqHlXdKi1VBHTAkxy9qLdHc0bVPSdWfxtE80LSYTJCUFsYM
3uN2kVuef/KCAHoMbY3buTq9bXFk4vIuhqi8HiVkokd9JGUyARW1IgImXtZliWH/BZ2HmRr1qCMI
FXaGiULnpMrnjKaFY6TB1X7wspjby8Se+SqtPPygrYRW0idT1Uo29TmsAkLBnCIOFbrrJc9Dn78c
GU7zm0ZNXXTTW2fhyVp0L0sNMCb8OGt23ukBNLcFDdiHpR50FcJsiMkb6dYscftLpWl5rwLGCqVL
5p5TB92NH8GMcHaosXdMFHODoCT/GRnJouUoA8l2/iGHDJcAVxEVssx4Aswmn8JdV2EvoDVaiv1m
0HsV6AhDQBemHi3o4qhNeN95M7/CVqTOgHrbDvVe9z6EA2VLGWKKVaISrz0oPAqj/CVF26XNvucW
bOkXNmueg7yfBOnAqIWLa1H7C2/wKFdHUwUIVJOTPnShDobhspsKV50fpJlxh/Q0Fvq1+cOJY+Gk
jo5UndLbRlhqKpCh3LVcTqCk3M9C+p3qs7qO9p81BtkkvNj5f+yQL+nrLoJcKNhZLTydTgSbOaoh
xbhmavxY5DfEftQeCExidaWud5BwpbVU+KniPgmvUPeEXiVuYXNqyKdrIW/lLrbNrIdLcap35GcE
6Dpj0ZnQ+Hu/x9hwiNWaqQYoKtY6Uslrgq3x/VfZiKu0xa0r/2pNLFA3iBbNIkzk5LiAD+NmEHxX
nFIlDZOyeUWOnDJYYIaibPkurhVBLDiymCyUbtGLyT8RAx3HwkWf00tVp/HGi5c2cusy+m5gUcgq
LtW/YpeuD/ugwiIdl5EZMGtHqlS+dKDWQyR9/LNQ92lQRaM925HdIG7zEuJynpHlewvitxHjdWtP
EJ6FWB4o15xPJbBSR/AcFDSMP0rh80QF74RImM0o5QEXjmNKePZtNXQN08w5bbrY1yBAPyR9wV3Y
jp2ogouvYpfkAnksOywIm/Wq07UhgoVuYfMCw1eknojsGQnxcC05OwFv/hAgeaT+YgdDdR13uG/j
D4K6KTLWsvfwTMAJWQr8kNA+1Gug8ujlD3hDSMtLMkDkFfLgV4oin/xRkT9WPx9P4bzV2Vd8bDkT
vyu2M1nnsnN532ct+uxu3zdLU/mPwMkzHnRyA3E0Mu3f1TnxJRlWoNINAKm6QpAV9OJEhj5td3fy
L8aCLsVD2FNTU3D2J8JzoUBPtztlb+s/oyqlTpSdsgPfE0BtBVNnaSmoySHOhG4tJH9QVVgAkS9f
xSyFBEIds+eiNRCaoNdLrjDyxtlDDEKNaJyzY956qiQHYWyqjZ2aSczR/vpAJHyTpq+jbxymApN7
rESXCc+aFfgsfUtqwKd6Qu1ve/JhMuXxTMNBOzs05R/Q4Huf3zompic8DPoq4AfwkGag/aBZO3Y2
bmSddmGJykmh90t5P+iwWfqhuEKgqZUabgDIlxtcZoc0eFI2uYOtVNQ6zsWpDAOI/vF6054Asfas
y9pATVK7LruFdFJsdav6IE9FMnbKXsVLM/EuIXZDqMfUO07sqLe96wTIIT/ih3pelb2C4RBOWnxB
c66EyWCYhqgri7qCd5nRkX5Kmu4LRqP0boKktLR+5J0t13jlMlJ7A6HnQoN51/qiSELUArBFDMBE
/r3QJFRgUE1BZdObxxLiCSyAA1Q6ezxod+eMPBExNXHR9bTdyS7FQbDDjlNjjDkueW5/LkOijsO5
bX6PhQ3bPp9pPtRTYXKPKXyQP3ym4hkjcd2YqxSQr4Zs3MgpN6lGS9Pgf5sXiYqV/gucApGsXVWz
80rpjlG5ZnAbUTSJrzbU2aeKUiXcZUs9bbXC55oM1bVrQXEtliuP5VbQtrLzExSjVMF3MhS6iLAi
Oe6k14wGoMRNQ3O5R4JUeqySInick6B7wrhNlBrQVytWOSp8Cx5biWpLTny+CvYqy83BLqBtYhjL
CfShacrw2x+I+GlQ/xCgK4LFO+3OgXtL4Y0WTrA+DndVmmKylqZF9JrfGBYJ+U898ALdQq3ENrFe
gqiPMwZNfO3DKQMtz7skwI5tF8UznK0zpkLE0qIyAzRkJ0XlNlFXbYT0GXoD5gFLefbFGj6AlsPI
wdyqsMOQiHxB+hbwAbJ+h0M6fFgW4u3J4c2+EDJW8dWTN1YNCDEKmIiCokrYRCWtQ9XL6DgzP1E2
VxE0Wsk46rjUe82kZNPjI9Eq1x+MW8bhpirpf7Pl85bWhGog9Ecyxkb03KUcKFRkDGCIyKbzvdGV
5kaxv3jppLpsiUdAcyzgOMw7i4+1a1ZUcfxt+dIqTg2A+o5EKh+3K2KTUawuJuVmh4GdJz05+HpL
KjuDNGxJRmPvWXP3bUMpdha7mdz/QCrkZLicdIqG5qKUqkPDqGuSVSNHeio1XTztlmHI0xayviYQ
mI0xZ+rpGwv4Y01/HJTY4sa59y258iG/PaXs0Z3zSZ0oXJ5/9VxOLiQ61l7OJwKZXoTdXJzAgSe3
IOuff0o5kBeEXcqr8RLX5/bhf5TJFXR9aCW2fGbI+BHzO4O5ppJwKF9/BXJmM1TxE/xEjhdAAayl
FSsAyGHBzVOkgD+3vaJ+t3ySFD8t4bByEcToyxnv0UsdE9sj/DL8ygazS48lv0ldeaDSxw8TspHp
2efFkqxD1dvwz4KFYbciwG4NJJKr1GkugHJnYbFOnUsfL42EqGf//zxJ/nc3maqYu6ORcOIP8RGk
kouDYzda24Y9y2g9LVMQTH03AIkXJ+ObL4G2/3TSdGTCZCb9c0pYVrNCNlvX4/+cOwodEG/qCdQI
E3WN6M5aRDWUTTI+FKPW4JSeOIso4ku4/yoskBUP/GrUIvz6BhWBUzIMYwZwg+DXWJ3dhTvGFRkZ
3Jclh2pUyklR2Ae3O2+Hvno0Sox12iR9guu2dHRAqEmr0IiQTVY9kDeOkhdfn1IiQUcmWjrOVtv0
q/DE+6AlrTmpoZzakg3FuhAk8uMB5vfEPnO/m515u8aASM9BTYyxhhCsvX1F0CcU/83L4HODs7EM
fHyeWVOMnn8QzEAkPcVUp34s9OCDDgIemUQXh0wmcoO/mrWMSwUFS5UGy/7g8q1+g9c6YM5gK7Z3
XK9N5tSTBuKebezPYVMQ9ueqrcY+Ct6hb9v51Uq7BQeI4OKavo65rXivGAGlweNI3h0zwgo5oogw
EFilZdZcD7SNtMRZl5jfKnvSpS+STwOaT3DWZYGSRx9Lda2jgM1cz8tnHVm8V0PHu0JJeyixy47l
NnMtiu3hLlJo0vbAwFI8spKCIO1FE54/rh3d+9kwHI4xRVE4FdDoRNY4JESx67/TPekF2dnkuVI1
A8/M71F7mX2sc0SnNjJ9GGCtLaK0nD73HP7V14CZnkgwD7M3Ig8Bgpx6GHZoHNd5EUq07e5/rGFr
neYv0B8TUEXlmbM56g/NgMuDV4AzX47M/gMlFvZs+pKZ8L3QfwAViE0tOk+WvyIxxMnb4sPRZQTd
BhB2aVFJaV3eXBkR2EzNaGqHcgzlxIB5iDjG5pAFZwNp2poosoBC7hqt2aHWe9f/RvOGdc/J6tiy
bJOTJh/iq40fVY3F8PzlUmOJTiRHXrObyge94NdhJCewQuE+sPi/nH+HCP+tg1jLMQg/AG39aXv0
3f6vaxqJYiT+/ogExX2yfxEjcRL7k5EFNA85beYjaLkcBSUgyfnHY6eOqQQe4GMzzp0I2wRT49fY
sF8wYBEysqQVmEtZVhNAPkRp08TJ7s5FAoBuREweVL10HWc0+3Olmh5HzYvjOTG2xJ5Bydfvs5I8
fK1wSQ2SSa/XMrgAStnQGnAEf2loecPh8tLh7hILmFt9Zefg2fEoX+f6wd+fWgfBhyScppjPVVPd
PzHmAGCDr6PvKLPQ933/A5PBGo0IxX87G7IOcvBTEXeeePdqczlTX8VREkHos4yDYKi/E59VpaPc
iH/shXUZzkt0Sa3DlCfe4y902TX0hCAkUk1hl+1HEItpUgaLYdd5I2qyLwaAeD8x1CzhbE5yHfz7
sbIISxZjADgd/L5p+K3wrCS/YUkT5QvfMjve498dxJJTQ/399TBGtAhMChojG3msJ3eBr9qBfxBK
U7xSPICmBc1nr2Hor27Zg7TzkC8pcMEyUvqBEtBCpGTmNy2CPJXRmbyUyOq/y+m44w2IJcqy5sTU
KBdNxUmpYkMjIjXTJ34JB5ssoPks30i4JoalOwMB+dMqzwuwCoDYXiU5qXR+wtDKK7sG/47RLECG
oLL+MJLg2OpMqGjfsIzElEi1+NIeN/kJgsCYQWXcArs4FUnC0S9Il3I0L5kcSAf2UtGAt3SKo2vG
2LGZz4YXIuxact6tcMqn11oNa0OiOOw+UIujlJXKPGlRpgYgpAxBnzwyJQEdV93hkl3zcuNJt8Wp
O418JdfQ9KfFgNd+cZcwRrqqTv9E61ckizyu4uLB97oNB0Ji5I/U2XWWzIu/6RYOXeVaKbFqE5XU
UU5BHy1GRpPbhJ8KvamRw32b4xT3UnV2UY3IvsRG1Yyw84O89ED4xQraigVJqhr5PVHwTcVbWfh/
tHrilVY6vrXGwEqpcxVYSUqpm+gTEExCUY2l9P9EPW+A71R9H5GdZi45qhgkrLi1Gd1RVXxO9myL
1ZQmNSrxeWrfYWofqp2J7RJdgeIOegnFRPtH3phFJu3drC7Xgij2Lcn0qtS9/bUWz7XjEPe8/ed8
z5bkCMO9R0sHvuAtcSijXOFBbATvMgLtde5aPEdu0fDOxQVI9Vcv9UfSboFdm+YM5FFj1sgHq5Ej
Dmrc+6oC+7zV+67v+/XiAxF+6+d8xdAZgbOA+tf4dacXQShedrTMuh0Ei+vru/fzOOKfMXTXssPQ
AhoegHxFFpeLN/ndKdAr3x3yQd7oI7PfNV/E+cN7njbI2z0eqCqaj2q8Ub2rLL0o+TAs73sAuKDZ
NbSgiyrqqWEBzC75nf4b7tNoQJMQMIHNOCjcxLIpaPAauCxPgUxJrGssERZDAXGQOWqUk7wyH5/3
GiXdMsIJmxZc7cTSeh+DNK5rJyYKfYJrWbXce0PoYlfZG0WoICcTx1jMbhMfzJ0ASrW3zU+S12Sc
1ltsrVZBZeiZHHTorWgLgRd41xNzY1cRdQH6j4Ppz4kkf35mk/J/wr/TIypzicHBe4enhZ/DJEHc
t1Icz4cXDOIM9C42eFYnKD8yaErYubxM7JFA1KnPWlTOh46Rx5AohVxxv2WWQuuksYJqwEvKK8Ua
Aro5UKZFcRmtXdyQRtZl8FB+b3zjjz2vbKgCncO74Q7I5M9mpetQZGSYiIEV/ganERAFVNxIe7KI
gykEez8uN9orQiWK2Fw/ShKclhhwzV73wxebi4LiFCPUv7vHAbQx63W2ZL41jl3nwqRSVkVYR2p1
JbtRulp1YZKvBGhva/LTbZY2kDwMf96S92KGvPmD9/5k2GyDspUDZSkjeTfcC6eW5lGDZ8wp2h/3
zA0LdkGmIlr9fXsPGKs2uO/ES5caxaVzRY+PqR+mucqhQOaW0OJVfDqWz0VtCRrejF4ukKK6K78B
G7GtuWci9riqxrRkeAUxP8RVglxhaIc9ZEs8XiD+hxIn5cgwtUTmZChjtfxtiiyK/nBsi0Kvcc+d
sGujxtUrquswqjDys6xEWdh9QvXluorgYgm17lnQtDAcEEvOmaEXgwMPW91ad7A5vg6Ru8GEczRm
3syWYSv0d8qCU/3sAfuyhAGelIV6M0Tnv1n6K3x8iYFk66m96Q3+WXGKy6xhGNyqk5q7myRRefv7
zE1djtk3kIzLaHze7Ux8R1ug2PCz7mCiFjD9LiRHVAWiuRAZPCM6H+U84QLuXWC7StSRwwpmKwCb
Z1GRkrMgswap8MgGQdXhnTJGcuVgLmHjaeVAC3R+1ihYkvooTNEfYKRrr41w6iaO2ohlg7ll4kMK
YCAkcGXKd2SbjqgZcSdXvdDIGzL8mcDoAmq1kKxLDJe0Ay6+N931+jmrd4r2UITqVlAoUHwT3qB2
aC5u74l4jOsGk4M7nZhFdgxOgsGl88ok6B2qlolTUUabYi+2OmOQWyHHY12YfEsI2eIVG1ASiSDP
dL+5C9p6GRkiG/jpiqNYBYRoPlQFzf82vgk4Xq9p4pW/dnQpXDXTAMceir5eanni6tERQxHytjGL
P72imml+7nFKjqo1FbFixlosS63PJuT3maaOb3nrmpH7zklqNBBXWAnwWzcG2i8TBtao0aWXqjDb
gqU6+VJp1RnxDN1ftozyVFhbdJ2g3d08vxkgh686YwLLj7g599mxUPYAFltzjOjdzh27zPg4W6oU
LHml4V42O6oe+Q/xYNpvN9wedGsnBh07Nep8DfF4GoYS4mhDRWlAUYizN2cIICt3WsVT1oRpqPkV
jwsVmYlKQCjY2nCHTf3x5t/3KnA3l9fgEjqXcHEQxp6UJ1NKUrnRb389Xho+Jg3Sy6B0wy7h3g5T
sbTK8f5LZs1kpUwDBOBBCJRT93hsdI5XAKov2/khj1NgopTTN39yp25E2jkkU0AGKZbfIzDXv4BC
qduVyTeZ6nUYzTbD87nEFPXa/N+1exkjGxKZDTi6Sk44PSTHN8Ct8MADL1Vu88JHcnYYiLnH4A6I
HHs8W6ammKiuKFylXheweYeoVBYg9CEAx6/GDg5N1qUncMXez1JT5xzmwsimTg2GInQijvI6EEkx
7w8xc2ig7m8ZZSHaUx3UvxuByBhbRl7mw1tQeDe+2atCEKngy4vQgnbw4ctgEgk+wIkz/h/lZsxC
5trrpBHFp2GzjEnnNbgjfT9qPLni0rARSXJiNjyihTvIxj6I/beUMbNqVBQrD2vq2XaJEpiJNg6J
A3eN81Z7EOFxRb+LXPZlePj7CvdeNXrRzBz+Pr0fQbIEtshsEF84Z6yyjfjn38IKjp8HOB2eLBVO
5mRus38k1+eqV8IYM82oulb2CVr83SVynQiaYPEj5QHkRQ0vrWEgMp+GT0NSB+5VGa2vYqg3z9yZ
0BJLf79ifMOaczqN26HonEThTe7Bc0SkmJpOxjfpY2QMjddQpBH0d25dUDnKzDZKudrpEMZXH7TN
W30V7KpKm5KAFOOzSKSlPtv0jir6grP/6G8thF6G1uyLBkVMTxtCIshJOYiRYfFir0Jt27xh0PTF
/kF447Ntu2igQjB07BDRA+RPvoTVdd0PX7bTdYa5c9FpFIzpr2ZpEYLtmbXPIVYOmAHr3p9IG3cb
AnKz1lA1IdSNVG9ShZeLelGgF44HfS7UXA5zOnxdFqmjzy3lU8Jav59rifW45kntTeJk/XbmpTUF
vymfaMJUSG6rusQNtq6VaSVGU6G8xK42rlOIq+H5zldQHlI1JxQdqMJIcsKEmasXHIsH6qURLJgt
hrvbBZeuB2gBZGslIyfxzaMp40yqsY0U+R4EHahUYTy82EUn9fxcM3hTGCTSH4ni8+CkwwGhvji4
ETgu1oVzNT5fO9tPJknizUWufoXv+kRQvQyU8+9GyCpSPwejLma+dugOMpWvlfEuGdaMgn7Z3zg+
IlLCBRI1P9IbRiOgJ1lI452Y4gzC7e9d0eFMiWcrcJKsL/tlUD2ImvDIeIzNt0SrAxoGrwP5HLAX
s0Os2GtTcMlowBMkFqY9ZAdaoUf2mL6DvETliqC9sOWZNS5VFgm8mDtGVc14oHr0TaPsi/BlZ2Vk
kPZVgUof+9Zr5cvG176NkSfpnkS8r6VdR8dLDnH5edU+OaNqzlQRyGDx/BKcTinDZXAt3bOYYy0C
fzEmkrHXQ+vM3bsa2MihFeYP+xjaYyCQQAOY0SjRAFGw3NpUMR79sVh6cBGTvXrk5BL3zVUs79Ah
p1IYksDdJ5kcELD+RIn9/Cf1Dc9WNzYn8XWlF0y2276xKGDaBqmBTpsCf2vG0NwjalRjK0FZ4SRn
0v1e7sBYAst7o8+dVCq/hb/SZUcXxgPPjD7HWhNB7YuA8hhLJ+YFmx9IWWYd1HtuXcXzimkY4Kmf
yJlnwcxOBM/Ggwdekbd8xwQGKufiYtWz+oMIk/s66BSEdahDzJ/Hvp+BDpFJdrZeF4u4t7BTK/TA
I1SZG0h5gkJq71t24FIxGcDf7ua1DEDn87NM5kWl5/bHXB2D1X/xKOzaTdERuGLyiU91tNX0zL6k
3ejSaw4Vw/3yUCoBHP7zMT43OhAcwIKnpHkeYIZg44fGZwB6ZIY4rNldepNYl2Y7JlcBgux17ZX2
GwNWAQiJvHVbz2H06/H6KfR6+3bDEsvL9UUP5tZOIQVjE/vvuX4ArVulpglYrvJblQaHsnLimRJb
pgEoOpqq8imauLetwTukEjir18olqBFu468XHQTYHTDGCP4Uztq0oY6D0A0vUtsA320IK/BlZPJo
qT+kTX4IpER4C9PoT+Y3lRIuYisLG92ODe6ROjjFp/E4ukMysHIDQH7V6K8UiQNASv0JiPFZwneO
hdndFDuqlHUK+fHna+qYHKVWiYDlOzpwqoM79ZS1vvW5tpFwBKVRV8GS8Pq0YNGiYB/Ef0iCm/9a
6ZsNrPWRW6NvxLfVSKaecElhC3sqQbDkSondxHOB2fE4HBqwf/bXpe81tLA+4rQJHdel97dXBkpO
Z49CxKDediK/bhssTGhUE8lEeRlu2h7gBnpZR9MnLcna8W6Q6gX+nbkMgm6cP29rz3TlKn/V7fCm
GzOfV9wy7bE3zT8jK3K0Gk5PuUquALsU9oFPh13nvt+8l222cnDynU37Hk2TnZVAc35wJK4FKg03
UNXq5GusjimB99WnjRS7W3hmLEmtcEmahNWxG8dolhVjPKbsA9IyJSYuojw57xJq1wmxY66Yr+tX
OYEwCTxAb9dGZopUcVodxLtdZhlF1V3t/40ad4ieS42tSInJ+STBi+L8bsEYhjxNQK++elbjK191
basHWP4tVSXabNdn4xaTkqtYJoQsNTo98AhVY0GnqA0ZDoZ6WGcdbA/j15fza7TRe0zzmNxaqvrS
Umb/3D5z3ODIj+fcDnR9zDIijii41p/uWIo7rYkPOfVTzSaGMUjtvplVp6kWqHMJM5Aj5QKuBHs0
3WwkRYzd4Oyu1DxdkYlpaHRcRtZEb5KKXwXl27r7YaX2swl+0AJUlkmUifmDAwlRzXA79NATfM8F
ppj+phJRTz9geG4ufR9E/fjm0idBBdUvqi3DDvH/8dCB0M5D/0egtNOuIirMcD7YAbGJibp8zMZ9
pcKi0t8wn3dkC9+TH7sV0yetUHXPxnb8pvNyRUBAWCfvPWD9Spb2hEtW31nbQJuQBWbgjAHW2b+F
A5Ctk3AQP9l8CAx3MgpYwn9yOtB/FKueJh4q2ssz3EINRSJH7yg6ljn2O2w4A+u7sJzxKqp44igP
vfxRF0imJnGpJgKrKEwKdtJMccVHvQ6qugwv69AmS0AKEBCiJRG4QxK0hMLbSyPDsz81PAPUxv3V
5rEsfMRWvzR59aHG5UVLjYlbj3LbbAkgAsRO/gtxL+kk1Hi3cF5qN474wsivMnybyX2b0nJKctTV
RWRxEwEaoX1HWCZKgOgONAux35w3/a/nwwEnRZM17gi6GQLCl/Luzh5+xDydf0N+fsjnl72Rv3H5
uG1A9VVFKM5XTJGJBY58nyXm/E8CtrsnDPbL0Z8gv6zUMFBO2wOY6caXNEwYUkBaNTNrYw9g3hyl
GrbhAvPS9LRcj7jo0v7g0LioHMooW7fWPwkeTscDg+UOCqoSFw7OpvdRwaUHYzWsvlg7IKmWzfsJ
FeyFTAEQcrhW4RVpDVZWR6NDXVY0YYA2nS4TNOXJx5x7HlJQ7OQlSBjacrrIkBeUSemnPQZAdc58
kuNJwvVFyk8E8y5NPFEmpGssXXL/aH+IE9fsjcjW+xFOLkiJG2zHmSqobpp61vLxXexNj0Y5jBcQ
YusFI4fSzmOImUQmSJIsUxZV6oWNl+ZW+5vxuJ/lnIM3+gO/nAKFR7LXnlDK+yKKR9XKk/e0FlxV
9kyCXI2be72kuBqou7XpDre+aIqDWBi53zBppefgO0BLaRs1h9GazCRbM4x/a3SePgpe5S9iEzmC
/n3jyK67r1+DxMMxF/GoABK6WpwDXENpbW+AKsUY1Xh0T1QpF5otnF3L6kVg43GvJR/BkMyg2kHQ
QUlBgcu55bqnvx4joVeu30XGZfLq0zUVFfygA/W2xmFUv7a3xWahgtPmgA1txJiOYFcluiyqyysp
aQ+6Fy/Izf1wNg7hDkbgxT8CtXOJPnsBmWT3zrfCTLqwtO16hQnDS8tiLpMwZzUsu0NAl7qGg8xn
Kx6gPkd0jQ+I277edKt6f80oGalbDKqJHG+DtFhg7CtEPWorN4jWc4cgIy0lVx9hFZ/6H/wwALFz
C4twA6LOP2eMAYtebz49jJnQeqsOr6AN75Nsoz729aRUqfph3N7PKIkzOw0nggQuBHAIuRS8ASHI
fx8wMyEZ7sqzZ0NdDDKmLfn5PBpzn4RB+2uG7Z28LM75cYsu7eJYMeRYS+LPxht/cqsiwXsUmc8e
CSGGwtn7xHiM2tPve2l3FE9A/3IH66OMAgr399cwJhKwgluq49+fJ/q4+v45hBYtGR4rhxG4cbBu
/S88CyV0E7EHhiawJe7qSSOuY/KOpsm4fyew8Qm+h7/9k7MN5WkPeTMAcG/RAW9WBmMhbjnQeMd1
PC1idRaBXb7bqHVuZHDVmbtPv9tHI0rk8nt8j9/Cgi3opZFtd3nRuwS3SzKuXZ2/j0Z7CUvJWNfI
iQl/WXJyGQJoO7fl5w+hNonfmt8NKGDCwgfxsnc1cN0JJZhQSB02SwHwZFw1E14CL6LMWuPO+/gc
qT58yHSVK3Wff/yZUKaaDMGLnIderXS2pfD5+uUaS9+4/nffEBacHCM/WtWF4jeG4p9cqhDHHJWU
FJNE1f/0t+Zb/PCS5274eScEsRBVSBqwjF63FggIzS5zDTxmTU781NZTtyQ/PduhDVxogI1DhSef
4mE/0CS/2GNMXl15YIsYN6jzO5uhkSf8iiNNSShH2hskZST5/9QFBrJalnrCXHeVg4Yb17cURrY+
vBnUMbYG7g2jlhf8WxXz7K2maDuAeBjcoQaeyjkHBjOJ0kgbjCxolBOQTKU5ia3saY42O3Vkto6/
rbkUtFDL68CarEy55V9CH4fVGc9CiAnnUpb8jXkSNjzj2b9LtVIFhcn6yT3kPYsNgWI1kb7jzAGv
K3T5ydzQ3bah5yi24brVw/HntQKkIr8tmBn1EVrVAs6SJ9Zfpr3K4wUw3qUQvXHXsXgFgI7I7Lbd
E61uWSfDwMEC8Iwdm2tZgMHrOmSUf5OYaUVA4XMnhImJFcFkdQtrl/q06mHQBN1cPI4aTWCyn0N8
LOE3AmkD//s4stV+dJwwP7FvYAm4Wx0+Hhu/mnvDi5Ynx4VbrELRqhuFriVxyYtgllnssJVjj/AP
/zO+A0DIuZJikUsSyQBCGUO2ZkXYH+Qo61fbR+grL7ukmUrwthEnfYIO8Cj+xZFwMQvVr66uLsmx
OxHUZizdy7t8XMmb4sOym83COgenxqXqDGFp8ukCI++iRO78p679rv1q3Gvy9x6hL4ZzO+ecDNIc
WL6Us23PJPoo7WV0zEpLTC1/lZAkWPNmgeB+sp+l2DLI5ylHXf6nbyesuCxvDiB1VpQDbEh6rc6M
eCAYyDCmPKhUcB1kQrjXMBZ8kMhLnSbuuziL07GM6N8ZYj9ShnHCmD72wsicHM3yXksIMDhvgyO6
//k4x/rMPQvjVA7V50x+jbmyM3SY0TPaVDXkcnXN8sps4Zf++5s7uDHZCWluDLGM64pbFb4+5ROq
IeQ6yqwfyGwPYWaJlGuoXXXRY0D7z+qBTDvldqDem1F5EIVJr7jp6GWHazzI+911795iWkB1yAgF
4j3LWRSNL11En0W8sIrShsLWSSyOT4EIGUjvZV9Ijf8zITXLdlc/mec09rcsgcXRqGokjDy8tRFm
ilMxgSMbJsxTUt9dJnaPYeYA0MerGcZABhOOAepe6c+qJJjuxKXy3feJS8iv0BUusBsALqcQInY7
xFlKwFf2W7JA4atiytLuTaCWg5n0hG6t96oo8FVQaW6OZ4Mx85q00AcwUIQG0WlwTKfmMu5QuAe2
EzHO8tDWaMkgfiJaLkAoLJt6RafG9UM5ZVVCozetOXrvLdg53d8VoeXVIx27yYD8GNuuFNu7ek23
1/GlF5da59IoNhx6F/1TA5a8LqxvigwwqptJxALqdLsfmzwJ2iHwKqHX+nDPJoCmVT6maiwTCeuL
SfvGeoaOehrJmLbu6rOL56Ds5RBuigTC+KhqksjndfomDLxIEoQy5Ty0Xqx7heAu/pHden96UFR5
k/BjDrlQEbKvRk99NOYo0CsX0HBtCcD0wT1hAccd9K9rPkc4cKs0m7zWIQB9vWKT+53JQ/GwtwLY
hChQexasm4J7FAqvM5lfPsv6FwLw9k7RMaUesnfoMenJ30qzFJgjAgn3B+bhViWcaII8L6XB4DW0
MyGab0G/6CpQGEYdPfCSqKw0OeB3Y2DbFnvBW81+YPb0X++ZvfwUEceBUweK0LDOi28INF/5C1+4
jNN53uEL1JH+4ZpKSn5MABnItgw0o6nVFj4y7u4D3AsYmfY9zHEtiNiftPbIWlFcHsDbd/n1wjoE
MDXbbKF7PefUxAhH0aodSXaiCkqjTnkcLJqtvEVActbSgd8a2udFIT9si1gN0A+qzSUAApo3SJUI
Iw5OmuY8N59yzMdiRIJ796lPiAqnWIpaGt12hEShW6RFHDKMF/RjF+hmUzf+ca+mZDLhGTur8oBc
ACOLviroOW6+n8rZ8evpy5KMGhcsep8taqLriJd+VUMDTr8uIjTTnDKtg+W//cNOy2qXaaY/wzBP
/K8aeuSaEC0ShWszbt6maLbk8+2E2li/K6L+dPTBlhHYRE+B5SHzl05mKGf+Tl9tcZMdsjEFS+HB
4ghp7+cEZqPJwIi9/1hs3rfCqx6C2a42e6Zi3Yx9+HkukjHzuNEYLCNZPLQ2+0C/MZIeN2ZmCRw+
c+Bgi/yAn6DO7WGPyQmcbrSDGywlnugFMzfUF3Tcitl8FOjLep1DNsckj/9Jn/FHm8tW4Sk8hLJv
mOTgsbs7VddK3lIfz6pbnGnOgzTqUrXAk9ytCsVe+VnQtmu3yzez9SdmkceVyhFbnhE1/UktVN7a
PeYDTK7kMre0r3+Dqi/mrGSKQmtY93vwRc/JA8WWovkKyCiHXQAeaN3hZnNbdDKXCr4JiTyR2zId
HyH0XOI+E7o+h/gDNDZm4JJs1VXxz5GSw4qZLKoRnM4dWSk4ep+APg5cn+du+xSIxGeb9O1l8i2W
1kA7VpG6z07NpwyXbxe3tNLZfU+XumYk5TrW4an/pTghj6gMEdnuaJRhZJ41GRIsgM95l7DMojEJ
BAWXRthzbQQKHPh5fYbhE32y+Fu3KYuxSrFKht+CjPWNJ7m5a51yJzMmrFyVjLMYoJni83BNOwGu
E3CLcZKw0GU12ocTY60S0327RGo7btFh3pyJGnrxgBkSo7DJuAsRwEbRZfH+WJjUHpfuu2tzhPdH
1cZIgXlNy1MNZ/l8Rco3Vnnq4HAJ6Ib8EiJ/Qy3M4aO3zgLrAB+12S3dQ3AWW7Rp8A7pvStQeDT/
Zt9+kN5nxlJTrIg9jHWsX8mYTQ70XgWBmi8dp1WuKuPYUAA0g6HZ9Bc7QRU7mJO8hvj7qFoklhiu
JLr2nRXJ0l22+Y8KhoMpeLQIG1D+nj1mZaiWtldYNPdfF6AGrEk8UFXfxueLPCns5K0aV5m51NLq
PqGuA9Eg6KXAToH0yvbr/+4THRZk5WG2InKTy9fNWRSqu2tZ0yjG3NE8MpGefjFKP2S+kAch+XW/
Z5P5k+ZDtp4qnDZIkAu400OzfTEisdGraQ0gAIKI6APoSZyv/iZfvGbhU5dRa9R4MpDGl1ooGmr3
BFMSlGwe8iEBzzP45Xc26MWb2HCdak58Eg64UnGBPVctmaLUZQKfX2nKSBUgAMrCsPEkAgoFgxeO
1Pfino7CouVrar3gozCRRY2CJotuU4iTZOQ/X2RTSdxaVigMpLebwTa+D/ibPLt9rT+xGwRs29QK
SEbqe8z/oxPdbbiiMgW67R6kxvLlZ4L3vhHuIouMDqO+fkxpe9NPVlC9mjq7QNuzkqcmJj5GKQgk
8RmNmW6L/w5HqePf5v+fkQcgd4FLKJ4X6hW9lAOd+Q4ISMHv7xFi6A0sXLcNtgfVIbouL6cgOXGZ
PcsiwkK/LWUGuh5eTcVfHZEnvDWkp4iHcxDzQBzQJnJ1QuMwPpleV0n7Q2E5/zQoZDhuuIf+9ix1
SS1HxMFLzkdbg+ZLtcjV7KUOgCV0OjJnOt8921G9CQ32pQZ1KPajxenuJKdWSq0b7W8P80NWP87V
pxUanai43TfxW+Zyj/OZDmXMKBLQuaC0P7kkWPynSEn0fh5LNM3R7iBqjdeg/FDD8x+8lfhMsAtv
sI24j4iJ/18fjFLRIsaR2luB9npUtiJ6xxlO1nsROsAWM5mYtwyu1Y1Fg0Gjqn8LLZ5nCtRXwI4a
iGSPbx5YN9HEPmVSPy57ru3qyneXFKGJiboIEBM75bvPbFenn+6KpIlK3jcQ5CsRk9hE5hDic3Ra
Tq4qviGKJue66Ru3APLdlHqnQkbmxh0rU6I8V4DGj3ZyemHPxbCZI6Zi3piu9TAhqQg4J8SHT451
FDwSTrWhWB5UgxYQZ7RN7Zw3IpPMjTznbswO55UbcNZbSO46SnwS7HzHnRDMcx4mQw5ovDOuwYKU
D2aSqVvAFx41cpSc0UCnIM+1al0L/Z9o+3Kjou0dj+qeENWqj1+ZkTySHI7/qTP3S4r+5LvJBzHN
8sodyDRjrrm9esZPjujPRwzeZe6Wyg4D1i5rRmjAli1qO5PhfSm4PmEKJtPpSWBFURxPtrw4ayHd
jWVIQRPJ5JpGmjQWLb1Ra3M8XWX61QlKCHpKN+r/PCegJwhtmnTzYNuW/p5+AOrJ37n6oYeCuSK/
fma7Uq+pZho1fG5aTriiorNZ29t4p0pWovlsViWiIuVQV37jbpIMJLzCW5UcHjUi0a4moJ7sM0ly
0K15srpN4WC8asja70JMVoXoPEIuHnsu+/8aVO1wSVOgtBvCW4uqOGxHSu/zxWqelJinm/UHBW8p
i2IiD1Vldq4Sjo6OZZgqrN0gYciX3FFubBCJTOG3CLnB44/QYbfIq9iDZtoaMPDUD9nyheJeDnG1
Mj18cmhC94hchKfFMXpM5qeW7RxpAMai1iuxqadwWhRT7ajkVjpJPd7c/RnEw3EF8cYwuwP2RZiO
mAul0UI6S8KEZS8AsguoMsDVV/MCFGJmFopMNEtJUHxzlzNfeojEjCOTu3fgRHxO3MG4QpeFFGyg
2uQFTP9CdSGTCrBMbfiCrINrsLTZKLkDXH1SYwlAaEXqab6PiukFrhjGSseHWQ9E7Anrkw4zf1YX
qMbAzhoAitOXkpolzwiXYkhz21bT+4A5VHuFC5neMIcVQFvTeizlQULv0ER4ERFatFqoQV8/25jR
Eyglcn3vJ6vArF4ckNS3cxtBorRR0cZOa2DGmxDGD0PDKMs+/jPMlERG5Vp3UBOL8kX65bw1ON4V
iHZfEQvPTFdxAyefY20xyah4N8F02vdg5AviYizBVhy0aMoaDF75zU5BwTvHsFK5mqP85NsvSGff
5c1fSmnrvhvl+5N3332skcFgp5Ua4V+Z7+uo2H8Df+BqvAvq0LAPjA7unf5lgM4W0bMZhAN4p+tS
zrQEhJ8SPOe4UoXAM06vqxmUgTx739FqII/Xyv++L2a06M/EqEfJM+kkOnUSI4JxcOQPJUwrXt4L
fe/OOlhGdg05NFl+I07y3mmFRswthL8njTSWeIOm0gf5Im5n2+pGBJyhtOqNVf1gbZHo4r9HBCi7
524QGb9TpiPmaLvR2jLcGPq6YJNYXtswKJXYrH3MUKV17VgiZe9efRDpKcfEqooA4JYAvseqZZhN
buWixETcO9gZq3xMGxZXZow9GKg9Vszt8cvenJNICMivSzqm1oGigRjD2sVuo6gyWFahSVeciXVF
siNH5hLQGKGQ6YcBbX9wXc/0uvl5roV26+KpuI10synuvRwFy2n21GbsngAFEiIu/xARUHN7lXta
ZX6i5bFmRDf5v9ss657XJE7vQWdsjs6j0+9GM4oZd0S6I5C7yzqeAJh47knOSsVxZtZcIwrQcZrI
bbBPCFd1fh7cf0GyX771+OEozXpmrHP4LAjeLjLV9JM8tbu6AXGHffl/7XvtVFLAEDGEklzuKfAo
WTEY1zpp2QzwOZapGoCAa9VAGfhIUhutCeFCaAWgChbhoV1bjwLKZnjNEFRei2SJh6a9PUtyghfX
9wir2xDzb4Ha6r7SUivHTICoEvtN8Wog4aRU0If0Y/GoJGrtwwl5adzVi43SSaeqLTUQ+VhPQozN
HqiNdpxZc02BltmaR0khX+c6qdZ9JcOxTu+Xpe+a4u/dpeOeC0ALfKmSS14kjzrPSUSO6DlKG9tL
vHBx07FrBpgt+OjgqV//HnQwVz46zyGy1czGRI2eR9hi0g1AD4gciqTZZDowOEAm61/AcXs/Qvz0
zhBI8YIcY/+Y4CjKcgcxiMpEa6qCfq58Vc+0Qz+exYuvBTLm5r8juEitDQozD7norrDbC5KYThM0
t2KFNzTnLvsX93aUCrhQ1HatmZOtKzP3lqQZEp5W9ZJKcj01ArU0MZa2jrkxxMvnPdz+gftAfBLI
HKXUeOCX7KKnwDGoSte/o8oCEQKst/0lhRzOBchiTMWwVIMg21bQwiGM8YHXqpfg5B1NjumRZx37
YJ9vevuhqmpl18IrWyZ81+12AnApXwHAcbDWf69c696hEtkxy0x1CTwzP/+zLjuLQcgulH+i3TaA
7gO9Jf1EEIrnEaIibSVWYLClmvR/e6j5h3Nst9luagk3Lej8qiLmaBdm4MZV1Df+NdUqs/LmHrww
QenEbN0dMXNUZA0z68oU9Crx5NM6N3xnxJvBpNPnEvotqGYDuZFO944BFUwdwN60Aay+Y+uhzw1X
Gpeig1/RlzbDPjHqzJhxhu0OcGlsNkPdB5wFXuAlPs0CgupfxHn26tgnHpNUKemCPoWfr0AmF3v3
oexHBF4OXSpw/9TZ/EQo8XA3PeFJGQEPw4GKdMJUPc2Xt/J2iFXjLILHlVBj7vXNbQVQuhh8rIlz
nLmlC4JoC6CTk2lef3Sqr4DiDo8mh1B5xSEX7lHxcitLmEcHAMQvJ6sWssqgBWEf33AeIRUV+owv
Rw9B8svWOkuXeocwgFsA1oJ16oRPgOFkmC1LC0rFfqWnxkfq0S3ua4U8dgvBMtUXuufjzmGPHlDC
17JP+r1wiNNrHrIULg4pSUefMd4cDOkmdYSbO3g2Q7NOREcsLxWmPJOSkqgjFx+376+EnBy2hQCB
Q2bOqiyYg9LLCLMzXCrTVclcJp8sfNIcdq3OB82oH1Q7jOlh2g+Yc3dcK8wk3lV7qqKUgeK8iAoP
iNpyQe6HbQwO1jC0jq64O9fW38pAMcxC26ZEiVDNEhBVDDbM/65qTI7XI1imducmlyjtA96u2Bcb
HDdwqzCiwUf7zSR3spOhORUzX4j+89dNRI5CXYMSF+URUKOkp0YKc7bW+fhx2qDdSYZONRDx/8VC
sfnuJNuZPjy5QOLQ4pdKRl3pK7wg1zBsIq8dyqnOtPnBao+w3NtnABkJgq0Plf4pYyjql9awMrK0
K7a93wxVoOcPWQScNNR26I4NFe6KdAr5u8x2J2lEADh7utmn26cLWQWMJMGyeyuvo8xHLj9Ce+sw
xmLv6mkj7mis2Pjt9bqMyV5JZZSy8Dg6EKKwLwajKWJ2fSAXMtYI4EV6MUv7vpIO64XiyH72Zkk3
+bkFw0mKa8bxtxHVmCEqjHoB1XX/Il3LUKaC1uvX/E5clwDyf3zzNP53uBFQn2vMq61YzXkD0PkT
EjldQJ9JbOcTt2GOUFpCc/P3YKoR5RQuMt+RKJw6gRZFwAkK7WdUMFCfnEEoJOIEaEO/sMgerp+t
HTGI5FLojP/fct4OI35nNeWGW3o+IIFRXTbJFoUMr/+Bzmsi0eQyTdpSAsU+30OQEArixUsGd+1c
ltOcyIpTafuzkj/CCyIA0/W6ULRix1Tq6hxa0JD794EzYGErtw0TxWef61+IDAl8ZeuVIUuZWRxd
hBhV+6d1tARQo/lL8UQLY2BPCu8X5udYVBp4k1gPyR8vQ6bNz1sRDKma4dEu7JJgQJ0RZ08NYc8s
yHEVpUs8QLPyb/qdLGAfYBkHzNmQjC6MQeHvVjIw1UsR5B8p9zx8pwMcD3K3UDkzK7xL2WBM+aTN
ZWlAa2Ff1qkLOOlqGg/mxC8ACdMBnpbAIwg10xhxvVR0coTyaPBKwTZ4U287XUXbruR7x5ilMeoe
4iOBQKccpjBLm+QxAvQUZfDNyq8DnJXs+cnVKj+Nd60kGddl6L/nTpAgftjXkXTOR/uhjhLvzMWK
v+IUNlM8XyxDe+ncJl7uWw9EWuuKiiD0BF4eSRLfUEd8njAZPorExBnKxlGYzYJ/+k6jnN3w48pt
v4nqBIaEEBY+Sm5U4TyWXOzyMHjoWVr7/QkDbo+bH+KGDN6pT9sFz5932RoauRsSZNRvOymancDO
A4NLeWf+C2WCo0/w9UIZYZPSvFVUyEHTqe+NffN+kbQ0bbL+aedr4zK/7bzY8q8yskKzp/x3nfbB
o/ZSxfBa1ghOT8qe7CW2Fy/ApIIcOeh5/MmyCz8Z5nQF6WisO92IJ7e32ZqzQopEdu5fUsd3DMbU
M7eiTvLu4pyqt9dKtWCgHPoMy7PUB7Qm092f2iGOvMwHB49AB2dTYzWHDNetJ34LKYDmOwwGugFX
JP564SyaxJdSayNG6eRpTquMJxFG2EPkRFViw2UD7Ne7Hgi717Dw2q/cg4pDlZ5muoz9G+IhNoyj
xSV+J+6qecM4EU1nzAzumlZHsnU+8DBsXK7xPbbEEconKi4fNGbkk5Y4u8BfrArb4BVu952imm2R
UwI786KZmCM2dcoXGtN+4ZFpJFbObQ2EtXn86aV2YERwNYS9mjfxKrFOL2WKmlAMJQGovz+2DhWr
QGR4U0ZtG/xeeIiQR69t3eZgJwo9oq/1wYAJCDP7T3h11J0v7yzWmOASdXTa7b7EFDWbpJcU5uvN
mK8xovVirwBUJCjocN9KRK3CW3YX3KEV+7H+l4c08MFAu6or3ZikfCzy3ALXK12pOQo8XPiUf4fR
pxPRDoBJFpkTtIdMyS8t8QjRjJBZbqBYUe3+eLz3yYB4tp8TQ7cdbTrttHDfTIPLi63tMjCn6QFx
9lQbijjC8abNJcNNdiLkUO0EsKAw6vifo6WEE+c+s6H12Qve9w7tXao30TZ+SwXrDi2RKIIZ7B1x
4j4mvheJXd5oSqFFlbRT/Q2rr2mVcvKG1Kf6+eP7Zx1WxLJn0BiDl3YTZ31+N1Y2R0Bi0aPEtWNE
K1nJeOBCpdEtrsKeuB28OS9/bZTuDL113Gc2KLJBDcuJnSEtO0PxNgzw4ah43J0HFthGephLwlDr
9FFb0ZKLItXbRFgmkbE+qoyUPXU7dDZuY480RLhhgnevRWs23yyvW3WH57WtDSpCVN0tTtxBmIn9
/Gt2IkIqayCGkiqsqNb9xan8ZGp6XxIh3hzKwfay1sFekIcRmwVVcUMFc/wEA8nRGgjTGm775gA3
3FqXxEXJM+o/kiutYmzZT6T+n+wjhlI60TUrPvtp8imkq5cuxS3MDl1LIB1spOwQTIQVRG/Muqvq
l/AxSMrY7Ah4IOr2WrmjZi9vIuo0lr0S2rhtMMSWTiZjnmjOHbBz0dZ543LqBwbHLPUj6UURrIM+
GplmJW4oprQCsUoHZrywzNG3lhOYqPOPWloVCgfGPHegWCC1IOb6CT3XqjJeJqJ/YGzo4sZ0i+DU
azylTOTDDusuSmBarcfR7VfZG0hmcGlIIcor5whRxMSeztk0+gG73RqwPyOm7zlBzjCWFVIaoTeh
Izucf985UGRcuTXlNdL5UCgvvzhPjtxYijVDU0QsTh1Ln34TKI5RaDFSYw0TnLiembXfCkM+eWsJ
X8Uo/uLlipD3f9hl/4JTXGxmU2I4ZeLNzq6htHg8+f8uP2/DIXri7O+vI4GbRDHktzuGjlt7GkkW
X4WuJ4zNBuQK0sI17UCiAjzJxodCAncSe9uXuJfczpCrhsKVDjX0zJEDvWxJuH9m0D6QGIizFCGF
eeLxSdVVFjM1DmO2bhKrxxqsBrb+AR2P4WswqeVYVulGteuk1HbOASdpdOhQCkzGvdBDf9TrvfBN
NqEgPQaRpNB7icjuFrcmWeYTmPZnFlXQNKHTV0xBbgil2vQj+mtMkKejhY+x1EDgvrp/zvMJGTdV
bdeSmJLYXa0Axq7aQe1vjk7EDbuM8HtbBNdVXvRLUWBvSGHqW2FDRMDIGjJxKIemRyRCwNO/n1Ug
jKJRp1tvztLPkXGzcWzr3qItnliq/g+my+uN8BO1A7RwKnZClBMz9MnhDoaVB8nVxuYS66AlhDmh
q95j59yJN7O0GSQp+9FEfpjJgBobxlX06wUC3N0BY+ErOC29xOH+9dt9+bsGMA5U1qJoUvV/RTXr
EvN3NHTP3R0fSeLKVvI2PfDwCqhbWcYOOoYFs9sf5BE1e/7aTJhsPIGHhf1FTrMN61Tv9Ir07cLF
5XWNPFwn3ONDKscwqS+6kxV5qjXEr3NjyAyRnDF5Px1FVcslvxR26eDTOh6URftBt+XCx/yUgyLn
yGhy5VNDM6ee0VgNbvplGj1B36f810MST217byZimhv0kvqyvh9JPs6gGyKpzPz/+/zYgSnKjrdR
HwQke4wumYTJmXN6NNTNHjclfKwFdSInrd3mGEdh7YV+TH+6v35EM4lSBNU8Qsp6pF9HLNiaJ/UQ
KuunYthTLZjLhvSOfMs9TcL+xgTlY1NugXfuELy1AXQYuyYWlmlQEQ7F0rAR5JreKcpXsAIYv5zN
AGc1xjwmFWbrbadHRB8lJURwnhkSCvFcAM8bGTxZmfFQ2qIzGEKTvywlATvXzALFgw9DgF5bAvCu
V6QiZD43jzd7GPxaOp+c2mxDX3xFlib7UdI6C5tavfdj/J3KRXGhPpOu80rpQqEZtgBGI/OeZZli
SIYYAOOdlXX6/NfyWh145XB7kTXw7P+y9POpV7TAIS14NTPOJmvEKZrBzj7kywObSiZcJKSkBI0b
y2ns3kC3H/McxyBj1bNMCQOiidOuqTbLAL8RDciJKQvAJw5u9aym+Wfa6FdssBdcRwb3c7bQqbjB
PkROG45ImbmwKgow2+T8wV9TLoF0d136wi0OQAn4xTxSmH8zXhmyOu8OoO4GVHfiHaZW+zJidfPE
9yfIkUlnrzNZl+5/smRVtkslxca3XcIgHg+6hFx5BWuCTrSHrtInvMnDaetVnGQoRbK2wY6mFwO1
Oc+dOCzQjDL3grf59V41mfkt1kekN3mFrWpm6VDF+9yYFF3uuj5X0wQRfu7C8p5wPnlXpGOi0skZ
avjr7u+NbP5iqGzpPvUWhPisT4mIa30jWhu9qmXIuiLTX4n6FSljQw7f+C24CY696H3xi4vCcfAA
ycxWlRrgOln81MB/1tV+dlVBbx/8Cdiw+8UMrbntKuKpHxBQtbsU/YGZhnr2MseV1v57q9aRTme8
7ELnjeBVfgtO4c2zFIz6oHTGudUQuzlQ8b54gT2ZfcPcXN4a1gm/xdHDwD+DSRzfI4T/IWlI4qqa
pGwyt8oh2ly9J+Ms4KTSrD8n0x16Hd6zCbN+9Jj0YjVa7NXrIBGuu4gF7kyAimr7HXAXr6UReZYz
2zxVKzIUMsCMcVWH485LKj3wjQvwXa5431bkrpZExsVg4cN8QDwWQ5YRexLdySrJbPqqKsNanmaY
cBSmkINJzQPKD4FeUd7WRzJFMtt/poxmwZtw/E6n9A4eqjyXmiXDBeAMWM+t6wx1uiEohlp5GF+O
/ZaBkghG7PREJVtmrQfkexJ+0hSUU9Itd/9vtJ/UGYFwzFBwg+kcs3EumFqrzx9/nLE9LvWZ1Q/a
MWtmLwuB1cY2jIESXEYMcSCDZRamln6Ewj/1j3d94AmeQ2hmsEYDAfPQhNLk1j9wlur1Fc105trl
tlCa7r0s2h2NA5BIp5oHbd/+fqcgiwBQrdt/hnQLwMOkgblDZTeUJqrpmbngifguv5YG9kH7wEjX
r9f/kDJEmt6WFlJAFqnG2vUzV0EfNSbohRkyHtcxe3NvsrVaCYCQHVdwOdYF0rwj7zWZBNPeddx/
hpMxZUArrdPozzEuLBb9hxUClXAirEeYBXC1p+2cI20NYiUBok2EqknzYNnosxlxFGXMJ5iJBFz7
uN8zKbap5rxxWGoqTH/nYPvkBQzthDL507gRizUOhZublXgVDfYfltIylMPhuDeU9VNKCvF+FVOn
xeZZs+ilJvbJoMWjiDQvb4NtPVgopQqiU7daGJGmItPlSmQf5pdUKQPwErt7EoYPxSpN9b2Gcdm5
BK4a2epYi6O3jBol/rolvJvepJ3zQSST6NY8SneKHkKOz1oH9oJXBS2ixliMZH8bCqaIWI/SQMeL
NsrD13HbjA6KCdNZvMcQtLwi1sY5Ctqu/yNkoCa/x2TtXI15H2KtOTd6QRXuu/pZ7/sxnXqU21kd
wK1sUHwRoytsBdZcJWRDjSWX+KvghtBGgysVg6KJzpiAN6nRVFCvxmUbkR5lV1xGpwEJ2AVsYYTf
c0gSuopFG8uzyQZTiHCJ1IWwOsliUroDsiSiQSJJIa9L6ZxI+mwM/BxALQhnei+XR23ui7NXzm/I
IBDI4rBwh9OXgMVqRFeG0LA58f2YKwET4RA2VNh6tnAH50Zg+Fl0T6ezMl3NZuRrP6yzwVyawzm2
nbGGqzaacJpFvbv19uuNTWf9vM6WKrKzaBu0Rcd+e6igw0iGgsHxzMxsptQhAsSOvYsfX7W11HRq
fLlbc2uf4h95Twjuxt6fbQLOWHyTfLgVxGzhKaEgUxUgNQLRxIh8eruoBsSsEkBhyC1FqsLV7Grd
tdhDX6BV/jMwaljMpc85yPpbiPzbUvjjWliAFnRv5hpRhKsIvqV69/F4ERG6z6hkZpF7dgm8Od5W
JYa5/+t5NeBy7bSRisi13Uqrt6hSXMzBzGnCsG91L7jA/lrhXunw+iKr3INIH0tYoUqcAYv5huQQ
HSJ6B8QIsWDXobqNjMnnh9ujw3hBIOGaxBGgOOkd4H1hBmLjFr/S0u2Ct4YQ6mSZ+70rHut9iq8w
MJ++vExnR0OIyHke0W+yGqxl4wsbC3nwbZR3aQpRWsGea+jw7feSY/Gu1XIOM44EYFMkTKjnqehr
iopitjIBC0s9/pkmX9fbKfLGyLlYopY7JG3hcPOHpBK56eYMCnOwRuzv1PQJu7zx+aZ0bygXpzmD
4KuqWHqonhMK0ntMC6sB7PGW9whIERz/vrO0ljEvKbLmZOrOCWrdh2jWvgdUC52C+s7NG5InwOc8
JHwvRzldOh1DlwDDg70lCAN6l7QPdDFZOl4leS7SL/u56kKQj8UOP64QUJpmbziE7AWt5QNN4/0T
+u/9e57wEATeSNIM+svaCoc9X7PD6iCwMwQrcAPEchSX5VaWfRfm9JGtC+adIgF2AmntDr8ak4A4
8mMTMgAqsAlcJ90yUibcvCXuHMadWl1PTCMIKcGQPl2PF3OPHJi39xmdwVIS3RDIQbGEi3MxO0aR
cRVfxpSZkDk5meS4aSx76fpZ/x7Wa3yPW2ro4s9hQLktcWN1ltBFGubxTGyh8nOU8DoI/kpNru2c
lpeBC6tlAGm3WdVWwwpoty+jERwJDP6Ht2PWzKWtpyL32xuZX9/7etlkPZOJFKIHGjh0gxCLLPe0
ryHGankLUDm9BgOZYzB/Nnsx73Vleu3iLideafINkHW1w3lDH/t2pahxoPbUvzkKGzPPOesIM6EI
ryC6o7KV3KFfsXVYdrShOKg88N0nP//L5RWnnLdxmVlk7wJOhHE8Q8JTN7PP/LdBPXASWEdUvqC5
ea9U8KDdkd63oJ5Z893RXVsKV9WqAP9Kfhgi4IL9J7Eh7mICcfk9atwap4dsiDTsWuYrmjEdO+E3
uQFJ2QcNMejb3pGB+5s5XBkRIMQnwx05KyiO8jEvQ1G2dBzvVl+Gt04G+wZ/hx+LiP+gQIVBm+Wk
Z5EJi1y3I3w1OpzaVhYE5sENSkpJJyLilBgHyn25ZtiA4/yBDXC7v11DUJDYCQQiDiNwvBS6zJsD
RnraGyweoDFDXJypcPl3P8B1v7yqzIoIEK8rypzo7pA4PVa9+kUPu2A60moSnE66mOVzoJbHYvtg
J6rnVfUq8DlEoO6DC5iYB6sa/V1aahji07q+V6xgcfG5P0itNWI6adhHIJmSE4tq0YVIHWzz5Fqz
pAwZcB1fj7hBiX0V0eCYaWWG4jmK/oko6QTRwpqQP0p5hw510v+DmPxJoNUnaXaeNn2EDePtSPxF
VZmMp8AHqql04/w7JiQZ+NTzhVy4nLEgE3aLHJJ1c0QrvYOq0rwLX6OWDwzzd4DYRwZKxOUnLDoT
junFsaqeO2ee1K6bJYFEjfVlDBBT/96QI6uuwIW/JBfOjiqbz8t6uBgiuLNI5n9kS/IoFv1k4Hip
Wn4NiFbBzJP5VOS5EeaOTVSIQiYimVvhKxgdHXW7GnD+CT/lYxxSTngrZ7WT9+u95j9MWhcfdBO3
Ee8byln/QvbFHj+CSfOsSOUbKvhs8GwugfA5QxLFn8efp4/aO6GdtGjS5Uqs07La5WZ/Yojeqdtr
KdQxbN4yH1ZoAf7I/AlkIxUzoFvMEt+7MWTVSC1r9tbSZ3+e+yLut+bciJiNeC/ejI2CZOgnq5pS
0URix7A+WA1ln9Q+m0glD0LBuaGMuKfKXCUg4d0Y+mEJH9/rDqu2lptHjSz7Yi49MEwbC9N6Izxg
2bTF2TbtNzJzxv98cmekD/znOj9wyDf98Oct1Sgp4r2e5sjkD2lmawnumTUI8w/Ry75JKv8UJjUz
bSww8a7m1xB98Mr+s+Mo9o9suF4T7pbtaK6KB3gtyCHjxRhxt1kbnr0fWEYHDh5Rvn34wc1wmT3u
ScK2Sdcm8E0MFavWlbjq/kaFNiRDH5Nm7wVkIS+XB9TfHLI4Kd/iE05conwCJ/Z75t/NC62gNs0Y
nRuCUEzsTx57/qI2zBzHkMcoo5HjYY/nqhkMlNlOSgN4VgihR67YYCQmLGppy4QEsohocU4Hqv0E
204LKN8P8SSwXIOqljj/o8FOtiQmQvWTVGO3htZidLTo+leBsEzXQ7XMuYj/JZHdx3HMuB/hcZ4z
iYShZcclN9pK6AK4TLRxbweyM5F/7sFspRhs/WU+Qlr4FJwQQtsTyPphc+egzuRGyYJ8xl1uE8Xu
zIpG7NjPgRxhH27bYDT1vwSn9eAuqwyK2YKd+FcjlhD5DrLcNPTcQkGFKFWSYY3yEQavJZmPhd5r
rZBR+d64E4Ct9JClh7x+Z0y3agoJg4I2NBZUDVg+KKnarMxv1W4XG3C2xx9seG+ggNYLl++YZZg3
6W8/j7V+v9+YacsW39rkGIW10Ef9i1xcxlYxxBgFRQ/3au8tto573X7yv15RoVWLu+/ddiYsgMP8
Rz6SmcDNUZwHpkLosT4Ot9uira4Ftam9tIX5wOYv7WMiy1t/trozS/HMqby9lTA8P72wi4EPMNMt
bKqELzYg/ENQdnu7uS+JiSMfT3XbbPfkCAbz3aCgpPrTAewDfI06tCzyU9UpkfR/3H4188KuT9Tf
OF1dIh2peYqCxXQ8xARl3Jm7P5ato1GwWj901kn+zIx33B6co3MstRvZuxWiNwdODTmDJ6arkuqj
sMvTSUz3ld9M4lTXD7eDIrTeQyUdJfV9tNUSYG440sEUVtvv5SkU9ZbRhet9iIVGRE8EJ9qvZe7y
1gj8+q1QzH/ewKIUDSI8htibldEfgCvH72v25AWnjlfaNns7lDxsYiz33pygFlsil2QJUcbhxoNm
s0jSxbbu0kX6x/J8pcCA/G/4ABBE1tNtYbLZUrP+OLhGFd63SfF+qucVcMX1dc3kqMU1CwwjEQGV
GM9hwpKdviMPvlhgxw+e5mtl/kZke1yJ4E7p+16cc1Jt0ISzUdK69oGih+6/ZHyzu/in9DWkG/RZ
M8RyPIFvwcYYYee3gfxHzHKg+dTImIZCaHxvKpab5Fu/RhT7wU+sjNnyrFTCKYk3FMbkox27ACTK
o0KqUFD/3DN9ck+08g2oQ0kz5mdusYPqeo6aqZqU5TsRkIOXvE2oWS5kJag4pCGpsMLqYs682Z6a
/2HKb3VqrYzEBbZp5f1AP3u0ga6q8KB0KLykmrU0FVwTe28d+uXPqTQNumklUPEPwP5WtwFTZiqK
s78mHjWjKGYDhxNde3CQ4zInGk9Wp7csLNsRZohblp1ko9aVm3oPxw0mvgf6w/+YfZsrggYsNY12
eUl6xK6JE3a9Mgkc+U/9iY08cTGNlMQu+AT82zYFWMIaBhwX2YaTiJ9NK9BL40ZHvmwaPzGkwMNl
vp5G/efmZFZ1zfti2Xzi/RiCPtRl/1o7bnCaQlAzVHk+I3YE9VULVDzmHTrIRiZ+wwLp0j+0H4bY
8F00gbpoGua/+B9loVRdwKohgDmeeEQ9e3FZGfD8+rQZTpftsN3B8PtQFXp2f6tS+LPi4ypqWu6c
WEMN7VIS8QQaL6xWmvnB4SoGdXxkpjESJ8gA/h5ZfQWRDh8iOBn1VIhHVHmBDrQnhc8njOkTCXfV
+QzkMsbwai9Le6gPGnbq3CNszU0owaTS0qrPOn+M3vZW+V/o1gXwTc7TAHmv4kguno2A9yLb2N92
+DaTMzduCZ9oSKGhAg/gapF1gEUKcdmJMaPruec1Gm1iFZw0oK46axLVS/lt/KDyaGPNudJeei8+
ZnxUV49FGjV4qdo/YdOpatNEEBd/CyVRgvm1+KeGvGrBd0RjqVUyXZ1SWbcUI5VC77JiwEOMMcih
jlEBV7HJPgmLAXG4rT3SHhg2brK/8tFivUEvPl8e/S/xL661tG1cHQWaISonnAs2WS2VbtUkmqDb
95aATndT0mNzgtxx29sc1nV+2rBV+ZkMIk1ABi6GMy2EItnh7ovdGb6ZaZtocoBYvBqQfabtVs+1
ntsGbCn2rmE8qgS+95IOW8T09Ly3vBqG8kgjw/0iExDi7d/KQiN1WtdV/it5KIiY/dnzjmzzi719
YgFPE6iGza+ReQ5Mpf5qJdQsZ9g38H5lIoJ7DmxxTOU5XN/KJtCjztvAgHtOmx5KkesTkz/uyzWo
O5aieXweHRltqgtpqXaXt+YZCoLbeWohv4iEqdEbYsobaDwhiBhqVhoEfbId0m2PLEWfSZEYkUnz
z3kJalTpdbW7Q1LZ9zFD2t9w+LMSpWxu2roUr/rDl3k8MpTb8rWinIxA9neI/Y0d5oDh41FmoamW
6uAzWgQtMaF8hrqb6W8sgeg7JRRC0MKS/agxnagy9wEqXZZ9qQ207sytI7Me51RK1jIAmqPOur8J
LYnX0uh9RuTQHWApVEKWCm2yFpIoMrtiAS5ctHZZpQWkQD1sJjl1SEtVADgaXk1V+Y1jOKceOVN2
NPzutYOG3bhc66VYEbIOPOOY8VKbCiGpvsWf3NsXG6u9QWw3Zm5x0eSLXFkr2MlaPRMkIyx8ASJY
VZPYitCU1uat0Ha3unXsC4IjPBncBmVUI62F+gbnAz2CKeJKImgT1008uC641dUmIgDleyMMHrXj
s9xOr6WG8FE13fx8PWdP/eDkeShodz/KPwnSX/B9RlNErpDA3mFGP/wjDvLVX8pzp5Tu2SUidKvS
aSG3CKs9RvY+mOdMv192ioZHGpJnjtvkJ2oEC2XW+feBpjXILy6y7kj9yiCCK8gxpXpUBJeg3yTj
gqu6pMwaMehUY/6fJWg/XmSDRI2hyTE6NOKo9u7w2UosK1FrcAoZ7ETxjyoM8dF5cg8COeEBM/VU
xL9ZV6Lmkz9JL8fo1CR03UMlQ6oZZuK/AUkZH1x1XbO/tG4PkzII0iSmBcFsz0PBObUd/eBgK3EH
6lIj11HD4QiLbPONSy1VKJvnH21wA0VsMF6rETtpx+d1S+CPIVm/dFtFmZU2zK1J/MpL8inX0P4U
zLgiNdlSf2LbrP5GMOH2erXD4grlMnOawkMSk8h9VNM72/QjfYfrbzCnxSQPyaDYzUkJI/W2M04+
tCu8YoQ2OoY3Gf8FF13SW3G8dds93yx5UxPuR4yH9i+HhNy6zAbnZJevRWA7azg0G/LKsND9juwl
tWq7xvAbpf+iVtnoKdCTXOJIM/WHn1QIjUIMVzj07Dx8/9cvIncv1hXOm0G0JCCLzGDWqix2BYgc
/T2R11Cx42weIea5z/uLQ9PSYQEdDOVxZfcjXQUFLF7+XdjnfnGkzfxdwOlOuu72bvzcAlChLviy
HMYSyVvFPPfBZjrjv1HqDCevYrShR7DsKjw/owF9slTI9V+tEX1cMAD/7wby/GIpT9Xvgc7ITPUi
gri2W+VpViYyyn53N5QnUOYvltfryZ9/NXwRI9xqKgVYUDD/ELA2a88Jv+smRvcD78lk2v3Lj8LB
8aGYAV3IAtVX1SN5vZ4JZuHOeuZY+WGE4huvKjbcLqMXVVVEOIrDl+PEmGE1edmYoPD4hlH84p4h
fBJRxvTAcf6O1yY0HV7DRkZ+c6F7barVgtRsgxk+cXgrq8WyTEaIvn8MsAzEBfDcBQunSTi2e8zq
8KrafT8v3wgDKqt0DV7LrhpgU6Ic9KuSyzPinvxy5kFIroXbvMVRVculg2FiCW8RJBxKBnD+79Op
96G0a9H0d8YPvqaZRb3q0ZIPXluKgBVity1EQGHbJBUa9Zm3T1cZlyjLThTua7QcLUA5U5LeUFCD
ZplJPl1YmIx27XRWkbsS1aKPiJWOe1K+AFlEIooR1x6l0SYZpZVEyL39K2WzUTYCvtLZ5p52cryb
ewlyugQfZVbBtqRPgO5csbEUdmZZrPzjzl3q2scC3CQbpTQUXutGX9FmL7bZpUhjRAd7kCDXy/3R
lexPufzoB2VABMV30aYlP+doxMyorbX2rIjYhv/fKLhS7+86i3MKcbE66PhmD5AE51R3jfqZwdtM
5xLBAdyi1c8doN3IWpYrp5CG1C2j4ujystlNBX7iTzQzwhUyKQXThjwS6A0aI/PK/TFrJvlIcQMt
Z/a22A9IRboLP6nizezzv5Jbj0IwC8JbI63g/8Voxvg50Tq0rACejMfJUNk4gphWa1iD7U3ccTMH
ujLeRsaRAbSiO7ywwlSnqTsNu8gwjFAsjC9AJNx4+0GNoYyPginLegea85Sc3+5fPye8XZEF/xeg
q/cAdRlWrmXi/y3IMw11SgOYvXhL656rVcjL0sjvtiqkAhq3Ho1aH2gyapghOSEtmwcDBxQs/3CC
483+lxdQl0VDN7KdmKsRdRIL2BC43IHcC/15Gdiiil7uEanB8Et2i37du4KMTaUHSl2URXl8MEGl
D1IMLPapYqteauoYdfcPpX94xWT7p+Sam8MO/y7FrM2WboQCrOsGcqjzKqw/axYou3/JV5UNw9TA
B6SxjkFZUUfztUrjq9x3mbFSEF/yKSyIc0KifNbvVqwhgsyAuDJB168wvvqPktnwNCXRwnJ+kwus
THi1QR/Im3+ABAXMn6U+lcyAYCVPlZ8j9ImXfXszAGVPZdk35d01HYpsPFh0RajbANUhKKdCCZmq
rg0Uwf7eOAZVhZ3FR2+ydeCl3UEZNIYEi/pVEKrczvk+h2i0w7LlThwAJTEJfMfFN/KPReVyH8p/
kcFfaMtjJaBM5RF4Z/G5nxeTUCFa73R1YFMrIEurSjN8E9gBBzf1VDrXG33e4Op758gLQ2GTljH1
HeScOSOpuqYfdv2IYgsdN9F80KCnn3y5hIyCVBvxDRtY6sYfyWfWiWJjKaqWiP+0oOrWXgagslXo
zYzl4FO+iuHsR2d8obh2cvbaaRkv0RBFFeu35XolWLApgzjy4z3wViok06yOjoGam0/14X7bi46z
NI2R6f1wiiLb+nnthp1hskty5mSY2hp1kAXmYld2XRZzmsJhi3cvmP0JTc36JHkLjLyZMN4uZ/3g
WsNOauSBuxDDudi5kELm9FgoI2cIVCQWantqiXB/cassdQ5fEApLAIaZpyGjT7+qpjZMrTJzVALf
2HNcjpIWpr+FnP7jpx3oyThJmqmb3k8EXTj6/VqQvNzZWgKADtCy0OOhrub9ye4ecRkHh0kTMws6
ZBhDsa4oMvu94fWrI5bFHrkPlw13BHChI6xqOq/biWlBxu0jij32I9Nqrpb38BZfqzMJkro89rw+
W442Bq2YGcNgZ2oDbvDg3XjkgwhoV0XQAt9niYFKzErC48dN9Bdd1Ww0HrbJoe84casA0yjh0mAH
h4bF4dRX2VK6Gl9HuhwYIdNvo7SNMGUHtLRPUGZBAHdrIuK6HhY97h675MX3BsrPZWTT/B2lRjdS
LTLIW8bu8YMb85bz9p/vIxB2JuMWCA3A4bn/61cAc7Nzucfk7ca46hbzZAEMsF3+xkoh5X7TXV4t
ZECik1+1Thhf/cSnvuH/86DdM80zhICYv2UZNeTu1OwfOrgXVRAVNJB+qnjXFd8Y1b5/fLS1VQr7
D0+UNHymtaevl6ozTj30y1KxfiV8VOSwcb7NTrObQqr5/NcJuyR8Oql/tSneeRg39sIXeiuB3Oud
TplTw2KkHjy+q4RGrufHxTBuS5CJMPXS3it8i9BRwQZycAi5ORHcRZeOw+GT5AjQppGu8Y3cZLy4
OlQGo3gUrzY0+Qz1r3xGzvW+Ia4s5YrMZXyDg0vY1V5JdYgHY4WdsuDQMXvLMsr1Z3lM86e9E6wm
FiB1GiDT36oJScreizH0PoaCgiVoE/qXGmpeGyLGi9MqkbbEgkdRZbphsbgsKck7lSGGSfftnpdD
FC09e2iHr117aekIksIO0SNtZ03elNW8VWsqwglOgcO/Tq1SErhtOGUK2+lCWUuZErqnJ1Raqcjr
RH6x0tVTMygpLERyxP9CwcV4tCmTe+ONdBE3sEuqqcYewD2fRGlYQxROMxv9viNnhv2rMKFP999V
g1diQhBbHPzPL3BtUJk6Uu/GSzhf8zAg9KE8OIB8OKx/+Mr+F5zX7NoKacCd+dkXl3eJYawRFMgo
xsmTbaNDoPiykN/CMEahUuCchyodRw9MDjd0zDreGvXinBUQt3zwc4y6NOF2UZ1TBFa/NDnF6tj8
SzQHPAkLhwmqDaBeImihqRQE6FTuQN5jHiyLkcJfm9GyAhii9IGt+H32QIo+20pS9rh+p7XKnvhB
XzPe8nC8veHKTRGAKRRNaTajvXfUnYPRaAVkY5hSNqX6SECBG5tA18oXyNF343+srsehE85TXgWo
qadENjsD9n+cHoDsKMTTgMEFX5RXSrL9mFlTVq3amQmlTFWifZu7y2AKuzqEKIlR5icOkW5wXjg4
8A2zNT6LYtQPad9c4/skpfG4ydLZEKCTQ9VXaq7r+G/YHTi8cuE7SPyDnQAj6t8gReLVXvZJIiEq
ltJt90RZf9Vd7+PMPYcQ3PLYj1on5xSZAFr3jQ+wMSKl6dXjpmMnrS4ABb0GOqMmsF6ouAGAeutx
McBLuIntAX2/U9kMt32wytDFgMnXsjorUaOenDO3cFvz6nfZ/MWa50BTJUo4Gutrx052e1dUOs87
MxVIhK9jSImL0YQ/lvp1wfzwhqnGXNmHcSdl8xogoBvRFO1npxht9UeD58Ata+9/soYgS28Tzz+5
a7WmyhA70abG38RNqZxSwyKxxCEIMuBW/w/4JAfqDTSDW/AI7iuowAutenSqkOTKTv/bYujOCYep
SzvFM5tTHl+BpqwJAQsfDzyMGQbs7gwF5JoTMiNNN4GV1w7Mi1cykfgpJsC5vX7wYeHR9rF4dSY2
GBc5Kt3rLZQPTqS1e8JX5aMv54e7PgEQx32e59NgiTaygR3zkXrtnelAOOgCPyCZDFJX2FoGsKxf
ajehRz3oYAbnQgIFICMnVjQ0Ii+i92lNCvLR2yBYWtWdi6E9JbHqYgKOWVNOI9oG+STR8sot3xXH
2YXD8iSOindNEZuIR9Y4X3+FLPx1AvgHEKO74U3c8bNC/wvWxRaMbRLHvNgpcpPm3wIfHsCWuThv
huWPx0aPvyo+/tXtojfW69X/65iaN+uqaFarHsaKocxyNf8/SH0ttd+FWR1I2zNXPYzrFgdrnSsD
ESc42gyr2qeaDMFnHuCZYTHlLof+V1kc+vhVW+K75xvasWafuzjWVyicjJzs6AAH6KMBlfU8hTSp
H8Vc74owRHCs5P4cdGvL4ZEoCcLk0OcDfQolpUn0bV9OxVo02xNDGnY2HxM6eBuC5h+Z5ZoIhiFe
4tHs7JRfN13rgJYxVumwYhQyeQbE7RLqtOd+UlyPN2BVJtuiE3rbO6TRDnQBs3WVowInna6rZRtB
pPQoryDPzJvDRlpWTPa7IwZ6lyMguaCWKnHBhNP9wHMrzI42Rpe6sJgFZGVgyTV110jfwg3qnPQa
KKcP1dkEx3B9MtP0tSekralaEzZFzL9eDrkAQj1r4TXF+3DvZ6Mw0PX398fWqeAN0bwBdk3qC3MS
d2yODIXq9wvYQYluL1F89elj7/47AiPO/zU3YGr+3Yp1xyyVyIO+DbpQK0htZ6YcGZdApvQZHCOO
6JXE0atnZPsigdS3TfEysrM/yTkwUCrQknTz6G63pE5M+jcSqMHjMOsv5VsrDujFhoMeILdQJHwJ
2UOap1A703pPLOHtsk+iV28HCM83jYUfgCIoAF7hSQ6O9vssV8AAG/xZzDb3VvPQ8vuRoW57pS3C
MpDSspM8Clm3sGzlXUnibfS5MCst7o6jJBusDwOqVEXE0QDtSaz8mRAI71tesoTwjTPzw4euz8dq
bn509+sAk7ZkKjF1uKZ3SBCN1IoUsh+lE9pt+I9gOoCD0AU0uxQ2BjeHyYg8Uoh7x6yIhjRYG2Cd
WElnG2dar2pJ9ZFMc8ZKD10k5eCowLYviI6mExu7/XrGwfKqqTm6Uex3nqCQa19GBL86gnCQ+w+R
j1CEoHjTqwjUt3XJsMuJHFfF8EN7jszRVM250smEal5FK8EhJVFgT4SWnOg4m5LVHiUDSO8e6Ibz
K25LSwQTwnF8zwQgL1ZMt6ANVTw7sWry3GGx/MExnzuMt8S7xUIzjLFG+I/liU17ALTIOon+tEMc
lzq3U9t2pA1BKcDliWTW20aRGXex1eVCdv0HgziuAqpUmWN7Ar8XqHcD4RBiPzG2HMoSe/um3V0S
kzhk8TU+zFS5ujzx8kLWqobOdCMstOIam8KtKlVFCE57ptPRFYJI1P8KgNHwv0jNTMWUZJtWp9p3
UUIQ5GsSP99MA4hb4tPtwArt/a2z6D/ljZCkW0wKKJm1KPL1KvE6SQCFS5CLShHbWhCeH44GHtrV
9T5HuU50VTz4a9G6x7hh9hQ36R89I6iSn9kpJLDlD1i/T9RdOXe5vyP7gJMFE+POYo1fBptrR76H
W0XNYt6plsgd770jNWnVXmGs0ZqXNFOP+uaJvgKFLXkmNeDRmEVHI/ZHcWtVycSH7BaTV+mUSW/s
fWp8yi6wQ9rNwcObyma4x9RT1+fcRYL9/pcnfDNBen6UC64nUOHxw3WEe2vCFQvs4j0vnGNxBEmX
1ajHSmkh0ASzcMaIh+F6vXn9kf3cFT+seMREwDJYxekm2xCqjDCfm9CRPs6yyRc6SNkrbjMf5p9R
+ljPfr6QjIwJ9Rs0IMp9iyXBu7Qt1AzZrEUhI1jKxqKrEdRJQhcH2G+Q7zfLjfVNR/UP7RL5GNiA
kJnlMWnaXU4k++lDtQ+1Q/r+q9ZjbMY2zbk+saURtXFPXIgHB1loQeOVg09aA0ncp0PupToicUx2
/nwawes+8JfEmgswJEbHmXyHS8FVmlSgQc+sF1Fi/TUqoe9oCdH8FYHgkgSBU5dpKsvmLJI0Y1Om
5ijG3zd636X23bT0gtx3/EhIDygKD/I6Ei/pSPygaH3VUlEOjjRMwhKaLVftKAVWzp65ZVkpKO9O
qnixQcJcUmNkbFM/ELbKCRPdV32OMKDkzeQYAvTO5V3J4NIae2o8wT2F8/HREBUeRnDCcp2pxZjv
Nl9isJeFWzkLuMq3bJTiZVQulL/eVd7yWEeC0JNFOqe06fc5Cr6Rd+jbCQUn+0Z5hlpTK+bZ34Hl
HTMYNXfRBfjMmD3Qi8q3OXsw+G0IxLI5+MU3hpSPJjkC1EJ+iPwJDv1AYtkz+W2q2DDKmun6+1de
tUN9a80JoCr0h4aJrm2iKmlPf1XQTvMr3ZAiziNB+ahuq0AuVWdGpMWZMSROIVVWGdCgwQ2fsZK5
ZOoqN2DhCYOi/BQ4OkbdvGij8zLTSnL7/XYWQUGhBVfWxT6Rz6TAYl31D2Tcr7dAxXbCynCNFjb/
POnQTOV6oMSD3zbxx1WR3B/DIDRnqTEmQ8CgHE4ZqvPVwXHDEnkrnTMUlTaJFyg5RA+fIULVFZew
y5RzZq5TEVoylF5/zYsqIn4GupQvq423H9+vklYeDw2g0j+fpWgLVW0awiZnQr6m4Ny+ku/Kgs/o
QmJhy4XGYKBUEIYIhG86tORH31OQKptdcNLGqFu4qk6blOgoIp9g2J2C0pLx3F1g8V/KrqcJat+/
TJupyCyntn96xlZ5kqTwvcVwoTNS2qYW43suxf7osTTHJQLDOS+JunzD70/Ee8GdgIjUt1W9kpY9
nqf4q/GcLAq22qwbBRlesm1nGORwe2372gyIr+fZjd3l93yBpJYllxA8vz+UeanMb+X10wXlVxZy
eQu3qKwX1IVmLjPQH5zzzDq2dFudaebmq8oHC5utBQJVUkpofNYcXwM1+U1Y4ibj2ePwRv8RM83x
QKH4ebqOkAiYc26LsMZMgfPI+m0KeLugnHabCsRQZhvm9KEx9EVkP84RIbh3GbY1AYli7O1K41hV
Hn5LF4cv1F9Lyodp+8sqNX2Gus4wmkkE6A+Si+qmrU2Dr3cblYk8dh18+wIr4gF55tM9AN1X07el
NDqK8i6Cc3/bl+pBeyp6ZszTWnbuHdj9AA8wkd29g7UbqZ1IJS9DnYaMYRu8WcB0l1zcYTWkoPHG
5foSAeoumv9gw2uw8qOVfR0UPpaTjfWCI04NeYqDeYwxpot4EiCEgGoVaX3QhGcRxMIHWuBQguyx
hDtF+WzbSMTairUrnL+xIqJ4WiAYMsK6hdBu3yWXx5fRbR5eKdXZDSv1xQObbFVURNlcyUdWSFWE
tgH0lmIQOSFDaDmuxOrRowlEidQfaMxtdJGBqoGIgz/AsyJi3drye6yI0Tb4GLGgAB7GlCSc/0PG
TNLTAtZcRuVNxCA8Hrb2BUsBmVkHNW4w83bZ2ug3ehR7wUQN7x9aoTrmiseiZm1m3xtFa/pTrvDq
w/OP7sY9f+ducCJ0zedPDAR5usXG06LpmCZgU+GBYv0U/wSE/JC+UT5et+QvcYor/UInEoFg+MB4
P0ISkKLGMxxazd1ts4NEnH+KGNFFSbTXTJfVKi8v/qh/4/Y0IHDYMjsvCIAeGHkA7kRiRrIUCVgL
8BNkAhd+Tq3iiompTlTet1bnQYzwaIAM4Gx6+GCB9/p6TBLwTZi25SHlvbs21OmYpn6MB+EsvJ6p
GRYPPGMvqkezcXe3BF59EllxwSHkGZ6TH0/KEgEd3+bj43/LeplH9SHapj8mJnTUXDFP8zwS0ldl
CA4NOLNyTfHk9jTI2jN2FH+rIeYUaK+Q5faYN/ZHKgq96Nr+0wA5WuD7E3Zb2K7xlxC+zmiDN5gr
Edh6qc1NvuUe3dKFkSh6haYDs8rHR3MEgEtO/S/HCHf1da5zFKLxMpDbR8RMVLIpCuTPZTO7Cgii
y61crNwBQmnDl3UDGCstn/1RbbvOyJIwfy01W1TVnYClcPfHZcasZdvb7zEbCRXHcTcAGTNsScc4
NX0IzHCRTNPQ66H5bR3dLsYPIoAg7tetRiqgradSn+qqrAPBT1tbyh8edG52Wdl8NdJuSnFO6Zdw
tt2vJrH85prvRwkCShKVUXLpBBBDIazeQ75+AKQMlgFFx+NEfq7PZp4Z6vPS+6XrBtzLs2+shHC2
GkdY9p8m6TApOvprXzRXWVgnVYlgdtDAGJUBx77n3PkuonRLFlWy+G87xKT7X84SRYsJKj/7mMcw
eLvKE//9SiLA6gkirpnQ4yL2nDI0fUDspC9gY1zOmHHQxf//JyHL13w8fizI6ct3IViYPa6T9WMH
rm4QimE1opjef66exeKASKyLA21s9beBb5aRIv8SjXPcigj1jcjzZN3rr5bnE4cE+/QdhHLNi0iH
FU2cej7GkzWZqHQZK5ygay+cQOSPr2+sonMS2EazCPiZp4NepKDBLgMWe9e/KOTFW1xhIveXTX43
5iU7RlXrd8nbJEqUR9vO3IdiD8MGyLxrQ1sCCfhzcwLLgHAeQu8TOfzCcxKd1t+xlOAHXdbAqDm5
yxbvWfSEEWJN6C22dC8NtWpyCxooGTCQFcY8JlwfKt4UmecOOXS0XxmnY0Qtmr4F090mkwW/+Y3u
uS2bH0U+8IBlGOiFvf8yGFujXhBSd921R1qLeyBcAr6pgx5jsLULBClO5Jb3ZJx+IItoxn9bP+x5
PfFAEs/yyJ5ovxKlkTMjyKq0HSgKwXaGRSOAoafeD/CewNomfQbjNa0zscxaWVpVEPQatJaNKPZG
Db2dYL7tlA+Pz6dyzVV+xzdc/h+dIYrI3EazCE4gnOvkczJViZdcE41YSSrQ98eim53545zrU0Ff
buNwRkYGq2PEPT/93WsqD1XoQ6xOANCT4oU0oQvtstpl87GQbuxE6qBanfSZ2OqTCgkuZ8CH6YHn
WiV0tJEbxwh+f/W4x5mOoviVBXpP8DH6aBuX6nqDWv5qNCW/JuBLyOMQ5RXVY6aFPWLwcVm3obff
56/pXjjGF7zYfSdM6fgB9BIKVlwvdgw/5wgxE6iBolllAZbW/D8mUysZZT2lYJvdufyonDJeB7wJ
h957EunxY3bCCZKX2UZ1JlBtsB9dYUgiezrzV+JDQnkHnRPaEjAI/+RjGG7CP1jNS9mMvbDgPbcJ
aHzKm/kXC66tJK0Tf7vM7KaJE1ybRhafhvp9HKKFo266rMui9cTmhUC7QAz4UvIMjiZsuKt/kXrs
svdtXKV9Sf3bGV8T6Ac25vZB7zz0RVmAVd0dAbKF5/gXyVvDIp1YKxYEbSofjYw8P4qutqWAKaaU
x+vuNmsaiQmIBf9yZp6qWH2RIaewrRBnmcIRcBWYZ3bG4B2g5FWPrurZbAU5u+lYiTPqtadm2yCw
S62soiaUCA0nu4fbD4DpTbrqnd3tRGGykUZZrflqyTED3drNu5zBFFXCUmN3LGVhUpfP25ye8q8u
VMg9YlsG4jx8x0KNA6HF2G2AGlB35djwTPgOgDiaZ4/nE6J/1IVuAGVXUCZZsoBSHdEcDBeukiAN
9VfoEVSvsjemUIBsAfK0QoLT44/P2iU8uDImByVIqULVLQ5mmmdTk0uvy2ejOMjpfuS4FTQpU6At
MFui8MAz7WkG1JTw3fHK4r43H1xk5PTeJ04KEmgEbGy+KdNN8lhDhuIg8UiGQHncTrxOvFG3VgUp
hCfz7DmzjMtVt2Xze+XCrjYH2MbqS8fA824E5ol83dsA+RMuyAWkqbiZ1mE58uu67EEB0U4xY9jz
p2MrmZw9Bkd/mSRUMNTTobbeghnKMxOIMobK8Bs/dOurVtkixzbSfdSGt4cXcdz3PGkbktjBuDfQ
6FTKvgfV4p7phzfYhtQSAVRGFKPUtz2vMEsasoCIJ8A8ofpHeoq5TaRZSW9O6gvs5yRdC61/HNAu
phTrIl3Vy9NyJrOuitQREsms0rY7ygRVh9ZU8x18u68wE4UvSaT2a5Qz/Thk6RHFR4oKg85LrNzS
BPNlQTvCwzMJIVztYlC0452hDpL+PhlrgSFitgqu6UTlmvXUFt+ohYFTJt30pfdcg3BUdmfwtNxK
botUIf6iWpOpwjT/eJdrN4XBDarGUzn8kXY60SVxi94D+2zy9OwCQay8Nu7pRBfc4okULBUUwDLf
jHRN6BXZjxXx4hfBAms+szy2389LdHRxKi7dLDcq7jh94uCc0Uo4BVvC6BF9AHgkzVt8sRQinppe
xG7AjgiX8SN6aPZO/4puh6VX20rGMDAfdwbKeJALyWhodsgHxkubuGJBzWNJCWdZxibCEeJ1dX2+
Nok9OsaI9Or9c6aKY5XLqYl7V8kmzDxLstzYQA5dudzt6C3HMHtpiGjGahglFrbVBy5pAzlHjtyv
r+ZRTHmFjqqWEi5uJ0epxZaHIjPgP9crjP8WaIxzSwJtGkhxeaZLQm/49Z25B0e9PzoV8Fk/Qdt+
Vf/G6xmfzGLrHjrK8mkG4CCiiG7Vgv+/5XvhE6f3O9XRsk+7dQu8OWoFcQ1j2zBGejxeC2kN+51W
OzOEJXDZp7CyA65V/iU+6lMW9qm258toK2O1UKf+Te1kwLLAM39NWM3sR+Ft0ES4/NtbunXin1et
vqQyqvhROEUpnhpyfvbjyj6bJ7F441I9b6v0gAkJdVTAtV/bSRUh48p7idXt7bWOqdLb5EBAbjPi
fY36azR3YyMUcOnYrpiWmmczYA22b1VP+pN3x2YyWbj5G6RHrioEJfwhEW5Hz+c+SG6+7c34ZHGH
cKVr8mQDDvDWSfVGr/OAjDWshDRfxupiFNPM51m+qXaK9fVBRllcfdkp83R6/R6cmNhN7zIULioM
JU8wVRww1xGIqjXux0P0ntEoWKLnUy8HrtJviSsjXu53da56upuIkDNNChbcS/d1khkA2+PI52h8
hc1wfqQ3T5xsPuBzrj5jwBEOWGkpgI+6GZDw/Y1rrHBi/adtVCCrT6lhI4dYjugQjXU9UcVMocaa
iRDNci2J1AXjzUAHHdHAJy7ZWIsLW/2EdnOaF272877sXaR2BLys6QA6uEeK6NhEI6T8KzPxHBTM
Ix/UTlqBKcM1XC47SGIRYhUN2ty3qR8BGxB6B32NH4D/qu75kCPpVcJGe7GfmmE2PmYEus0ae0DQ
FTi1CGyzcz9cXaQkKDssXMUXVJlhj7XQRmKDwvPiZDwAOoLazyTLMXcn0Cbon5LqaEK7XX7J4gc9
K6z3CUEDbv2v0IZCvOIQpSlhPN7WObbqSD1nf09Y7ymmc3FiplZAw8u1VUzj6BPaRRXBicOj4VJo
qaSkUA5NQP7NodCJ7/Z6OJ91eGGiB0ESjId/jSO4dL+Q+MAwnMELem5ZKW6dVjn3JWtq4DZbAPLC
+DI3VaaX6mR/6wdmcGSkuJ4yq4UaZrIOczJYv7Z4oGsNznHlg8f52VnBsp7Iff+7cYYmprTAUyEc
oBzmEC3ulX5smbxpZh8eUui2x2X/j9st2ZhEZQteQIYuCiDETvDU/cESOcO9J21MpQRoasiMTZ0s
nfSzsZaU9sDXqnJEYpUdpH9TjHeXYROcnlaW5grL8pBzmeI4JgWfyyEnqfaU8KEJaHghuKbOF1v7
VWvGOc4kGctaZw1vkwwRBS4SQKFZxJ05BDMm1m36ERyeZDoB/VGzmzhfn0ctmni6mP5z2uhwi5kM
lmvLahz1vT8be0v7PTCq922C2B+BwoZ4zNrx1jvzk7zU0xZZpahnqPZejEBxMwnf8/zx0Ws35gQa
7mcwXNnLUAL6B+1DX/PFmljOaYM3ULMhkmSzDncdPl+BUvgo2AGElcFg7kqplZm6Pa0WF8NEeGSa
IKLJYm+zFnhDFg24Qg7ojXorN1NkaNAvOaot/w5bpvcDzB8jaldnZDFIZCu9mtWwzsz0Jd5D+U61
140hFOqxfDgjGJBrtJtSNZf4L7eStjwrehjcuSPPlYOiGAWrcDlK9I4fVHCIgPVj3Hzuj7P5N1es
XwbL8xCmmHRVqOxHanHrIy+deY6X6SHyNkYERGyNErDu1hNrSZhIxVz+4G42X4aBhW7/DcLsQlUy
IWgO2JUA9jTaSDcFj1S1zmyZ4L4U7Mzm1QNO+b7fITTiyWDLh8N3IWjEcRQjWM1lbMJ8FyFj25mp
02p5YTHEjhroganssgFseUKO44RXoFxq7C5Fc+o8XFwBrNy23+dBApWVs/1NlakYX39ehZAzBqvx
mF+v2gajt20MWQL73j4xQ/TNWkzFznwy+IISzJUumFHJ6itIlzL8Mnc3AMo+ooQzrgSbxGlm/fGj
XAT5MnVk4S3nQcSBYaBZbEZYdl7tgi6kU84Oeel8+anHYY92IKM7SFdSr06fnRWHuk9kemslTfig
DK2gym6RyBV4N3ESJ+VNdOJmm352wqxaZ5kJ03swlUU8MC3gwHrZFo43nuNzte97rUIwynul6Ezl
6qiINfdh9KB4uxru6YNJr/vnIp8UZ7/FabCn4k7B5qMn+jNgkvfGeLEU16VD2zP6iV6hUrR7Dyl5
RUhiRILHXqqn0w8OFkmdMa/BxhpPlBCzsiCAQo0HlVbYM/WtcpyZsOx9e1+k24NFcVukaBARfWVT
wqQiPMz1aeC1xZVTSjRcVAKkd8pJUVQfEkM0I8uMuXFFKAwuImTNp4wwHR2yaWM2wAbhiyxKqU/C
VPLDa7JMh/hHa0EoD2Gi2JYp7+lkODJ81Uwr6YtfTOZgp1oVaZWcVzcDuyPmCQ5BiaeUhkRPZyGV
9VhcW5c8jYCatApjb/cFO2SFyzxDw9dA/gn5WmTHPK3hRfn+zr6SYX+yu2wj8l7JnIEwgBLd64MZ
Z9bG39x5DCTORfeS5Otwfd6IxQa74XmOKaujhtZaWC38jmBvUYDiPwmuOcBxzLbtFSctpK+XwMvl
+vtgUIrNObunIMrSSKS1L3Ro8/X4vlblLpNu+/U4ndWA7+i79NgLnczOfCvU+Tod09n4pAox3q/E
w7I4l9AgGvtgzspKiHNCMDjBngQtOnpU5yWPgIdJZrfAuvSFQN0ezOaHV/5m3raazHqQq7U/SzXI
NjnPtXI0Fp1cpvSpt0oZg3XhfuoLQAG0zOzAGYRdiAmKj1myWwhWXejuZwcSaJkc+E7SeRTOlQAt
ggTCqjKD0BgLOpuIxmIJLWcyT3C+Q+8egg/Cv9UJtw3F9HmGn6HBVvh+N4NogSfNIKnEBHDOx8ad
CbAMf8xQgrsNqA625TVUvAsyf290OHn0AQbxzK4LcUCRHIEKicx1vjkcEWP26SxLDcARzuQbg2id
i7cod8BpEhomrJVXXpUrB+3FP5mz0WwUb9KL8QYgSWgJyJR+5cY58ogcPaZfiUIAChu+t0G5HfdH
Y/Wgl6121PTSd3i+9BUkREwcmXijPQMZKozPFrOXf/TiLVpoc5Ou5htSR6gfvQpJlAmIL8A4SOzr
zPnAG72TTqdDk6Gge7lRRrxPBkyZe5dj155yv5TIG6voZ2RqfKA+Uvnkwo+7oMdEZ8ec6Q3ERYE3
JYH8NGPXAymgA3Ggn5hLSLxNc8tRHKleoYG98g7aPgYXebxXbLJ36riwK5/CT6+PIXrCT5GgFxrP
5yKqI4qOb01Qb1H6/rd3xlFxo4KtgFFe4WJv4tvUyNApgGo1cg4QeYpTYrhph9URQK0DqaxnyZle
nD2fESMy+X0ejwW5BL4Z32spUb6bh88B4gW5C/IbUFKtXMSkfCcqd8D5b0JPNZJZKyjhKgH89rLk
Stgv8l6xdAL30SyrHcJN00BIN9AzQZ6kOqzuln/adabR/EriTf/RBm9QMM+lXyJmcfbM5aXlLRKl
Yk5yqxc9L2D/VQ8fCdl4zw5g7XQur+Zv4LCo5dJi6avjD0whDijH4x+CgJy1H+ulGI1NBwScWvi9
QZZdzhENHbLg2Bxq2OcF12JTAOH0UUZm19eD5swrLF8FIzBD1lU5eLV80tp5DkoSdhsrHnRprjq6
Fk4iOGrksDg1JDyriogpQmwdemJ29yBCynS41i41yN6iE+1w6QbQlTZBSbEJGp0Re1bCBu6ULLoF
IV6jZ00PMI89ZdSoQX9JidO0Gszd5+9+aS/hmr7Ct3WWxmPFpQQE1sRswwFpRzN0wBqpC0l+zyiX
besYidnis40Sx6nXp4lWkxeqvcFgGIcyJ/QZflpkrg5kHeHREf+vU4D7qKaqst4qedb/j8/q2zNv
GtfP8JrT3DrGHXPddtsCkIIZQpnwLQaCpXWo7Z/osXTVrvElNAa1i8LMfDHfKR/sEnQSjPwt0to5
6lDUoPevGR0Pu6O3XLAja6GzyEaNMYk8g/Ch1fl0HP+9a2Mlwk9XSgrncUqcvRHH25sbBHUwbNyy
wMJ9hKjytUuP3GS+8KoTUmzPb+ZQ74lcYcuXbSe+I5fmevTqcAhx2NaimwnoBOf+XlWH024I1f3t
QXM9ydQTQNFZS//Pl36p43JKofukFR0bUpaHsSr+KJ6wiu7Iwq9j6jHy7u0HTTFSMGKKq3RksMBY
HQYHQMQToUaHviN0yVIDvFrGJjIBvrN/UbrFQkIy7GmFv3KFX1QPUwqSxElHJmEC/1yi5Gob3Xuv
LbkwSlruCjseL01aw8geQs3YYH6fDPMVHNgwoOodfGNT0fcpkkH+Quyi+hSDmXzTzAIJ3ICsGZPu
ChF8hnMqLWju9+t8PviJZ9oG3i9polSj8P0u67R+o3no2jBpT2/LvKOkJByfNQExdkPmGdYw3tyd
RPHy8G25kJkQoKg+TPjBXh0NoLYGX0t1W9rXgMwn4fAOCIKSGTkMmgBWIZ7XHkETE/YrCrCZHoNI
nr0zdINK8cIXyaT6LKU1lNqUmZNFdlqTyDLVuuMtbyjBp2ID8z3OfCbcCLbeuDmywMA8A/p2l2iv
8ZuYFGvvHgHrLWXRNEWicO4MEr9hysb0OtPKVGs9C1g7qdjZmwiZG/p1rdEBLt8F9OS3w8alcr6D
28yP+E4P+L+HjByXtf0NJrupAqEauB/cfHHAlH6VrdTQANHEe4XEqpo/9EyWR0YnvyCt0/ZchGv6
fSGRhGWTYbN7H4IFYLNj62jORZ7oBxiQTafeKQU7lMXI899J17wQGIslVaYpikYNH0+NBvDM5th3
2OgCyKLSmVcEY78TV2/Bwo3Lu4g57CNtnt7q89wYUmtuGMa+TUltB1GlxZQQWO9d/yXhlJ/PANaO
hW0HwGuxD7Qo4LPaqOfTk+dVM+2mAdF687hvqkHqb2r2Ou61cNGh7zJG+3ZomXNisBjSYpgRdhnk
F7uG5tiPU24gSI4oc3cXAIU1EBaX/yBEpNKS2vW8788lV/xniv6u7U7r52MmZ42iC/eQ/JtqqONr
YHEtCvc1S4iXdhRcoSNDI6AXj2vovLE0RVUgK+BLhZlcbZLP+REI+iXDpTiPO8Fo+7CXjfatloBu
cEW8kSVuELh7lgMhiWMk+AW68aQaLVszLqt33czqADVj1Gsjep8uAWy6jf0lBw3qQcLVHEo5yq28
XbJdmiI980RzA62CZpITK5cUx+Wvm+L1IeBgAV8bqrZU5bp5NpLnnVzldeQRSqFS2QNINgfLqvzy
lv3qjDmTMLyv2dtBeU7bGREC5zbxi7X4T8xO2xoMNURGpf7NxkvjY6alYiggjpVwwF9nwqlTkVM7
ZACJQYUlJ0eacMurwK+/E1zna5js7PlrEx2ol8YCtnM7NVZAyZmnDHVsruLAoRYRGNxfODdco+lk
aZjz3tlPxJp8F1hFFi4jl6c9eyFOfEVsyuoIpgffcBAk9cPyiyfsHTz02LGmbQwuVXUAv6rk0ftB
Ue7TJCQtSie5yul1BD4KubTDTK8taCEG0L52JOrD3pYSmiU4mLjDL06dZ2PP8P4mRaqTAxfuPmbO
ik367N7i+EMz2ki/y+0zSN3yUmXNAF9Ct6ELYjaWcckSkIubK2mzBDGnQZQr1ck2Ccr0oX1VF0PV
whXGkoi+Hi/s0w6Ro4t/Ww3WHuOHdN4vaCNEbKf7b1tT7mHjKPmPiJE5xWh6dFTcmMj0xsywlPBb
IC1ubPBNB1NIAdXQfWMoEHZPe01Sqq49MO0naqhl4BdulN5rCvpOBjRQKEEu4aGR/XrVhz/4tYxg
Kt/6wSbUZU8aX3GgreUgcUNqIJStFBmWt0Nkp9IN+KijBbbeU537tZK/bmChhay2nQGz7R1tkPdn
1TOh3l0SSf0ioW13htBO9yplTOthGSYt9xiMWEbQHWlBhuR+30AfL5S6dpUSZhXVW9J0MYIDgZGx
fyLlHEmyu07NkaMijL0N4VQaJaX240XHnCZeHJ7evxrR0kW0GciJu6AztvPqFYMxFxmAlv5O45KT
ZkLXjkqy566xLXgF57Lpu3gGm5J62ZySlQwVIlHrxrskzyP2v7aCaFiSiE71GGz0BTlWjg3O+yeL
zJfy2NS7EqdZHXwTuIUANvapJQGvbUmkK8uHPq8//uQ8bfhRIhSbHeqhAXudf7UFdG7Jic8sdyvo
vWAF8dbCkFTCpqO0cgEowjsxsFTTSq3HRJLYtDPwEm+ztjwextWf5lpgfFTMQzQebSXlo/D+N02i
TSMoG+8NtvDBWi5awG2v9PX7jburYYo8oVNhjxJNwot/YI92vsGSErNRNhGi65tvxw2uJiwcQfy/
b2TbDjTWR5EHjTiqpsH42cb6ELXi/3l5oE/wqq5nOMeUQkXht3FbCuYxEIW4DFZd2RDNK+Db12SB
T5+UalTaNq5C4vOuUrmg720PgFyjLGVI0D9m1WdkTAGuFPVwuGgw5U9+pSIX7u2Wn1dIdXwAI8af
Umyr05GeYKQQRPknO4Kbhmwp4fm16SKsktdbf9wIY5NdNkXn2s8VOdtRQhPWxKTn1EEOLLwbQJDJ
JeaGxquuRaZEJIuMOanmqpvojrInJKC6TiJ0MnWyn7PKLlwt7lWSJK/i1Fz8ZCEu2csXzRJgRVWB
vM6z0ZZ8ROC0uV/mfzupDalf6D8fR72Xqo70ySm8AcroiwV6SlcHJyJV7tJ2bt6SaoePjOre6u9K
e3G6NO93RYNOhwOcZcuQKDqqJKNuPsZnjNylmjJH+XooI+6hth3xfuvoUYkM9xtvyvJQ9l+3SVas
GeX9XBdixteStIXWehrUMXnOl/pzCkf4a8fZ/fGhE9SYjU27s1QBPfT6ocOgLCB2Dn/GcFq42R/Y
k1CCoaiLD/RI1iu9YwfUV1dozADg+8kWehIv0orWM0xYvGf354opVz5kzbuaki8ckPVsQsqX4FuA
BeKQhH13UQawP+8U5qFHBvs5YgWUvPZmuiO5vTeeIMVVI8pEkXAGTDgSkl5Y2MEb5xLHN9gY7tyI
tgKL8Rs5OCwK4rZ+/WxmUp8ey/WdKFjQVj8Hf/djKrhsrmw7T48sGD4F8+qeoZlbVGakDHaXzg0s
yFVweexDzzFZwCcAvhKdJaVRxAH6W8Hs/jSW9cv7c4GiHcfd1LO8zg8ezZnewFkQbFIESknRl4JG
O+o91S6KUcrIafEuOtP+92suG2OL/SZXv3AV+2K1sZfTd6c/n48F09/9AXKBa4GLxRieAc0N/nfH
A5F94t9s452eDyTmxURR/iYBMjX/gZtcVhuolMvO6Hb2k4J7EvVFNeNi9zAVOqFmVpCx2q/lVA/a
+RQ6AZDjOEa3hEwUZQf6+elwPCRKPKrRn6tNPsWNKJL/EqOcNH8ITb0NHsMdQGTOHnPk3LyL4HUD
qGxF9p36cJTRBMZ2vtsL7CLQHNTNAX+6WBb6YYjh6PRUbaiDodi64NzHkNhmoYPy84Mh6UOC5wys
XHdBaU5Qy9NBkjELhLQhYjbidueGyn8yag8Xz9K7XSolUPOgO7mhfRh3gPwVP8BBHZHitA+38z/Q
tycZdVm8Bh1bHR+in6As1bLggkyPZ1SfCk8AE4vY47AeyPFNRosYrvkbL8baGZmEGStjZ59RO5MP
eGEYgjOnKtbAylQ9fMKqgzoBIaVqy1wwoQP8RbPC2zAYAHCge1mQ/cZMj2oDTTX/06gWcjIF/arX
vdm10Xat4L0otOu1HGjxKhK+mJQc/1OYsR/U1NIZmi0g5WgA96S4nQBsNfMV7DQadgjYqmGqQSS0
1uc5V9RMojHrybb1Lzd6dBOsSLu+8uXjWzVIGnXtGPmemQOV0DyTR5JURune4caIgzLMxIcQ8do4
qw0XzUEiYlgTdL03pebAvqrAJdRn++pLk8HU8d6+cCtJI67Yt+I8IINmbd55a6YYeGbYn0lk3xUn
uyJ1e0eAkfIbXP0zg4973Ky1cw6oH8ZBUNv0+EtJuG6OcQ6B32jAXQQE6aXWpjJ6HX8CBYpVe1ta
45wZ2YQcwWwp7RNb8ArD0SKBTtbm58ZyDFQUmqSoFWgxxWN8SyERy/2MSObB38nS0DI6MCZx5tyo
OZ1+AJFtgsT8DodNfmjYwiysQdd+N61PNI7dgZAGYYN1qM99b9Z/J0OyOyG/h9a8nf6/zp2BmkDi
RawbmQUZtKcQb/dvbawJCFwgLfZF5XdDq4Qxt+Ak3MZpxbD/rE3OwV5SuaJQFdSVr4BZ4bhTq4n0
JJYVxxIxSKUR+O1Oui0IVU/NmMqmVfLW+wliZKyQVVruEL8zHs1Z/yqPw5mwEIX8Iage4s+5frPl
b4tuoGyWNt26hpjuwP7yeoLBuFOxF7dUPux8GS/xIYlVAkqARPJC9Ks0vFJjTTmPeRTrMZ2Ait5p
28plM7lrNSuKI5g9SxzmiLuOpBYDdfKNTth1vP1EfOC9bFe2BxnjxoBJCx8ypyphxtTryI/RZPqp
ec5tIBvQYsPpWdlRBfSg84Piln7wxooGJP1RJrusN1I42I0d7qHLUR2qZaMkkwzfCy1vmEM+ENfZ
EwkqFBn4dXbLJ9dSRN42AXaCSzWZYVnOUSxqi/OcfgucsSvwC8Gn1SLYIBLksjmFybKTxc/ZnTo5
wakHWWqQzNr/d7On+e3i9StwdnVRWqupJMTjzFuHViDzAaq66rSAXSLq9BsTr8lxrfXbeNQrXWke
yrJdNWiD/NCSzMaiwqoLyAixSIGlOZtrCUXIe1GjphM5J/odqqp5StOyD3jUyOBgdeagQaUhrxx2
PYnbRVuWs76Gr3lTb/2ext3z7vqbaiN3trnZWabQWtv3PNVxFIwSyhKu5+8PK46kOaD/U3rB8lO+
ZAAxunZaah8F/lrq2dQsfWt6tawkL6rJA+vo8FoGqOUiPvSaYOr3aCekpf+dSCTlKm2AoL9nb1Z2
oVY+LkEV0G1cZMjo+p8iIYqzwtNZjTK/cONNQg+OYs/ZnbiHFtYMzpdLXTDx7sKUXB762MOPnqdg
d9ptXYB/hRodVvaO8hhmmxrE/Pm639G46PUOMxAR8qBAcDggrsFPVjeYBvtiHDkd/NqqKdotXIRr
SZwsymF7ZidCrPBVDMa3VAaVgoIhlvEeednkbpks8SKHiC5YYzKW/rlXpTe3Qjxg0CCgYkFfz8UY
S+gA3PKDGZyTDmkhgk9ndAcCzU0un085JUc0SdKOJoEPcK23GPkowkVLjyIjnB2Vo6d4REezltUe
6Dh+pzc+CljoTalV61NQBQnMDMl6GMm3jpTHGnZvffmG9QUDmwMh/AKjQmUY6vdX84g039p7+0Li
ahR4/wawm87b7DDLRm2Sm6xHquQwlZXePAMK+79ZBJL68kPgJf4j2Ks6cgrdpa/7wCit1CpFdMCV
L3IW7sUtVzZQP67DNG3ph6A/uEgKEfuunLxWfU2ja8mBie38i+N0MphGp/qNZKIKG18pS8zQ9HiM
AA9Ed4jvVc06O547JkKnMnak0cMWC+i+YRQrEjLS2SyFIGG9bX+nC5t5jo0MPQl//xqNRK6tRHa+
ZEpthEtndWEXzYz5t/MjLozhups/apddRKvfrm00Dd+hOMWQGtVB9ZVqijiRzdI0eyWKvPsZiYPX
Cj6+QpNiMMwZfTHb/DxlwnwVfdKMV+ElL6tJlYB+j2pf/vlYoESs/rdzDEzh2InaXAMYBCLlCR3p
Ju0SoMIMD6M2tkmJJcj69C4rIP0blfxy6VbOE5HkN/oJShWSBpO+c3pTDlIHn+rXlXGgObXeQu7A
BynIzwNJxfkA2/6CC/2BQqzQJpSrQIpuK53FBV0fbFbAKX3KqJYxiBdbkni3VlrGmeyWsKHbHjeB
TczKRJddc1Tuo6kdkgczM2uwjPd8a5zSIeUfHxVIv1gXlelUhkiXX/Ri8587txT9hWmKf9wzWBrG
vv1rdIysifiPKfFaT12A5ODbCAjo2rAd2Btit2Avhc12RCGy3DSH8yXKHlsXlRyfXG2ux6WeTXzb
AlD/1RlWAeS8bSrf/ls6apJc9hpXbBPaKEAZXuzg1esIxGDkaT8hAeIl5SEzTm1ibYEUVKmfUoRo
lISyKqFOHZLfc6/+z/fwSzTyfzReO1/3GqAHWVSVYW4x/Zsr4CQ8X2Cq4ZJCE5ApAYzc2QPtxuyu
Ov/XLggfpJX5Dq3rp1fs5w1UUpu822djFws2jM1cvGsc7FsWvj9UhI5Lsmj84+BK6ZIHS5bX7CjQ
FTBBPvncOh2qhZvsXiymJxr9WmaNbWY/GbmVrff4OKzQkTP+TtCyIIsY6m0jdtoElUQhzg+yj+nK
s36lqlYICqjgj2UR5vttQ/sUZxd1XEMFevDPEEGcaZwWds1c0CIL+IanFPKmML//MPDs8/keeWNz
L3lFO+Mndrp8a+r3MPxkXTPBRzwd0B0vXi7EqmMWsv9625IZ4WNcrBJlPw5iaflEPqw5nfwYYWqi
20n/GzZCk14IYzxbt2BVZjztVBcUY9bwwxUwjM5efVTEraaxfRhWIyy+TFtZ4S7CTwEkx/I548tj
kYflGqySrKHPGPoxIZoomF2+u7HtkZ6W5deLwwgEUh+o67tGRwkMjockhu1L1zcn4ZQVfHrXvw+W
7DkMKn0ztx91KqGA18W/nrzyuZoTtUVq9fDjrjdJo2M/tzKpk2UtJafW4qFU15AuLS0uD+D3LNap
0irrgAZHE27Z/8NXo+WwwxfMeqVsmkVx58mNkevsqnBmLNY50ac2BCbkN4v6sPqIPxzxcDeHi9I8
xpfEYTvvRfspR/6AAry2zaQvGq8mfJZcN9+Q0hYmQ3ngrRSttAPmPVfy9imckZFkqg/hNgyQTdRT
N1hZfDpJyxMTNr2lF9fnvHavqbSVdtPej96y3B8gzifK4ysK+0jSvk6mTx62+09dR5nLTkEOZFz/
T577M+Euhkh8FkJyF2ajMG49pPOn1PeOpp2J34Gh3+J371WvI6dE9eeUZ/zFz/AKArFSBA/DgFwp
lFpxT7YHoR2VwzAVAyd5Jz0dyOAGObVeWPHXZ1MzWHTIRXf2QkVMNENJ9LyAFvoZVDZxcg0n3qGj
c232+7U+CI3VKRqaLj+0HZcf6F1qW6T12fzKnc91ZJtETmadr5Q5tt1mtGlX0vuiidbBbkTXe5BB
o/Ggroy/7XiNoMyU8ZS5N2OinMFW7bSOl4vqnlEBgtdgMhEY7TnD+uSDBzXwW7GENqbye7dbPt6p
k7iB+CjIvQZEiq9jerI2S/cBy9KcWlWQSncfOKsy4zCytcVwUz3xFTacG+3Jj2dkPg7pu04RSQBC
7wqY8n3EqYQ/zautqN6vaKXnC/yjYXGh7PX4q/sVkI72DhcREmOZOO3e6SY0RC97SnG1O0IIdJ21
hOY/EUoCe+6VNy+vWT2l7E9l1DLDTFkPX2r7M6oaUxlnjbCOTnuG6bxCL+msVUSD8Yh5jp19fsly
1qIazIg2BRwL5ojAQdbo/zDEC8Dj4qJwkcC5XNgVYWCZu1FHzISr46cYh38wu2dH9cg5mG830+hh
m8S1PsbQHwCfWpN4ckRCQzXxUXaEdWptVYk6GihW2lPcfFXt3Cj9PwfFiKfwpTsJSxC/7GKXgHrf
oUWn4qKTiWbd6ykhM/kpralUUq8mgieXecZ3c6EqSoMqK/A+9d/aPZUiVeJAXAfqt8Cr7/u2uHVc
jqOLRgweIaCKwboRcLocxalAL4gD7JNwgURq06TtidJk8QQjynxqVyqG8srymyWdeTTfmJ6aQOdZ
bxLM4YsoetBanWSFK8+hmB+1KY9dQge3i2KNr5vZq51+K5KlklUZq2MpggO4sHgJHdB6Tr+7LhBb
S8MwafkLzKeo7VhSjOb2pDuoOtxw3pFPqsFD5XJ0BQ8sNOIDYpamplR9dhQWR/n7n1czmnnO+vdl
3TQLd+xNGPe6YB+LD9Y1JfFsTi//PCRFleI0NS7Z+b+b3C3uWCf7GmqbP2rSsPf5Z136hOPimKtE
hrLrxRkSF703GQpXfX172cBeDo/skul2DHqknP38dKM3NR+cjbYLfIbMArLfR38AmA7G1ZKyRr8N
wCsQxMyMF2XIFCytQZnkbT4IJ9FftsfiFi4RPovL9z7lv3MSEkrKnpyWhoLeurfHxc27h/0baqPF
KmHyaSwXDwW9C2jJSSbxkYTNsAIeD/3FlM6gJuQGOUI+XF8JBKRIgWBMn2Uoy6X47BMRr++H07WW
mStoF4/6UmvNW5TMj2vf8hfAmIc3uqH8GZ6vujm/bcrcjJf05B7EKTUpLlHZiCsPA6OXwMnHygla
XISrOMYKrNxnOti8fodHE8fnl4RtGk6ixQV3raV5kG7Tc7It3q93ghc7iUlZ+18/nu/l+eDRvXPN
Hqzy+kRiSKnhp/9S/yMnxtEwvHlva0tFcZUJgMxa8OeClW5CkheBCWQv2CB9HY+kHBZBdjh6OnJ1
P0t7FiPLtkfND29UpmfOVXf6GKrV8CW11N+56wvDPSQLo36eGmzVI6BbkutqPrvYGhbFxPuOAaHz
cmQEsJfEHijnxXy5OKSOkE1XI72oTU+G+Ykgvv35yZ3UPrWdSKLFOx8UHue1HW+avLtI2FqOrnzv
BmnwntOlnCADxy2Dx0vBM6ooAsaYKCjWIt1JbIXW2tJRjMH9ADt0Few0slz6k2+KGYlWOFbuFW6M
gIP4z4anmZTY+A7N2qreeXqVV0Pu12HajeTQPRFSvLBK5xCvtn7WN8fLAkUgaPxifxRnyJTVBS56
isynRhEiNONpRUCK8iC8K9cTSTSdqREmxFvbE3MGN0bsfqpVoBVSmUxr0k2FAj2PmA9iWmQyttEQ
qfc9FYyusD33X8D+ww2kM2mDaCPJhwtNLxArNaC4WOCU7irMVce1nvuDSxEWoPs2ZBcjV8RLANqr
msIOiAsRP8BDWzyMYDVioRRLjfestGBF8z183apwQx8vK3b0SIIyIXWMlNURXiTBkFWIA5clrKdp
1hlZhBzU4lQbo86an6hyeH0HAwXSRRPd6AnN0dGAS7Rdsf61tsNPJLVg8Ixv6GBeOyVtPLAgSMnw
/9JV/w9iXrsr21UdG/l6Lr9gP0m1CfA4rpKlBDUDFtpYt8vmLydeEe2w6FbEbJhDYR2Dg6+m58mP
3ONgmVqmgiRMpKXbKqqtOIhHLWhbO+p18UmJDTSvcN294Kb7H9JYT4xT9+NFRRMn2M+tby3NivRs
gdd71wceCLQew+gfb+xxmhNlkfHZBBTPUP1HzFDzLKC1SF257ebjhchFfKFI0zxi0wgKF6MyDLwz
FUchjknErLd3WeHvnsDbA2/KMeapcBZSLFX4wXuV7RIUFGS9DcN/3hQhXWRthOrrilViMlIx0Iaw
WsoZErMvnF2ZEiVvlkNzkDEXwtPlNZ2aN2Hbx6Cxut3aoMPjtFLJMyYMO8u9ONrZhHc0KRI1rw+s
mntW/CM5LwOiCONgCOpW26YLvJnk+bJpy7lEYyM2Ddcc5HP5yrhBe7QV1L1D+f2EQmUokarJ1vAl
MV+1pl3vOnqcJK99ZOReOz80PIgZ+QZrio6R9belzXFuLoZ6sInIvc16rYtGKWPQBRZcs3XQh7WP
xxdgyrNzEKNfaqo+E4AKIYmS6m/gdSq3wSoKImYshmDdu/J2c2lRKld1+whs4BxumCHAp+JOK2ff
RKGdRUZiQwtl8GToD6KU6oYBYEiEbZF4OKmO6pQ/HA3Y2y6Z+guD7g7s/VnfFYKIJXvIDl1jw+HH
VFXVQgorbR/bEVFrQvO1cXVXNeUdpLA7ODAw/BNUm626I3fY3fHBzGqAGDY9W81qpPm1q4c5Of+Y
5nsu8MY0S5h+Nr1hv3KVcpPNo9uWezb+RnVkYJgu2Vdq9A9BOFrxJ1MHgv+y8b+9bnmJEs0YcqYv
8zeQEvtNzLpY9Cl3Uhopx574+TAZJf+h6wXOLo8C7v16KLvM6KefYBHP4wr/q1d1w14VozAhI2BX
2MQA/G0n2BaEV0M+Sc89Zy/HvVxGXAbQNriGA2FMhHe0yVucxeKmGbscwcYK4pB1bqWR4U7L+Z6N
WrycpwhJm4CxuReEVpdbmTdVg2+JP+qvkEKcFktuHDrJ4v1I7+v6woDaeM/M9MwbdNgs+RDIpRnT
Lu7nF19B+tDhRAnrYP1CJkhVZJ29tzHmWtMH5EhtKIco+2c5ITvYuE9Eu9Vn2qUR6YZ9u9yO5ijz
nnwqGIo1Tdlk8xOJvecZ05f+skTjw9Ym82oGoFrP/z0VBop3rKSLRtH6NuL+4kxzVwy7BEnI3MMW
VWY3HPHqQo9mAH1Lron4TCxb75JgH3dLUVNwScNXFyABFTx95BWiLP3X8ISvLu2RA53ausB6QAPf
QKOHqvMA+WwrwqgbhOi0YCF5V8oNZFjZg5mASREUtfRBxk8AF94klTYQ945D4CE4Y25A7G8Z2t+F
wWwW2y7LgfK7USmIGFv+4PkvvhitgrLgcGdH46TkBnsvlRc4IJUwLK+ZeMolCC6Siq10xkTbVUIb
XQEPdXu+k1ROzr5FiO+F+wc2DHi7RxJbqjroGznC7SaRJqQ2A/6K7oVr1YQh4NzkUEIWoMVpQzw/
fjNCYjbVNVXXYVsy7eSBqDaaR1CAjb2lTOQWDMhv6L/wlJ0hSopIuuelnNloAbxJatsQAfieZV0Q
Ex+FzXc3XZ0M+m8dNPwENet3Z5w55ir2rflxux8piACAkUv4a1RXONWrB5agZYYUO62lPF2HXdDB
itV/GsVY1VlXTOJDAt5O9nl+/NSo/Bn6vUGIVfadg4ck3Qw6WVLt98k5RQLDIJds18tBcqU6vUxX
meRuIKRA/D/jLftdX4TtXHxbbTqIb24Ph3/wkGhv2WO0UaBnUr6NmMAbz+BhQxa43yokbI6FfmFn
uA9/6cUuoPhi8QxPov/0ksn2V/HOEmLqtqP5rI1dbkUYuwzzQII/rAKJCEk2hMoMwHUSbMPZ442N
m4jztkdmDSnJ+4DC6d3th3vyJ+Of6cJBtkv0eUoj+uIsI+EqVsIdP84Yr+rKrEglESbXTiWu5c8y
cSx2kCVduMoj3s53aT8bxmnJ4x/Vd0+JKCYvLoUKkoVYYME8C7ziwClhXkexQyjDTx2j/+w4hc+o
JKLh1cE9YU0UcYii7GbxIXKE4mZMHrlZvNytlv8yVmmafRkPyUCka+xi8JPkVriWaU+JMpIchRA+
wXgnFAnyfgrQxc2xquWxMp0yFmdk8GIku1K6HBhID9Vo1w784fXcYYt6j1B1e/cgZVnjql7kYHBQ
XESTFKWRN/5+oSWfOK6u4caH+uLx0URViexUdYKLr7PtQc/mq5CoCz7iE0OSxHvCUH9Z/kIbnSSH
3PFhfUuX/zcTHIXdkZ3pOSQQzttIVsklbsT1k+T6hRCe9iE9aFzWvPzAOIuSA46owQ8PsXQGO1p6
KVGyNRgogg/xht7PNjhkqC1rvgvMsYHCIRDOR6zpfOFBU6aFPmRM5aJunR5LzWXoPHaUlQ7C3kPN
SHpRELN0rnJoXalW5OeI79KjaKr9C0E6RMH2RmYlfKnSpNjHK/+6TtU4rUwrsVElonkoVqUDf9a+
hzZj2/vEuGy33FIrW2qn3uiC1ikCcHo7OHr/pdaI5o1rbkHmd3x8tfsPAOfTXZ1SuRtzqrkDD9Iy
LON4ELWyAnzwk80s1NN/eem+/adlZTErL5jYADVuFX6w8Q33hw37/kFAfmqvbwnLeeh0u/2Lh3+f
+23/dpRzwP24YqoSAK7JVYg7flEoO+huNIBLHqGc74Cb/cqU7bHafkPysBY0ctzOHKuhSotQYZ9g
gkScBl/kysXPD0oZe57KnzOHiU3QH7BL81oxek6BvoJOJPjGvuwQj+TVQDYKPzkDWNtyMbHs2a/X
MXFzVsCLup618roc/tOKxMDUm00/cmQxH5nIo2Lb4HKKIVE/Ui3Dk0+lMFvjK5RCFUZ7LMhn8PH5
MKmVs/XlwsrvMs34Fxfz273vejaNTILceNZZqfSZEXfOKHD1GDoZdvgxMtBlTY3flMw43QNO/VuL
zZTBvJaCFrMgf0XeFv/YIhNhJK/4hKBzFgz92v+cKbfGdD+QwgHxEuhKKRtNYVwJ8H6MGaIx56fT
8w38P/lRj+FKWHkyYTNx/8daMp1Oe6opBlo9ANJeS377PLs3z6vhi5Hp3neF+nvWIAAcdk0gUkU/
kMdKEkIjh9pdUYHeFE71Z/bZwnLldO3EBMewb5SQpNGYwzOZVfQ/HOkKp6tIZRC4uIyT5L6QiVfW
fZvWsJpf1Z8A83gyQjaupUjHlhYLJJrCnCjDRd8FiVtUYHI5zUT6SAQ+FMrthVEjZZ8C2b04pB/U
STGHASJQoQBIrFtpkcy8lRwGe1jW8Yjx8zcmV5OMhNgjMC62m77867RbL3fVC7FAWkCUV01xZSx8
JdEP1b+x1TNLolGqAEF/gLziM/OdEQDe6VdlhAgHV9xt+YB99ZHt120Wza85u3yRxpibUo622evw
zKS09xgbYpnOuAUm7+OtZikxGsf5BGbLHSMpwpUJNlIyPC2fV4+d9s3sh7GEEFLrXcn8LEevxuxt
YGPAGdCBvM38xl3bfUW4P7SPJ0p2QWCsGxqsmNhtR+ZqnD+xhNvZaf/p0Y0E7GvIGoa+90Fmy8yA
EhVfd1iVEMSqiFOn7RN+Xwnb38uRhS0n5gHuTvpkJbDiCZU786TkuSNgFd//3QWiPwSEj4qrbgyd
FpgWVVVhvpUQXtJeQw18pW2UYR/Th19FHFquqMHGTvjuuFhE50+mRXoSYP5xh0OBOPILo1vOeKpJ
Lj4SKYkwY+DCa3LsuZjmIoiyAVK3yYd83P4+FXCdSIaDUEZd3IsBdHNrWZXlfQv3ob3/IMR2LXJR
uO04wD/uY5L1zuNDoXGHZU8L1V8t3SKDFW8YbpeaJwrGAfwvUNk6qp/5M51wFgG8PZXxdBLqGk+G
ylIs28FQts1LylX/tAO/OPlL6qa9elaNElLWIGk2OvYm6g6KR2mzIQr71CPwX+Ur48Qz+nHB9N1x
W9bH87PZjLbeIiVtbcxsrh6WFqyTpoawswCcbqYpozfsL7LcVQNAEQGDkRm6D5KRzl2xEVoNFAO+
vkPQ5WR+E94edJ8FGCrkwyXX8ZUqBbQsMdXXuObX0Y1WgmWsY9Xcf6NGAtcL0I7v4QnLgU9Tn5hS
nmZUo6B1OBHvEdL/QgYbD/b8G8faWpjxx7EECIOHpII9xwv52U+2TcmC9FR7pdBLwHOSi5CMQp7I
ofhiV8N31+hVyzb0gjGjjAbgUyGbTqDbBZDByLILDc2CXv7utkHjp0QZb9t6+Re9GHeyZKGA1Rfh
/DuJhfwaSn6V0JFtErnCEah/AkoEroBwjmzlVnYS4as0ltRXtm934XQ3fO40OmyItl4NNQtjSaue
PEWblWSyW9VcRAMy+yRsp1KqD65JZ7vqyoKXoTDdBnvJJqdfmkpLRktZ41AzbD9rARCk2rMgWeoi
rMvap2KJ/0GLJwECkL5dAvx8czbILkOVdKNOfOYYxgYtBfh7gJk9Qib/i6DrB+5N6VXh7sKdyvln
lmN8Fhs8sMoCYqwq6C4hxhOskx41Fmx20Z6/BmQIrS11F1PtJZ2VLUBQT7sh0m7ikBHUtLLiNf2f
wSvc2Q7PDqyMRpcg5o3Y7o4R4Qq2/MpriHUxd51wRKF9IPpNoosUOOYaCit6ip8mKYPn9bvZDoXD
VaSFClVUuMiXZFt879emFtDCnsgFfAiVbxCQBixle6F0/3qc8SKcB+rN5+djeGXs761EzwF4Riaz
haBb19kF/e4f4+8MI9oWZJGqf9Lau+DEMFuLEaTg71zKEKF77rrHjxXQluZvBWyZTJJCDpTL0fLH
uyKigULj/lu0UnFGOcOFGkIKFLjP+rmKipSIceoFsx7woc37t0oDCrUtM8dghbbUgl9qRWUDucei
32NYsP0a9Nwz7nMq5cbtksgQaFMxqD/Lm14aYWiabcjJYlH+JmXnIqG5jVj5ubumC758OMWY5/Xk
lb9n7m1rHes4yZwQRKo8K7g9fNOoHqeyYuwu9PZut64MNYQj1zEdHInM1km+zUqeUavdlN8QsVyx
UlZUxQtphCBbooFyGNKcaQ00fLtHW4H2bfFDZFPFRtRoyOY7zFVbwYrTq1IvCS94v/fR8T8KEfAM
AnPDSVfVQfS/jxSxzdtzOnvBYXZlR4PmXJoFBRZM50+yUOXbvHqLWq+lEhEcoqDIebABDrC2/AN7
1oldIWgSmaTm1tK017/TEJhaCHxfZpu2cSEHeFmsVoIpSrURIfAOY9dBzCoPjjmwRe6z+y13h2G1
o+DvjiAC3t9oMFW6nFS0jL8nUme68fF30ocDD4P0sVJzbMWnkUrR85E8Yf55jBxWeENJvFT600QZ
wUb9z8zyUwd0iD8WSYZAYn8YUTgVwi+GAlG7Jo1jDEIA9bFsnaBMTO3yz4qWOpJsngov4abBYBV6
1vcf8wFjiytwkOiTVsCcNnGY9yvJjowBOb4h4UG0FcW0f3tQufPtFTt6hSvSu5uOeifLfb5/FuyQ
saynCPYWdNtN65nTHXBZJDGouk6KpxxpHo5xahcqdIbOJun3q06+MonH9lpf7AqIXfMcP34TjooA
WkUVbUEpXN17+sLipOa8qhujoOrhBGbM2E8RqVqnxyDkMii1q18WJrh4RIvmyDDiug4nkFSzJsbt
mTMLqH/UreOsIkL7HiCrZzCucdE8kN5OCiKIMgJ7Bz6EU8+baRH6y0FScx/KS/v6IY+Acv6pruf1
4X3DoUqd2ng+L9Fxo5QywKKTbTEtGZtjcQ7/5GU3JmYtqHOYDSEFV+ERlkfpdgk9QdAokx21Bj8I
aVrvHnRkmY6LHvKewf0lSaH5J/8c4gcHMd+0LPMfwvbQVkFvhPL26we/rr7/noqquQirYoD9ro41
8g0y2XZZF8U5vB5kNWFLwAJ0J6vEC77h0KTaJRSy8jA5dRTB0ov9z/QN+C1/OB4n2w4hYV7xSdX6
hrlnW71Y96gKuuB8IqkJ5ZJDxo2puHLRUI9KSObwigl1VgBGla+JKlmYSTTOv7vf/yFrhR7OmlBB
9ASKl9hy8XXZy7l49r2y8qPcXjujCDpdwIDcn01Yp/4caUqlXn1ciXhgqhcA0u07EsQpMKLcKRf5
a+iS85QaoDTuYQFkaxllpjVJ/ToKFaf5PM/8+zRfyCebIcJscIUnZPLF56YkMNvu3hl54U7OHAGP
2cSjkg+9dwLea3sF2qsUeNv0UXdJwhfRhxymioC1uehVvnWiCJ+z5KfuG6/TLTTIbA8Qxq2FkQZC
U9sqoPLb7APc+5x1x/Yccb3hi59IWk7z8oNBJQlIsNnEjZIR7msyybKxDYiQLLCb6w1tApAgEKYd
V4yCjWpeBizw1pCSuqCMRms2ohhn7J8X3DcyGUzMefcQGyIp77cc3n6bOXlE0FFPkSdi844RixeQ
n5YVpXG7e+eiAWGzyekz/a0IDYYqQAXy8UH/S8AubTMU1eXq0tIdQpKHVL+6edSPpQD74mNfKlTn
yugRRO7ef7TqAMKxp5ASWR5vby+A0BxxQwh/QWsdRJtKq7pQRkORS7E+EUElZHnfssz169T/bi7e
ubZfhQaOZ2BVMtoZQsWI8e8uO+LsVe3c7TVZKzpltdlmC07MQ+lr633EDLZ+StffiA13sCxleQ8W
O1GTMDOAA2xPXc0jPjemuKjzI+qudINoR42J6I8i+JK0RjcXtcff8tJ0+mBIJfns3F3S8D0ORF87
X+AUGguN4FTKgYOs9AsvbzG+GyDN+lhOVNE4XhvHr6379wB7ngjvW5O+AVoKIKDIIzF8QYxCaAmG
FhVWVjavl+W295cztxlrSgFrbtRz9RIFJYzILK65vy+h3TskbuzdykdFSpfHLyj2DQ5ErnCHoS7p
qxHbpBz3LH3ICmVs2ZI8zUwZ1sgWk23YuB+yA7Omz5cX0d46DjHJ7J7Q8WnCe5UrYCBKDdfcciKq
/Eflhb4c/Gr0CBtYJ7qQcRwgHH5qydaO61ePSAseQZwlLqaNQIixsaTGqDjueNrsIv9Oc/szhLw2
iRSDgRB3MGz+FdYcYMOJe9SbyU7lvdOqZOFV5RiiMv0hn2gQAuT6K1WLSSz4d7kf7geKrBhDyk41
avQuYyWFbIrihED9Fb9mUstdvlXCjyUx+X2z8XRejJ5S9RkzloUqAZzDScwaw7/FPp0dcaNcvcdE
6UfSPFsC/wYn8PXaQXew07fg3I4CAiEnZoJxPNIEchr4n/9/0gbkIyw0zwmw4DEEXBumV9f1iIBS
FKaiXIRmr//vQ3TD/8V/XIEyA3k3H5jvcuYAj+Of8RAgCEU2MroPXGUxLk7Htr6wIfJAXnhPTt7w
nLraNs4Kk56+YtIeWbvqxnJyilahiFxFVGBrrExv9dxm/ybI6seO81CBWOaT6NbpQsnLvkc1297m
v4ZLmtIIoD+4iS/nLIHUullFIEG8CEv7FZRh/hcVNZfhcAXHkIUf2qqTVyKcPmAtojUbN5irkpap
/moqGiOiC9n5QLpDQmXOM3ZaDlExMIehWS6kCReTFTcJjuHSJse3iIYIxcvLKld/atmv5ooUDYKp
O5J/V0qkIeca+EHnQLwZ+QU7NhVUGtdk4YUvfxg1j35Ril45Yl138HV9ZYso6q5GAOPsBgCWSO/I
itG3mHt18Bg2Mff+ESrdcn//pKtilT/Y9z1Xq+ap8YqUT0raZDLwZQMPcKrlJxG4/WGDMIsyTYYr
ePc1iy4ybbSIRZFMLk5gTkmnCH+bf5Y8YfNpzYCVNIDarAW4u/7l0CUxrxbigr/ZIs8jbKUVlccu
uOFkVXdY6DQnHua4ouCfQv73hnK0Dq/GsgVg0UEBcFO64mK5wcKYQjm7CdSrVvc4B389cclN/BJs
rD/HskwwMkUDbpQQDOkGsComALXl1s7YjBdXw/S7wVM/oatPrtU4U0zr71poWkuAI9y/BfVC9Ypl
UfVmqXK2Bz71TTFSlh2dFe90oyE30JOhVromI0c0sqKKDUqRYuitoEfgj4+H/IzQrqsi/Th7jdMH
WzBjCfOzjoi6iOnUYF5bgzZZCOLNrKEZMnAKkBKepglUPrEHODJWj45Rn/xPl3X7sQA8/NEVyHqc
Egn9VsB1tJFMhH5lbRJsknAqtS5qZJJGgHH3MQE7WFwpOS0c+R2IH1UizrbWTFT2Lh4F4cPalnHW
MeEgwIka7DoO3RCtCHip+M9sR9zFA3ubVfONXvoFa0w78hSAour9Wj4lZD/FD4lRhXHapy1it5So
emZuRuW8Zt7q0Xlpoca+OUgWWQYjKjG6707qYa2fAb2xH2BVN+mFGrNuRDWQe55fC4xWAo2AsBmJ
vDnIAbeWhzkAJINqf+D6Cf/R9LyxwFh6NC8Xj8H4+bv0eH8pqorJopPDmvW8rn7qzDD1ujJFEy46
hJXY7kTHx0UbWwtm/ZHQ7jM3YyEbwjNAEu2etLzTmch8qxnQx1l8kAYEvZvGzMIHxkMCLJ0NbC3v
HOcXUTLIEuwoOLWzuSps24xbY/5FuQoew+UAIAb8KopSZXCqjz/ZkTgHYvAzXxNz36fvS1n/I8aH
1GMoEythQI7p/CLkTYBGUVJAgBM4Ahrl+P8AGaIiTpZ8EPdcaxf9I1FCVe41FXl1q3tOn4BimDy6
pfU7AW2NHaep4CZG8KtdMaIjw5G7Z/eT7OJRCq4G8pBtOUEjwSM1sua2sEilmdBFLFaNwZZxnNO1
mpaLEX6YwvY1Vd8EN2IxZjDnOwQ7tWsZjnbm64z9vCCKe0T9QcrNbLqL+4BEboXMJWwGjHxbYIzg
PR6ft/QTQunVyKZBXxTXke2CzmRMOOTwjq10raW7v5zlmusKn++pKwRA3F1R0T/F930DQmP+5gIo
NYoVrxG7hTvp/5ny7TBeCGrYJU4ojdo34FOqucu9WCP2AoXqi+//KlL6KvYUDU4PVr+EQUZ9ZTIC
gbZNPe9ZUjT1wgc6XYRLcDI6LAFVabxg3SC6THiYXeSAwXBfN7s2MtsDGxdNtWfNZIx6fLA+Dxd0
noloNJC0PeK6Gb6fdyWIKOZNzlKoBn8z6AWG1fTDUxaLSN30iitszcEVuFwtROle4Mjppyw8EaEP
JjJPoej2ZfEVty6N7v3R+8T8flsVVriY8PtL1vi2ZUDbbvrswKkayutJsg4NnaxdBdIpPTmxdC0m
ImCyAYlAG5djgV0vUKDS9DIIWeTEleWPophRQfmKbK8XN+bYVGuBDako6W9jBshSb4V1Rxo5UMAr
oZzFbxx739eHbIGhd90MfYMoa4SalSDi3EE9VR/VgIRwnsjKnUXA/g4jVvGjYSCn++o2SzQJPPmP
ec8cS+0Ve417atWJg+BkBdkDm7BaUcbnf6VgS/yABiS69p4v53clv/qFNNUWR7WA2aLVXQNH5ZOk
2AOHEZLB1hfLgUUUG1EiesoSyCtpo6PlfiCZqNOeJPT8ppPI3GElZhVcU3i62aYFNJQdtbLm/BnN
oYImyMy8xBoXAS4dCmnXf6xLBC+MbpWdLMhcbliwNtjMfkBwpoxor5aXv/tzXpYvBt+e+QSzMR5m
KJ98S9ZvPXp+M7CODzu1Bkgu5lUew7XFPdJhWLIxh1UUr9zYjeqzKKTW6JqVLvpy86MJzTJocEuF
mUkO9g8MlDXtH7SGaSvGAjqu1/3HA0ZMUExblaXHDmNys0teON7BNWOQUuo+1xkGJXNfbKLswV/q
I8mf+IBSK9RauUMJyCnjusgsuX7tWQ0urJE+ELY5l4RjnQ6OhKh+AJ9MQDKPQczF3MPLAB0g6GHn
n721hDMy1GeSwxLOguVU/u5mwWAo9SMq4/CozWsgqidgXkKhU0Cz6VjEsxtwNKz3Yuehir3DqbTn
FEF5TdhAClwh7M9prwo2SAtAnkAAfavZIFqec9F3kVAee9NkUL9KFKLrh1ZQM/WJiugpJ3/eiRD0
St3+jwvmDkQsSc2dVIHtXY8xJ6JZd98GFU4lOG4LbCsEBOBfPbvfS6g4YiXi5BTm4sKCoVAZ1CX+
Aa/BJu3+VIV1sRs45aWwL505eS4NEBBb7T/R9Ll5VwbKglsoJDImsjhNHSFdnaBVrKaK4fI9OUJC
LppYEPbCRw1bCQnhDdD8GShjYRnLUmdzom3MEPA8TkHXxi8nJXl8vykIxdUPiRwYjLaVTe/TaCxg
RRJR2MVRaFFkP3W7o7SnDv4WrQLGX1ZSn0F7KMjAiSqrdIw4TsTfuaMR1E4nuM84NzrvdmaxJqbv
zYjc2nA8mbI72cONqTyE8zytawtrSbMTae8kWVtKiHluGkDWn2yBWgmQEoENeLSJ2AfO4aTLv9O7
O9/7gjYzYr7sqAfKyMY91sp/wQ1y8Ejkzw7gX6m6J/MsRLRY8bkpisC50v58tE9nRB1A32jAmBGG
sDoxTzXOQd99YKBl97Gnt473PAjRpPBY0l4AoBMvb29Ea2a/jLROR7UX4drUToh1m139FWYAiysx
OWxfYu7BzmRZrGBuXLIVqYUCAvvhyXB7q903HEZDZ0ydl3LN5rJx7JJqaoWgfXG2zMqHU535DuFS
3ren+PuvCVSNI1pqt7lK1pYJqp342ZEtqWOHXlLf3KR1gdLeLVIewgxSTAGmXPdKEjma8sWANnwj
8qU07F84kf0rFLKfTh7gzaLzTMiVCICclODV09lTjyLY4W6hAmrUawibKq8IA5NhLLAhXbJkos8a
VSIB6PaA4ik1xk8n4AOzLfXEMO63TBIKsTaP0WyvATHIyKzCHFhxmk0kVG9ke3LhccBTmopEFi+0
cY4cFqMXZ6HuE9DFMr5sqQfuY4dYewKnCN1hBbr2V2jKA1y0b71syVX1DCq31SXrHuA/i3MqtCiH
fqxe7T/BBY1dp3hD7/va/SyX2ks02jT/HnOo5pSzYtkg51dXCGxqm+ropZA8jmuM0EGSHD9HUVUa
WoQnmDeqaU/7EzQ6+ns1HUjzOChMadC9cAUUL7+775sMYFtwZkqanBwIJCWZDYV5ZQ6eK3ENb04L
leFLpAY9Q7Mnje60cnTSez1J142QaidyahEmWGwJtTvN4Ugup1lZ6WnTbAdq2im+ciqxq3i3OKz4
39P0JBEJUhpFsQ0Py419GnmiiiVwSwCY7e8ZOxQ1oLJZMQ3Y8qj1mpsQnUSwYnWAayYECg6UBXNz
tlWP45zIzbenAv+A43Q0iRePy0stQZPRk/Oy+ZDQ+ff1Eix/xsTUgctL2fr0dt44O0PTJLDLc8bA
khNnxMypu3aatMLC7vuiPkAA7GLQyLA3LUEa6yf8HF411mYNlUxMPqzRn6qGuZPdseGosp/0HmlL
tmB9g7lDzksufYIeHjLznu61IJZZZ4uqnT2McLkxwJYuSH8FX3nfn11Hg0SVrPt3qfUSP5PfN+QC
ZBoPPBQshNcw2/ucvXsAjfuHXUCDZ1BUBAvuVU4OifrIrZdJpWdLY1H7Ggwpi0ec+rdaMucSstbA
9/hHB1xx+VkvxtPGvLDZoBtMwUnzqvlyHFqMk+t7rYkXxRyAkzarR1K3yxphYZ56dQzech16+Sxm
Dn+TldS+hJ/Dcz605AaktYfMkcpmsQ68Mu/mTxDM5IgBEKrzmwbv9IKQPIYQWAO3zCON+UJ6U9IV
5bBK1kohNwrqjcDa+6I6nctVSWDJ+aekiiqZhwG1y/Iyhn/lNimA6054Ti3v7RfwJJwgUKHWE4XK
TmPjVNcsRNtQFm3J10UXTscC5wcryhT71vVL1w9dJGnP1drsTS1AymdLSoQjk9x2JL9vOMK435yP
2YGew1aG5Ouo7BIDiIkoV+YjC+Gad/a9m9i2MI6HzzlF9uFFV40XDv+4cyECMzqLeieKafUaXEhH
bTv2PdI+GUz1BZ4peuhG1pr4lMjtOy43c4NdIFSoAJJX86AJHhNSgNweoxeaUohsXwc4yuC1G1px
JYJKPwTrZMQjTV3+2sEC6cUrejwqhIPyhywv/5Jgd25Dkz5vXj+8NOUiqSoDN0zjl7DnlWMfP3P/
opoDHLJXCw/aPoCMIw3kyS/DTxjN+Pf8LvMAl9id4IGwlyROTNsGEuXc3MtXZ3oSLEUx8rJs/ycB
GWQb6aZe6gVC9I8CSjrjb+nRcKvGq2JtLqJzOQt3y/QBFCV/5QHONgYxGJ0CuqfNa9vkfIvcyEte
rYC2a8L1cgrdEVnPYRPV+JdbT+2UsKCQxe0/NzaEhBqxxyZmuWPZddmK+cXJHgY3CW4v3usyaOOb
c6M86U6gMc05Rfl76HUHAJhrlZXh/mMAgFqe69hTIJ6BPpVd2BLn0wakS7B2KPmmQcQfOMtQdVuA
aDDhh1MzhsCQgo6W/pUVI8ukaMe4X/66pOnLiw0f1oneutZ4bOoVE00cClJZhW7UQru8fC+JFOZ0
o/EX/myfCdpSjI+3mIA0T/alwtVqGSsPZ5BA4gsNSEUJp1PISe802idQ4360OCg5Fx66kZdhyVU/
3+Uv88IE61Eee6w1/o8+D8O8Q5jwmiMTxzWp0r9+qqueM/1B9d/XI9YAZryrNIiQ7jzcSD/QEA0D
OLDxIYxVlZ35IRNNKfceB1X1iN9NQ4WFvGmx4tgYwfRtyXH48aetFI2gVp6oRNleDPZI4Ce33SGX
NeqVpYmm2Jb0CH/vPrbHUz6eI3WT3tKkI5f9qxo68vt+J/zg7PnuCBl4YVat4hn30m1iIBbZyDFk
y1vtUYm/pwYRZZ7d1wCTsLWh7DIPXPr9YmNQRPOBPGZBVAHU3ZYZ5CEUbifagGBzI3EqVMJHD829
FW8FR74I+D0CWecYcRQx3JtWtuwYz2ktHi7tdCp8VBkGc1SzwpsIsQpVzx4D+4jpA2wqn+gACLvx
u+pYACsSgjFT20mJzbFHxL4sZR060tyKhRq4aVwrmu1B1HzQ9gmylthb6zU9prnBJIqEKkutb0rX
qcj1Hpu48aRt5t1IbCmDxJtn92he5RTP/2YMvzG69BkyNWhE30mHzk5GF+mjSrekNj+dL4lss3BR
k6mVj6xpdCgu7rubmur3crGp7MPr/Wm2GZqsbqqJL2+NF4umLI/kmJWZ9VdfeJYJe1SybX/MNCac
l2DAoZo4anIq8v6Crkw/Hd5C0HWdCCm0YFM+Uty+fDSmU4s2PzuFNMG+ezhoeXS965aaEYi1v56Z
JzT7Y5l5liLI1XTClvDGLxS7Zh+gEvmAUoRtiy7TVQQ7Tc+OlnNNreaCQCH6vI/CS7NaTlIRF9SH
PQyWX6oQCpj9FP82GvJ0HtSsgYutKux6kzpY8iPENIoRuoHMXsH5DAk11pCzonsCM8oH+kgqhGfe
DmPmpPJw9vcEgBwSLCw3MB9+X2fP0OtvwnD4g1kEjNO65x+oONWBKOsDJo+dnDeGNMPBnNVTN/Nx
AR2g/PW0xaE2+3VFDHFHjKcQvwooULd+C8AhlOJM9IGR+XQrj4NgtLhemnXD1Db4ZnW70zu7osCg
99lh9BWBmb+2ozZx3S3lW7yAssoqVmChNVuqfmkj1tO0ZihakkZztptOTQ9eVo/2OzrU9iqoqZvt
b8Md/0dQU8B9G0Fq/IdDABdKid1tGd1V+bo/WksUksYdFMGeWhTzeTef7A1UvKo9TtZBkva+dDVW
+z0Ad+nAFXe82OaDcaxkqdYDHD+zA3FkqTe4tbyKhiLjh9htWTgGvGdAe+s0kCL82cjJoFAfr+Or
JbHdFnZpfceqj4lR/a87yaDheyGh8e15e/OGqpvSP/qofwZrUYgwHDwAl/FGj/xFg2EGSUVzK9O2
+k+GscARSqVvWgWDpBmZIGStyI4IEIT499nJq9+WmiZDrNOunvn4Lt9GSrAGctl0ZKU+JIq7wAwR
9IjKObZ7pMJWsFVx/SuR6sCvmG9qK6FmY5X8Z/2EviEnZbcpgpDOf8ZE5hRkqy9UUj5T5IhV9/hZ
w1EcKGN7Alu16yI4sj4FIT4KeW+tq9kCGGc6CA6HTKAs3N8fJiE8Rn15kfF0ejArwcRdzEnnmIuQ
+ZbcRli+LCiPSzEFz0Y5r00sIw4lrgp76LflabCNR+sBopR6V2PJbcpRI8CvbZQccJhSsUDRqJPv
K7QiUpNgC4r8qptx09EwEdD3DtE19yccDURN0jU3J4pkItaWQDqIovmIoqod5fK3T7/l/vskvEPz
ipbDtaYKCOEtnKXbrEXMHrKw8hC0+oDheLMyDOOCD9zG0+TVkoSBFwgPkaH5P1kUkWlRa27d2JEF
a2Vd7uLEojzA17Vg+K956stARPu4TFlrAuMmw7tqmVPU/6AtVyJgmcdAkcSmG0i9MMElsx1dI5FY
VWYW48lJsp+CwNoh6ipUdHR52OSw5wGpAlqsq4NHfNxSuQD1D7dZw7CG/M2CJO6dO4CLJ9mNEfFV
8PLb6d4s+xfwwJ/yuy13/Fa4DK4l+U1dedB6YfirP3NUVq+iWxcstbJGq0nSZlyWr8w96aAbdCzo
sBorCXa6lqqxIF3uUSNVfSKNVsZTbnBbX+jy3J+tpZKeRmkIzLi9Q8IRKALIpnYoZcaaALNgLi9C
d7miJHi/6eP4yLQQzfr2Tll746CCxIg/XUw52JejhuJqzWnwWmH8Rpv6L+YaNMILFG5VeH2KjuDN
04Gv3yOpT4ZdgNtFGqUcaMwgUADQ4MIQfUDrk5B5IrpCvLoXady7W/UfgB6dpxZ1tyYZwuNVDS9o
iu72G+gxPPStBvt9BdSTye2+lBm79RTKsGVaovOyjAew6FOHzaYRWwxr6hLyNQieF3eGfSxKJHs/
x6gh5t/Bu5kZlKNtEpp/kX/Uu2NXJZBp1YPp37Be9aYVZnav+hPQyjccHCZk32XDUvFwmK7DMMnD
D1RXoB9KHJFMBo3yrbUrBCyTxORP7KNOm//55tt3Q2kYWytBFmSZnjAog5eYKoPxdhxgMIf0vwkR
t/AMK7D+qslEqOICfPwqihVqb5+qMuN94X5tbPIlS+Zy4CiKJ/cG0Yyg9ARZdj8i6JyQWE0p7U24
vAR08ODIpV26J99uLUBStj5/O0FEFIIPOFR4X6z73lChUdvcWbj+mwfLCJYZK+OV1ZsLd6IxZ/C8
B+ubfp400Eqn/92gqgt88KHzdfwcdgZFkRUank4jE2zb23fq6ds4+pbAkCin45yYVPGsiQPYWmOv
zv/e+FdjKjy14XuNCSSLh3ZEtKCiigF4DS8db0qLw8myaew7VieNEypSJI4rtyi8gqWaa1LN0YsY
rKEDR0J+snJ43tsT/61UD12XQZB9+39qYfIFMR/rx4M0xiQLhP3Ga/KmULGImIKcNHgO+7Ive9b6
bSNvhuSrnzeK5JXr/bjyjKTq+voEazAfVKQwpI5pUWFkyO/H6ljbB1j2H5LmZH32h2d+4SR45lNK
2lOXwQNipMMHmz+/qekrUtMseV8zjoSWKkUISyBLgkPr8w8I7Cixw/7npMPSEiXLmHH/qjindzVT
fYkQIPnXkClNP8tew1uv5miKY1J2hAdVuWRMEgLEW1kcEKrGCzTg1GQlDSFeI5DZUZBHO0lW6pij
h57dwJj6Aq5z2g3RkzeUbbMQhbo3JUb+DzEotHdWbk8JSpstp/dFqgi62VtCrclSc5PlONTfe9UR
9zZ3RxAgUIBapa9cH3HjmKzLPGaWjGNRE60618Vggf7sZH1v1Gc06gWZqRc9YFthujRvfe/bjQ9v
r94cYY2IYSMRX8+9NoWpRn4iL9QAoApEkBcjhJw/D+ZQXfouU2UOVRJ+ls6xl5rRrcFo5X3+D1b6
SslfnlisWypXK86Uh3oMtriN+unIAlEv6UBcBHJFniN4HsyUqu6JJI2gw72XJwvyiqxMXZlWDe2U
9WTnEUz89VPvFxurIIDHf22RfzCSvQzzcwG5dhEkbM/3GJPpti7GVBfQV7i9mneHoq1Vc0iq0yRl
F5Wv/aV/Jh8hJSmkJbr5K6JMgCq8FB0FCIjm9eoLrjHfM5NfDZSWtE5CQhgO1BzZTj1nnRPsaN+g
Z9KaK8PnZ8K0s7ZiZYBFDa+NYRTm+NqBBXef3QZZ7Ds2cP/jLck9sS2GJ/gfqdwz9Xq2kHGGLTdn
z3zAI8ScKHAnoRCObmyg0aA9KByv8VJtbHntcsqcqPqn9D5daUOeGT5PMz/CsD6pBQMxhT+Tx660
ikrUSEuFr3EhYi9Lqe9KnHbPgYZDHo0G/QJs3VvbBfKxMg2HtmObvVbJFiNpFbnWOhVkeVvcx4GC
VOr9nIYbpUw2TngEKrLjYxG7o/K+6H8fb/Kk9Xgn3dzOEGqy2xhsXBQGeWLtMASAngRmB2FJhKFO
s7H+e1DeDQoxIxbGuO1h0Xywd1j2DPugFSUhln7MxALxOsdj01t14PaK3zx1g7TtuUUCh4eyo4LP
yDZibfX2tET8pUA8afCAgqda8UdD6tLuy8FK9+qQnOwX99x4RZXJn4XvvKA/QAIU7u/UVIrjuE4m
j2aq+LapW605YRo8q5DEkG3Q3Iwc1ckdLKv03NdHHjDKP11irJCpv8Ur0eKguiyAlhCzW8IOY08Z
gRvQWOVcm5QJ43GawFSrxZCAQPKoOrALFPiQ8P9SH59g4bcudEkNvTUwP7QRsnaEgsohgg+Z/j6Q
rncEBPH8/hvq1+QZFjRfw/gQhS8e2GNaP/UtBYwsbvEfTpNj7e556zzdA2ecyJhDNCB183VxjWcp
9qnBFwL66yQ0EadkGhyuXjzWmXra5DiKyefGM60ytqa88TL3h9z22NUybEfrACUoOi2sQpTjS63N
VIRd4paPkk+2BbPz3tXIyWaJKOcYlnnv9Q/pmbqLi+lIOsvYyOZSUtMv4hoT11LxwmAxjeW5QFnd
s188vR9Duc8wzsjIvR04vSk6QwqGNoCNWcd7iSzj+EfjDvVKoxbiUljpI/3z76BZxzngc6Uex865
wX3lKJc245D4wuI4hxho+X7sN609XBeJG3wT2Jw59t7pEROIrP89RsW3SiFcG3B46sJP7LuaHRv2
6277CmTpfaDBO5ornvPSKDc5/cDXEuUPYvfHLyUuPQ/r/E6lnVOrvP61othVmePLCbJh6PFtm5NO
pho5GRnzxHbPxXoZKv9BwwJHZVt78SXIw8we7+gle4E+o2wTUegjMmCRnVGIKHyXkNz23GFXONPW
p2+F35basA7NTi0uRpmCOUIhz96c+i5MEhrEEJKyv78Iw3bBLzpTKRIchRktijG+/1LAz2NUif/s
0Qz1KUvB0relRatrl+09lYcFz+ANTajCbCtlRtoMH2MFP2Rqx4atwWaIDDspbjgc57L+lFH8Y5nj
RZI6EyoaH4zKvoHPl6LefriAIfSP6F0QpK8pPGpj/qfodjvqXV0w5iKh/HlQkYCxlW+cDDxm97OT
XXvB6BuEM9oT+MhV3tprBIcXGGsD4Os8kyAhi/lDYM6Ov0UW1JZBupTQsPxroG5Mf/HeFwyv89NT
Kw5WaoSmVfYXo+hNrkA1ZuAileAazFxMOBcQ+xIuwuheCLrJ52WrLOUXAiyifzqUUfbhhLbMhV3z
oLfiqMNBiKsB31Ik8pOjlhfAKHyMUem+ayrqfcBBwnA7Hc4dMk1Z6A9TE++RumFMt0HKUuWb0HM0
LRVM7gZIWFMgPRK9myUN+8QcvOs6IWRTXJhD8wljsGrU66gdReTQgURG8x1/gImB9FjPXagmmXuO
Cad65hxavWGFdGGS0WnwUE7TFs+Zm5cngW6J8JWFi2u7vpz3a948rUzn9aSnEq0deY3OT5mZQS3/
JVKlahJUZ/3jH9UJITZoIjCg74kGndPDOWlJiXyGtxb1Ax7+lEiI2xRK9uuXa1DP89cEiVomBxUU
53R0Q10G/OZ+dka2/Vdx0qH4Bfv5iUXEd4D0QvjX8DOQgBHuIFRJaEWZ1Q58pYLIgqrwEmPBrBvs
SN5sgvtPeYLWwjNxSxoRoaL6S46MmfrZ2xIMkhXOd1neGf7ETERFGLxCvfwx7ElAw6VxOZEIa9zy
kvQAV9bgUKDHStYA3apRITnOxRB3k0y8UOGRcFVefIryIl1BO+DthxWsXJKs5t3gZHH6URmmU0Nh
d1wOpBpdty55uOIgT/1KZp+s97454ODcusHeoGqWF1wRQFsfCOfJqG/Zxxwm7u8eWtnorKLQ/zeU
dPbH2/Wf/cFdL21S95jt+YHEpxG0dEL7fcMGUfYtINQ0UANgH+sGMEYOh6fNVxCoNbpH1iUata2z
6VZqlqfeJ8ySeXZYuUn74e85ctbtvVm/QUyTJ8Y2iSCVyicg7xXs56hzbXjbVE09N+K/uAj7jefo
FmMhUgOI7OedRjOuohC4HBLfj/AZ2vcxqZjgpgQm/H4/Iy7snDQLXAKMXxUvZ8PY/lT+yp9HcHuj
RW2Ouw7eVYAVKqHqz9tDq7b5NA+E3xnSNEfPUYXuv4XrTABpNTb6BqecnbWmIuNFpFWKzoIxRTRZ
HSjSFoWmCsUSvrg/E6j8gnooIRB84HBbN3YvOr59X0Y9FRLuma4tiCMcf8v2Ores7xFmMqg9Z+3l
I3/xHt1j04bXPNHlkigqJObDfNIlJ1+LM/0MSvj+6WVcDuW0rEMx9RfCI50Al7h2kEgAb6x9S+gs
CtWgi+l4nEq8c30SbOEFF2sSzI3G5zS8F8CYBg3u0Npm6bPm6vCUOHN4r3TFizH/tHBPQoLgeA1E
FSvnAv2wIf87sIO/YaB2iXj95ISBVIUSvzM66e19KYHYJ2jx1LbrA4e8qdeB5ICiHsnzuH/72qJa
kkBRQiAg6/uFT0BmdMhK6fZEf1Ktk3vZP+K+HGIaGxP1dZOksdpD55mVE2RwAbvGWm3SyykbKijQ
nmRIFQ/E4eADcukniZV9eDVeQVlewV/3T9jUEFhtvmMyYkTTZ+0p1Vw9makDEJmubzjlPfE0nMCu
13Y0xRYqIQxMQTOiFqiDr30o9a4p3Qo5YKxDUf7UB944+Ao+XpQzZojbLsJNuxTRpEmCJ91p1THN
Ubjx13GiBiC8J8hLI54TV9fqq63fpfKkVnLWrAgakZ3vK5pN5XyZJgYEVgXcCGfizdd9urlaQvE8
YKoKZaVHwVz7CAuKcD/kXGUIdoZUiiDV/6rB9haLilznEsWY/PkTgjAQHz1wxAwtqOnbKi7kIXZt
z/3QmF6lZW5EQt7f4Y2UwdZxgdL+5CIb7Sp0mc4ALQp8UTpeSnhZeRwQ6tjdvCBOtCBcAqhDS8XM
RV0Uy6kKOhyLd88NWvCdx8jqhMwrYqBgtH3qxCUye+0ZgrJf7t2+2dX3HOBVgSKrVsh0PQNtEcA5
4/Az0weBj84V0iOuJOO3MKte+2+cbEwo1zXmjcJ3ky7m3fMB7KH/dWGYqYaHeW2u5XVgUbdiu4TE
DIbpSfRm698hKpY3wDhPp73gC82aYZvupa54UxCvOYx1LtTzuBgZddQWXpt/BWFuKN0++x563jqD
PEp95bAteo2j/nmcWHO6caq7NxFWIp3hlyBPRv7+hxHAs2zeMzA80xHEGBksTFR44LsptYNwrBQ6
PhDD21/HYdUdG378o5HwUXdwvNuHRxyDZhCBlyXkrC9J+g0OPiP8PID85rAsW9xoZN2g+ZL1M7g7
smUwgnf4Y7b7vyU2dowKEiGv9ohyERA012QeEUh1F8fOWsByMOLD+zxl0R8B8IHGErwLG3HXYgUM
xTqKDUDrJ2BRTWL4rKcE7SiyT13y7Amh24bF1nE4BuaNMx0JBYtMox1L1jlVu13/upyV9Cm+EPNN
Cv2FOL96LTSD1OX4uJtgJEL8TM3DpKNRbnbEYHwrAqsUdFnCMQxT8hV8BGWeQlyEHEZ+j7V0Hh7m
hoiwuFCfW1LRBNE6ACh+pbcXjefI5+g0uyTJdNRePSWQcoDx8pB5fEAnP+DQdMQ9txiLHmkQ92ZA
fX4Ogv6fOpa/3bxEcbvHk+uY8Z7sTOHIkggxZ8XpmSqrmVFZqK6OYuphMimodbLSp41Doxzy/x1v
u+q0JBu+eiC6LTRtOOyP99+/ygdTM2ZH6rqasT3ExS7CS6UdmW4R/vFMNROgw4Fw1P4MCGCcOmdG
glVDJDfR3CY4Xeuu3I6Q1iumtmdwOh+SYhs90D6vLmSZAyNZYg1j7nYeJNqmkhS6qtCaT7zpIBfT
EfmEZxb+ONvBdF8OlrD9Z3zX0qmQE0VjZa5G4FHtpww6NWqOIkf6CVVJwX+cCX+hghvXS0535gBJ
ObpYNRdSXkDQIaxO1SmD2451E/YdMBXuzaOmerTQAFDPcNiLwypLUI1sEo22zcYd5DMOS2rJTqVD
Y63fcdGyGrQRO0FNAt6ylnUbViI+ZKeA3CQRQSHfStRVXwOJhEAW18P9CeLvZZU4bACJQskAVKt3
3iXaqXqwm+wSDXVQezOFRALaJd8AaefilwFR6x0wmwXlyy/3F+hlZaWPcJQy10msNyMhN0MEV9yH
oq4Y0Z1Gi6gASi/oLNN7cr1Op84eo6/sOTnixOk/dE/9Ca9+M45oYkCMkCAgoyPTd1ch3V/FASPq
DgybFDw1u4bP+SrLEPQqaU8welmgl3GtDwzuZs/dkFXkafIqfTaIuQu7tkwAjVLOvDMMVFwq1oan
r55aw1Wx4q5dfsrC34UFLGCsDPafrn6sBQza4dg5kaZPBQik2o7j5wJYXTDtMsFZGWep+JFzmk05
YcLIcy7CTXpoQpAYqNeEadzZuEbX+qswhZH34QAEgK/t3VUc1HZC6aFngJjEaeg2DWr3mmtctgNp
R8BQwpCnVQZV28LiX2vc3fGC+FgOAgt0la0OGVdFwvwUpm2XUptoe3r+Di/fVHBzo/RHcxVb2fth
Q/jC+Kq/DAqxqmXZl936uKON92J+7Pntxw9crLbfdnv5JPg4OEcqyceIhlrphjn3JdyxtKomwVg2
38/6xVQyYtdS4qbNGd+tDTdpGqSMrPjsobjEyEBn/uJKtchYUYGdi4p1tLUJQ5gUpLmsCLFeXc6q
L2R5CxnL+XfKBH5vM/a75/uarkouxSv65Qvo3R7RE1NJvIULsz8QDWEu8//ZhrnMHZToLH1ui1Iq
/Xly4cCWx/VQIxG2bsaKm82aMBdWdeNLcvqS9K15rDdQfCmyUV7Y1uJtytthybVWZfjpibD4dTbj
3Wsg25rsIBCFO/jtS+pQmd+W7x6uoUwYxzWPy8m5/bUGSg1z0HRwF3vPfGXW+ln5MbWt02byBOy+
uqtnmeslCN3BHrOWrAP1elwhpWMx5G3eVphfv5UrjlqKpyEHB6lJJWKsGSb1DvNcRp38UrSvjz1P
olIpMB5NM+rLdlJm5vAmZDn83cbznqRXMOftcxr1l4FfKE4pIX75Zk0cMH/ChA+LONIo/RiAFfdN
mIE7IDtqKvguT3Flc4UDOXG2+7tOew1IHdOySacAvHEWGTTknWx4pQcwHhjMPPbdU0k0dqsYsrzF
3VnmzjwvzlQm6eIojN0qP+utz5PE/q1m0bLhBpgCmr4/WV1u2a52uk0ioQFv1CCvNHNb1+jSsLCx
OOiB6FKGzPPx/VQPtWlK/aa+cWPsgiBjptQHEZTtSRC3fPtdtgYRRy7L2h6LRJNBt2jbTNc02wvq
z5++Ldfqi+MJGLNjHqwlQaW7GyrM3cAb+dy92fU9Z2kZhcnCe5yTSiC0OO2ZP1sRXdmbm/hch/UL
EkjrBq4jX28yNSF8DxUI0Cniz8s+LASKUJawtu0pFiK6lQ+PyYGEdvCaotLxM2CuJ2zmW+erj6Pz
0IqcdD9vWtnmIgQiGneD6TUZ57cL1+Gw7aGVJgJEn0jzUBiBFy8qTaHH5xPu7xaOHS1wzLjtkmVQ
0g0KzcSnQ0S/xkLpInUbd82JC1OfbcjOQEJKle133Qy/mEIFsnUPfjMjnc/oL8SohwgjOBVoiM1N
nxSBUrtK45njFIlmsRNHpEol730SZEXlxXzjTryAqILlNNtweisxJdMZE31QCqTPR86nk65Y/+Fh
aW9nTCayj9YS40ThDZwqWAZWYgIMw3xVK4wNjZs5w+r7c/EWxvGqQpnd2HJmgcfohyABkTtmwqJn
9TzBMaoOwyBJnCOiw0eZ6F6IVf3lsS5Vr03P19Dawt4vvAQBaOo4JmbjKEy+cCj2S5xwdms7gVke
vNmeYcEAl4IvNoK4E030C1XZyUdrCM+dfSw8+Q7IoZ1PFxZJCIVoFWrrqv16/buKU9uki98GvTBr
FHOoEO9lud4MMGe0Xlw3kDq1Y4E/XqrIDmcSmjQ2FaUN3e4Gpdz4AYgvShz8UUrtO3Ip0kYpIoDK
3y4eUF/sQVLWTIC1ukTNBBzJvoyPzkcPttbiNH2Gvg4oLdAsX/pLJErLoHsLBIZPM4eBGXJCAy+q
ebg3s6BLKxXYhHACuRwsqDECqjsJOjy8nErwMJC2FnbfbDUM+kxsxTB8uhqPhMJP0cRrlZpfXY41
SCecj8eAgl82Q/35TZ4UDhRWT0gs1sMH9qZ8OnHlV1tMKzHzV/qljcQbODFhtFSyZBuJMb0mzGHt
/OIrcruHzsLl6jpW/cPdPURIVRVoAuEH15HxUqo1zmahGYrfFaiFzhfl4F4FU6G/IhKnm+i9RvCb
aLo8/TYBW6b7WIAgGeamzG0mU0T8mQZVR9IX4Zs/URniRxyu2jd8Ahkh+esqCb08W8Bt+r/HAG07
qR2JXsrM4qzLaCKhxGuEp7hTSacxaFnI1MFYPB3n58C76r8n2IdhYzPQP5CcPszsNbXIGp7xuDP1
2uKS0DVsbpct5OIA0Glo2rc/QJWc0pRuiPzHz3OkFYaXjScxZDy7DDEaTeCNDpHvfVA8vCvAnsP7
/1jp942caqIoSAynOjHMogyr2gfQqHHFclhbafu9RGdrBe0ChAzIfjxKOqZ7RZfPsEV08jB+e6Yo
UsJwVjT5X3iDXNCObfJVly+CMCDlQIPQ/1cyqjtgC5EdB3oL3tAZprlcyqAlf5zLakobDxsyj5q2
36rLE4yor0lKZR99ZjEpYS//dR2/udd3K/dNxPP913rheijtkMloNiox4PSEKwskPRNwwHur0KI3
dot4ih1TwgWavnOZ/+Su3NNdoSMBbUhvIirmF+ydcKEqZKzH1GNKKkOD/NjMD5/Ws1a7FSPNV9dW
VChhMTSkdQK/hyhFuRx41Es0c1jHvRiXZRyhj+9CirmGswWRzn1jChfbyOa2XondD7Hxus3T7i+D
4FEu8W48Pz1EQbXawGyq0yUrCY3Ugf+xzZ3kuD3rL/PTMpY+Szx3rSUkTPgONOa3OcTtC7ldH9Cf
jS7m+FeDUYXTuDPUiPqysXRsrhjcz1MfcfnhSUfSh8u9DW+gTpDoTtR3AwaQaea+fhce95fIPoRp
XSGF96PzygOHk8NgwownGLp/HVtkMRDvtFb4VHz0mZClxh37nDfbaNh4QsuOz30PQlAzPmJzSW0y
XlaiFmVjohF2RRgeUNoBpr/glK3HSS5CNu8O15P/coUkfhkAuhDpm0e3zkq8kunVVDn78P2+1EjH
z2h3y8dI4r4eVOgneyiMaZTqmcFH5QQKx7bJZcq9gVrbtj78N5FqvBk0u7fS8oPheMwnlp+fbtUm
OcF5xzmRlTAZib+2s+Zvj25NQxjtA5FCWPOSUarT2pd2kLRKpPtmPtT4jq9HfZW9oFYIHq+3Pbe0
wZ1GNCeElK3BErnTEiYz87bRzmVk3PpsFjAArTb1IxshS4tdUcfCa4ykhKrKvD6jtxb96E826SOF
iFIEMr0HB5sxN+JoexjX3fbg0qR+YmCIsPDwhKicWkCEmiU97NoZDeSDzBWOqngrKhj7tqIBVuvM
z0jM9edkmUfOXZwgJV2LbE00Ngc1dSsvagkQHW64+sIF9ETOk09Ac7cBVGFDBwLPe+P/hixXwMZQ
hOVABSo83NCZ1MqIxwjkNFtRfzKDzWi9k6FCzneq4iAco6Y/SBQHJBBWQ7zYegB3XCeNlolcx3kL
Ee693JJNqOckjTJpbzvjhi86tf/aH/pMz2ONrnQJuQmB92OOJgXAJpbs7pejlmDcrf5ovsOMSEZP
0NUMyyyWDxQO8x+G2oAuhuGVj+uAM2/9o1qPet1eU+VbVQ/tFz5uisxkqnXNmRv22G038vK+Ezs0
XkXzYbCYlaCf4gEVHP8a+5Pgcyo5F4e6sl4H95dzZxPnF9FKAjrmMwiz36smdEwCx1XEfxvVT7Hw
VnQ/LmMpsoh2AZNR4OhdgsG5krWYB6Uxl031dzhIFw9dJd0QFEXQlmEN1dZI54LzvX/eWTRQmkl3
AuuS0MyutmaG4fO3CDZWYimsBv2bdVPqzy3PbHOybN/9Eti00Xpt2qe9LDWhPY0VxcOAC3DX63jm
RY0uNEuixuOtRcLV1v/6YV43TgMo8in4pB1nOKWEabgbz+gw+g8ouk2+eZzCyAnltHLEyXImNXH7
2FQS/nrYoUf1EqEzqikqqDHfr7uLqkZLcG6TTa9lejy2bZuBHnxD5XFNzd+3XgRF8wYBY4f0D2o2
xzknt1SS9zLEoW+yPuxXBXnlW3ZNKAAp98xv1ZyBbic14RMOIFJPOcVWTHqVp36zI62MI8mNS1rU
bIKBqkRSlg++6zxHWDRGh7HtNXhdiFp006NcsbJxm9+O7m6Ccs3vf/75MSNzQEshadhiTduNrt/L
9VBwnWa1UA5lK7spJ65EdPr0anaBv8va5+5OjfGlhQarljc3H/DgDj+rK414wuCqzTy1abocbWGw
R5UWBVA14IwodeWUw0uy6IqK64/SxXSxau7o42c36bxdbFahGIvg7dBF7IsViYglSAYgdn5Tb8DD
wsHj1KaykYMDFS/xoForXsmUvLOtRsy6K4myngKER/CNzmVvB4HvjIROPVHHT698xj2bGmbO7X5w
4dO47Ot1Me5r6PzppfD5TwvAedWCgqcTDPBf4myUTgrLZd1somjyaDJlIpUJvdVU86UeaN55disF
WBu72ERuEKtC03CFFu4H3QI8eH2YNOzdH98TJHp3g7hrooTdni4SD03XP06EpqGUOSz8FUd51/2I
NJVmqolSd7yxM9n6B09oqPd5TEdIDZMgvHlL1oU07Ucpl1DYKjc1UuFXjFW/XMUERsUOfJEDCEbu
P8sK2/evmx1mQsgoHsOVCTjYPXf56TaDVlVQUxkV2+WJX7f+Ybu2IA9GxG3ce8LmK46/d0ggwaDw
KEkdLSDYyig6e8P4ZiQ+ICzS5ZeRp2zzNCsfdnySqlURC1TlfEU3GOOrovUVbelE/7KTpnLLT+mD
WSWGpXWFbUts8QpgriSKJEWgrhT8InCxCWkJXEi24YdrfujhZDJQ0G7jubxSevXo80ryX2msPAf/
MnUtrD6zJ8iEBajQp2VN00PXbIUJ8T+RVQg0cltABPp4362M2rdHmw8liQOFeHJ2IPpuVhWkQIuz
t6TydZCygoQCMIkPUuueAvjXZ919w4Iye5AjuZ/LY9cpy4Gzk707zLrDb0i70vCwGZHHazRxeOxd
oFTlR/QARaXjCRER/CZtJ4688FJSsJMFTmWtMKIQUxMzgVg7zesYj41MbgbtP/uTFbcH0yErOraY
Scrxynlu5DjlA5sIssztHuXkJW4mY5+I1CrlYlXSE3vBWOmH1g675zswouOY34fVw7KfhibHZpIi
xCbm8eGApyj3BWnw8Z3ijy/74FJbPZEs700ejRFrd6TG3bjJsf20fVj/5a3CkB96zW5JMLercleQ
pezHk7dqu8uZoC0nTHuPoP1+V4EIqLf9iZT/tuXOvtlx26HHwfqKzjGxTdogeebOusacOR+pPubR
PqVI7JxPYgKg8g8dvdrjgWJtQEP2TbVd7xS+v+vcXjtwPnJ3iIiNNynOTXm0YK95rfujx6Qjcc2y
MZrqiKL+mJuzYE2GylgNg8SU/2Av63VhTZWsoPOvQSyzJlkWldhwCV0qnsEsg8NNRage2qYuIyJh
pX5gejUlonRHVGsT+bR+jQunj4uf9wYIJbjIxS1Y1gM7Uui7Mgo9MlAmAs8QfSGFMKbBvuGawCk8
MHjisRKWKsSSaZoG3bln2TSNeJqPWCMPq6B/a6lkgNUXJ5kKMyveX1lfriEA0qwsr2qhWUK4KvyM
hFqd+EaR/tkiGmzUVtn/cx6Sjgzz//b1T56ir+4/P6XMx2HWQk8Ry8IcGPgo1Rw3EooFI7MfpJky
wV6Ax5lb5aJe6NHiA9jpWeFX2Hl+2H2Kmw7nAexTxB9zgulJInoh5zo3SfNUUrNHZ0pNjK3B1ej8
IK30dHRN5tomBWIcDQuNt0jHsc0x0fLov8JcnQWsGNOnVvVQLTuwH1hq0fuTDXf4vi1AZOCgZlVe
MP6cA34nptTwdFOQFQ1z+AqgoeM1DmRTGpsQGhxIxfgBI0xVQWlOdDCK+D1uHepnSdWQrb9v139v
JByGSu/EspWLMtx8TMUcH8coMC9ALOCtHRv4wiPjl+xzFC/MsetoeB3oflMTJ6C6DujiFt/YONAT
+foGiAF9P46O9dN83tF05f66NzgVF2XJzoUfxljdpLJE+yP58O205XDRPNCL5Tdxo4+R08V2/D8I
f19ZIMpskPpw2jXfsNuJO1HDeNhYUM2p6MPDlwdj2Tw61lm2HiDOcNND2Yfp0zNli3dKdtKYDc8u
ke5KWnb1UFxEXcg8QsrWfa8n1fsvqwK21pbVohEZ9QPUYdIuVRsWy8POdSA/sWqhEPUFzVQ+UDLP
SQOdKvpvBX6AjHV/Z9WFg5A8l9Ez7WWxoOJ2TUtJZBOYm9xkdjne5rGWiT296faUm3G4V3YHsApO
iJ1f+uLcptET/Bsilp+yTV0kr7eFVz2Aqhl/X6tPTfmWuQreUt9rWCwLvm5+fdlhMX9ZHhUJdXoa
ZHQU+t1cwvPMp/c/srRfk4Cw2lZ9Sxe1z9BDFNH8aygY+RlTZuSvBdHUzk1yIxXxbN0c0oJmX8hG
yn660UTAOsdG0cwG4HVSDagDKHNL+lHU+PnyMJigpzPcDDtjvpzDH67zMN1HAzE9th8pGWZ3BtzU
loenMZLHpmC93v+J215f7gGGVkxwHq/XB7SRbW6ApNmL8gKONUx3M+IuTPd7nEA9DbutAZP+uIgr
sOD348bbt80YMfsNvYqIV4aQCo3uhUKtAnPX+QdalbLcPojTyZepqz60wXYDwplB0IXOy4R4KGN9
9o+7wByUBlEJHBMXt84q6Stpp2OnsGhMVG14l6ym+jnkbrvH0/JfjapjaXiRwY8MqMaZzh4+tfrL
qJEJ+UDIeKpfEqFfQgn9omPUWOks3icZcMbTGJ5EHu/aXKh4AN3ApFRwPAonzwEQz7brXbgz38Gt
P+GLncvOSSQQ5eVh/rXLpmqG3SVxi4JkSQwP2au8cPfWQtBVogEhyxPwnvZ3ibiq1oZ1abp+FAyL
wmX9mp068xwuPGYD7lzO0WA/MJetgoJkBFyoB93iqXoic2cmqQYESNlYWlANVEAxLXlRP+5gXMx/
jEBj6ogH2YCrU64i/6y+WqTH9/4x/BAEj5Q4HMCEs7445QwJKAs4RF0+VKo6AvVCT6LIffQc1l6v
OySTHsYbL7K8MSvSKT2fGd6nDhVkgCB8pHZaGnDzuGsDeQ5ZOmgUjkRMRcAz3Dg0DE+goVQRrdlQ
HHMMjfhnSo7LIz0EhOIXU3TBXpczdSVhhuiIlkFCpOS1+rOe6VQi2XBBkGHnQIRcUs3PEaahY980
ytyL43fu/DtS7vb3q8/aWbVgf/1XwjK1FaYRuRxb+k/7+Glf3lMoWqU3SPc0atgxTNu+MY/jX90i
UqqYaXF0CHN+g/tz5MHYWWofDFzaA7aXtPEp+M4m6uQbzLcZDKZPREOxQTltik8ccBt/Vg3wijmm
AZy27mdSRnM9Vq/lB1w6IrXqW0SH9MNz9plMf5EAeEnKxcPuUPg66SIwK3mHNcfh3kYTbvyCOdGZ
D+ROEA8xIe2YzQA/M45YtykZG4mXtm9pG3zlEELN/SYD1RxDS7X7vKQg3KVUNH3tdni6zhRIusbB
fqnEQnewqaAKE8kSdAzd273YX62YHgy+zZR6SNPmvRFG98+9l6pkQ8iKuEvbQVvzC4Kjy5skRCST
sZYe32ONEr9I2BRBUX51isD/rKM8xiQb75DfDKxABhC8LVVwYj9sL5jnrcFh2XI3V84yQh1eXCIs
KwKQokmQChNRsFCvC8kHnDsiIKATiKlVhrMJfg4CG1emCcC8Q26GXhmaY+IZtiXLlhMYxWmm+79z
oPT1fL4PTXs40CgQG2j09QW8QGfDbGJbbpMO2s7r2oYttNvVHClqIIalztlDoBJoQwLEcCcLYWCv
zRuke3k5jK2+XmBSy2vTE3GdINMZ4m5naBcGDw3oRflnMhXSq0EmpXAo+F6RMxuE1fZFfOE44MRD
ZYcOKvkvogkAGiIvm9Fd1CrVPhufDEiax8qUSLAxdJ9bbyepcFOVGaBNlQBsLB49q/iOpl53IT7n
xFvEp51nX3IHxGCmAxUNVNLC0WMwFwVPzVfAw41KMSz/Dj4it9xCDPI7ELGUwuoJLThufeXHJ9tz
Besd8RH9M1N8GlE/swWgXM1jsPVi6qfORe3LOw6AJh2PJpOUjCNguiXmwbaqLMILenDgszHgpIrH
mrG6zugDQ5Cafy1omlpUnTOwzHVBFONLtT8mgB6vB7WMJ/PcDlGp1Puk9dWdstKzsNFm9z1/mLK7
GZf1wfMPDAaJM8ceCw7WJBgfAWTZbIPymspuTucFwbsuSjR1seOWs6s/jYsZlCzr/UAG8XMQboLK
1Y+gb+L7r4kytHZ13VLQ29i+7ExehdlzXUMvBpyroK+30fnJJHt7cQJz1TA9H9t6Q5PKeTl+u756
coxvq63qqg3WagCOXoc4nZSSvjM9wlfADfP/ElHbc386FCYP6f+PgYtAtGYP4vOzeIxl045Pi7jP
whuJ4AbXd87TGup5qTqDfyo7Q3E7wb2cQ25X+jQe+2Ivjuzkda0GYYAiWPiQHmpk3ZGaHtkygdWK
crXVf2qXVFLcdqia3E7jL8N+6HdTTQrVrEnKB2bxn/cI88BB1zWQJBu2VYASnAsU1wk3fxLQDxc1
EZ3pRa+cS3rjDIP/3vrHhwh2sTUnuT6PZUwU5DkovqQMml8FpUPtXdrdIeF/lDtduNILUNWSta9T
zegFl4j83BnLROujn+wNm5qL5teOHLK5cifthj22FRfxsDHQofzG71D/dbTqpwcw5xN7s5A4D3Ee
H9URlCEYmYSydxZMofrPaJNiZRpkqwhZ7V+gbFvvsb4/A1ZKnxh9jsV+YrKlABTvlwok4IHHrPiT
/WM3SH896TSmGMyYd7xkp4ELwtnBjHJ3ECR39oITVkTL3f87/Mu1I0bs9WGaxXcSyrObltkPvpc7
6iHxwtJux55z84aOJRlcaPlYW/+ZHHSJGbIV71SgFCId/w1PAx5i4RtGrReNJaN6qciOoycuENCb
Y39n+eCoGl3oryNJY+jiCppCFwytqrqCi3vs5owqNK6kn84qCzcPj9GYgNypl7c7uSbZTHWhWX6n
1ZUaHtoSq2SmE3K72qkKD0luof3rf4bwq2ghfsIP1isxqb8psT5kAWOH/st/pb6afOWqJ9UpQYRj
9IZM1GB3I7bqgwSM6BLrtrWLXdgMgzu1E2pW4qKh2hGk27Fqe+FceYcVfHMP22szPPcegIU2287I
DG+mXFZVURABZT+9cNJP4qqnPSuVN8lyW+64UAR4Z3xgEGgE8aEi6gl0FRGLRubEqPKB8tt2pjc1
CKFeN1GcBQb9muno6NsbRhocl0PSYmchiAvguxf1LTdc8K7ouunwgyjZ1cy8ho4sv3VCEJtQEOVX
hZCy+IuA+Fvq36w6tBsgKc8DiXl9RRvhyXfn9TVPiGd/2mg2xb0T0pB1x/h5dhFM11MTo0e+W5jp
PHdc0H3vzqbcroifEBKFz6btDgT4jxGgQ7rVGvcNTbRV12WGRE6PWjbORARtSRkMtJCgGTjQYF9i
B7E1wj4fjEpM47t2BvfZ9K1p+/9SG5OpmzDkoSm3tX152FOvmbdoLFQjLDZHSP+FFIEKJ+JZ+ZQp
FxknEEnp64pa3DHQK9ID9lqSNeXL0s5JMPSwoMNCEsyekNPrm2bh8Ws/GK2hcvlrTtxk3NXa3FW1
IERVfnxrjC8tYsKprQ3atwJitcOUcJohUiFTKloGqgbYHK9v5FDZKzMmBU9KsW2QOxm37GMTornu
a7x1KuvpdseB9NKQekYjqnD/zDNWXhPyc0GViw68/E7mWMHyo3rpQ4j+b2CZQZEP3SzFx4gXum1d
nZaaW3RIZfwToPFxs30c53VA01NuG4xCxiegpD6fTCNmDrjUIekVqpWGQkU3LKDVa7OZ+9Gm9QbR
de2Njq13PNFIheDZwDcxmz1BAd7jzTFu+JEv1fTjUZJxLZuh4gKW6TcJ5q534GV2p5SX9/Irp/ym
LrVVl1pLNyL8TKV5qoT5XUXnjdczoOvgyEAqb68UAmsDAWgHh+IaqDV3LaDBnDlRRYBTueQR5JDj
Xi7NI+3uIEKruUUZ8MTckPU/ofwm9dDGgzz5HeW7+J5c5poadRP14CV3POx3fXONgZsBUy3quWWZ
BdtR6bWmVdW9khXswRPAVQcoOUYCOV5bs0pnLgKFyZnHrnKjHxNTaIdIsMHwfUsenMjl1SV57f9u
S7R6wW2Tr+8pdnr6mHH+i4wTZHMzNL9AjIJPb4y5SRy38yMk0q4+iunLx/mg71H96dRwkHmn9L94
VZL8ws+5ZuoaM4jF9VfRKafOBU4qfbqNPngJZ2XLSGan1lX4lIB6lE9NTpL6l7uR+2RxUVGYt6H5
Vjv9qmdQlPk57W7CoPMANN3EeGrgF78zxZhWaNez3LX31q6Sbe4dvO6Is7dKGUMMWKUx/m7sUvid
wPrRSyO4z4DrCR24WiT8Mgz2Z8tMFhHVpLvqyhzHR0619O0o7EOxofZxajzX3Iix2PWTW9aKqqxH
725vUh2+XmrYvAeIVEJXVWna5yOP2mhUGCLVsdCBzsqvhF/EZOEEzqc2XKggX/R6UEKws5SEk2jz
GTSgA/6M7vVoQBKNpz8KvH2z867g5mt1jriBzd5aOEgS/djfQpQKByIBhVQgWymRofQLgFUKnqzD
7hmiwPdL5o9EX/iLDIaBUhjIaYKVb0xSnl/Ks8DLCdNtoRSANcnMmDtAkfgNnSfF2eSpQWtTK2L6
KDv5SOlDd1SsqV3fp+dt82zZKElDYezaMQ0hTeBXByq4YoH1HidX7wHd898nQsaJ1eqtI83wMC8t
il7JXLD4nX+QXcAuVHaGE5WdZJdogjIBuvf9avfd2YXFmWO7ezNL1pqtbNlIt9RrO6HoZaJi/0hV
tSrnZDk+Chyge2BE9LW1lIm5BjAJUsyXN1KbifXJ/8aXnQ2uNog4vaErKjZcW20sw+WFVFETBQ69
dNNCKMo6OTKoBQ5CtXpXepv+el1eD57WENBSfXLg/TG5ysaLAXzntzZfFx1EgkC56dYN3D38Nj99
x3PlvazfSy0ZJxJronAf1xVM9hsehigPqe+YRCnRyIBk0icxURV8mSDIBgyHq+iYuxGBBrwnGoKW
AD3m2Hynh0II8dJKuBmqOVOVePBiiVTUYUUy1BGKUImxf2bJrKP4gWxrYsMSTF8dzyZ3t0u/xzex
Yq9o4gE7al/2wcwsJTSFY2ptpXGvEUJUVQk7ls88BBOJcEKtmtEB7vxYsZozplBlim8qroaUtOsh
Ad0GS6KM1HZ5QbDRjLbvgbvldzLe94a7cVp8NDidnzlW+YIXMHSEdB25dWeklExO/vILqawUGjZr
q+XlsaO4tR4cyoBs502APc0SO14aGgWr3FUWFk7IJB7WTtNJyEZygwUTXl7SPNMdMUIvVFqkJwoZ
K25G+CBwKbp9ngR7U98rQAklWxQa6FIaLZH20i1itPFdbAhONw1Dt4j2p2KVnV1yGz4ACyB6eD1T
EXfH9PDXiKMiz65JaTiiUv/npHiPZyWghsDyin51UYBWy18iBD8CB/0rORFvP3JojbXatdpzmRHv
IugUrYuqrM8j+0KV2I9aovI5+ONNm2qioEmOpk8BZIyzYeqxGxNo8j9QTir05//ZWjGWbpvR0Ipe
mpihpScdFYkcSUQ+D0HrOuRillxu/S3xJxrR9Lw+WEnOZs2OExLnU5YfluXGdRJXuniRPY/byubi
kHXWGLirp9O23LZpQ9M/FPMQiPLA4CyYcHUCivG/ZWXXXRWAljC3OLFIp3I7zcMYjO/yqy4aJ2T2
rD0GPnvqwJc2ut0hhmXAf0b4KPJioCRb9n1Ppb1GpdobmbbgzBTCAQ5W1t8FvuLB8MT1qf2GVk9D
uA+UC7fxUdE61I4Tj0hB94sThbbMWTHnNJoWrMxxGqRxEFNiZu0gOs3f9o+qok2yrDoOk2EwZ0ty
Ax97AUUa3KFT2dQ46+lhrTNKu2FriueMkCgQMtx5DF64aRoJNUSgAonGLwZ3T12Ev7Voe4R78JA/
ZyX8+RAhbDQd4rT4cy2YLqsb9tRAx8Ro4f0ruEy7v2wy7XGCNUN3FeM4CxlGLcEOzbQ0uglZ3zrL
0TVHXkn1u+B22jkEyzMCJiYEANhXeq6srvXLV6l/Atuhu9FVZ9YAipmj+GC77KJG4ZY38fKr8KmC
2aC+FPkLUOrBKPiWEDZe1+Cwy4idglFF0Es0hL6kIBlKfxRztpyRo16DE+Og/G2t8YZxvRunSyFI
5X0/HRzqfVt41kRE0WfYMrk35Xs20fS62/wsEr8eyCXaw0wNq+o7Q1ZKnxjfdp1tyaM3HW1YcdTm
1QhtWzquH/gOYkMxCLVlocSj1azSlHFCmMkIZvA4Xq455Mwz+H20IAEvcSbWOH9r2WAo8RFqVMgJ
y7Zf1gnuEYUf3fgYiCaBuFQVmMAYrx+yi4RQAxEyOv7nw48DgFVAoR/nQEmQn1GZQdPdvbfzfJ0R
zC/4lixCCkUDlD0gOPzypuTGJG2XGRCxnzG9SwFDQQvWd90Zikud63t6gystruxIX32O5z1UCE20
sD4RsB3/LCIWJGjDJMPRH1v9+75ygsga7nmg1AnvIMkSwVj0pmV+xr+N/qMLc6g/XBZessvQbxXd
oNssqO0CErLdDDQXa4RlhLGJY2CTU2pjWY4WuxOEHBtjJUbPWnkeDAlQY9s6gxNely5LLsj1Cdt7
mt4rtDMGSF3r/x9YjILpHU51hwFS+bEXogly9abUYqwGjpekeBRAvcsLV83TMTfATcTBJYiHNfFB
zrErHvQa7IZDMof8hroyOyMu7u3n9j6jCXbot2FAg83PO25CmCXYyJA1OCMmf7Ir8M/ZCQ2JpIsh
/ycPaixVf53bTFkmJTOTchA+1pxB52g8UKDzMMu4tcI37fuHM72uoFMUH/WVYnAfJsMU4ys4V4+j
N5OKMn4KN88iBSLo//wpXgYlB1UgsZBTRpbW7XA/i9N0dt+MWvpYdupq3f+oOuCtiKF4DgBDrh/k
C4Ny9Hd9b1UxmtVtuEVP3ICgoWdzMW0j4p3BWHYWCGw0jRw1LOekp6tTy2GG16roV1SzDdPt9rZV
s/E4rLMjF0FMldAVku5fGdataf0SuzMgMZw+xShrUajbVaJstbP5ALE2O4Mibj1bucbTAX5XA94t
zvIhiwmObp5N3b959doAUlydjzRWZfFsJWAMUNU4CA0UkHaqVu/+faKtRbx+m2YrBTW3apX2mf+G
1Y3tIz65qwIEDk+jPztQxkH+EvXW61xa4AwjNdqa3d19SHZnKUBg7HF+CIX7KcU1NXG6OWe0ExEx
QeLKq36InVjo3dD8TXVv26Sxo4OyXciwyXRthJWvN3WC/FT5U6m/cmJGEa0660NyHAPQ/fNDptbY
Ebs77O0CKtpQZEtW3bKLGlWmJAfiTqZ3i66tMa2JQY77gDbslrh21G6Sd1DNX/X+j6OXCjsNU+f0
euXk77GWev6wlUAKFQf3Q/Jc3YLs+05dQqRwL3jOVGdWHRJxWYE2Q5D0JhlJQN0nLVyfflj9P18N
4JSdQSEnDG2kipKc6xlAg54aohOy29gfYZO5/Xq0CvLXE/oO6lJAvyC+nGQyk8ced9gmcAD87yL/
6KeZeDVi+q4fusb0l0yJxbBgCY5A702vX9hHhYkSL/g3mMQifhpz7Kc8tnyGeyli9G47X6LgOE9X
Lln0fv1bNKAJtCw+DXCjuXsGxQtGdo19erPOMvK2jZlYKkZffyaLVAeeCXas2Hxx05PZmmOb4DXe
HEkj6Uiw0adbCnJOF7xuNA9ea7la9LUGjTxVMu1ejQZVHwoJDArabhAdNWM0kbGcospDYZtAcGaU
c0qo+IWAp7zAbeTJV2bS2a7GkICDLk8BD7ySJ3TZIABhHrv0qSy4kz89JeTzO4dWmTq+51ZL/2xF
FIrz4mKx7aSNDjZPkvQPvz77t7YuaLWtcSMD1zIBYUIxnYUd6WvY++bm4GJRKTevMG6nwLBgboEL
vZ5X3gtmTroI94i9fgjIoWjtqc3966iAV5PYAOZuzZCqJrhGzUJ7y7U4LnUspgg7GxHY/8eB+nyy
kSzsW2HZ7H03yX45t9fTYWpZjKNIY9uvozUnrT+aek9GC6mWax1FLnXn2cHiXcO/kaSn2EhbHbZX
8KrvpNCwu9BxhO+zrqcIPqRmdR4rc8YE4pdPEkwPPfBJOd4fao92nr2+bAbu/M27m8BydLgsvJeo
UsRyTF6PxKffD63sVKCtQBIiJGKozz1rz1id4783W7RpkVruLNk/Hdbmx96hLM3z1RCTcEJjdmej
DJtn9Pxf0sigPXL8iQNX2aCkfu6sGaZdaO6jJ1oOZHHQqHA27nLPAWN8H+Ai9cmevVnSy+biishF
uYiJfELXH1FqqUraUej4VfxWPzrgfZhWVV777aIJB0JA9u13PWGIZCBCrT9LNXcNvdrStwWwWr3Y
LeZWPzrixAb5kaFLnvDdNDLTUmjnURG3vKhkMgudB2oMJKSvw+N7U+TXkiGxdHObcDALXbE4hYmr
RKYZiIRXKYinwhNglJbt4KI/8EWubrI6IDppdEU1orR0CMNH04SOwTC4X8q+wryBA9f7+Yo+vvwt
8upnRo9xBJawWjONba8BxMX+NAYdO9vAh4KFy+bDEhAwVZ9O543OFIm2RH3R8VmjbXXUsVLPQg2g
WHGhAtWjm1ZSPTcHc4jj9AqOmZOpX3wcpwV7mGsJQhD3T0Q8suz66VopT9lUk5pYQNdPIf45Wb5l
f87C+wV0bYn4+xOlJPUGeETe9AxO3ssH2po3hqVMa3JkDoEMzzoEw+PmSNBkaNpF/OvzSyagfucX
s/Z2g5wtdysyNXpTfVsBv1PH/xMDVsAa+tKQIcHFr0BzxK2OHGMnMgVKZs6ajHEMyFqztNWGIbSm
PZrcr93p1YgH4VjfPh0Z2HyVF1OtOQiVtZbCeroWRwdbYf9Mkk5YgxvBzAh27FvuhshP9kEtipjY
xek6zJLsfNFjRHgumo+l9NB8P/FqrI2JRHcRJsqfYfWkzl6I2WaLFFdeS9XCvew7K0tvLUt+MrxT
Tt3Cw/ZzsxibSTtJNWjK6JlMs772K7oxUXpKVjlW1fvg3Nqs+KWqs0L2kQnfIJ54bDtO2NuwxmZa
UbYEMt45IfqLya2cU3/CKuy+DluEtLVsDH5FFp8vhzTFpiWq7L9cUmZtFnbTDYDBFyuRIiwAcF3c
2FRohuZX3dLSpRvILHnPLBLB/TKKAMH/gX0m7Zd20Vrf6IhGFtx5DN/x1TCFOW1NuWs94RroHq6r
ThpZNfCGFu+FJ607hQd8jtKCvYZph5g7wegssT2atylHfniR7ZW0mDogq5AHoObGLm9Y/lW+AWsM
8ziwfH/676cxPsu7b99n71AjBG00Cipi+pFSuRXhXGnosn+vtMJG2h00BdasmtAnMNzeTpjvipg7
9TSzjph2XyXwK6oZITkWGAv4oRAfDgHEOIz2UQSxMfqf2p7cZuECJdohe+hWoZGexN6mlTqgqGVs
e8UQieOFS6j1xmnfKNNmXy1VYlem9UPf6iLh8kjOBsTeqim0WS0qe5tfxdPHOv+j+QfqjF1dceJc
LGlJE2cOJZIsbWFwpO3hEdj36HfYMtL/vNhXg1h8wZYx4W9rsocaeVuPZL9Rg5+HHbOPWgUkRvXi
7gVdhj+41xWyWMEgqrZfxuIT03cEL2CfXSvw28+p1QkHPT8qePvFbgV4TeHeyQjSTQPafPyaiBSP
cveoxQYMMxAzaHi9vJ7TMLNwnnd2fPmNz23Z4zRYqcLLT0me3gG+S14QQDsHX09bcjgoz1/EQI8h
/pUho9q8hs3JLHNRgNwlgu97Ia1lCZ6UMBZ/A9JJJllf5+dN8Z0i46wV+H54SbfhN6lzbZR7YYLW
RRCUVxUCI+5mQKSRe6Dpi4To8fU7F71EUfEenWGlj5/zlkrR8fcq7XOYuHnZdArMNKkZqRuMVRQd
4ztqy+oFEdnlHGoqsEU5EDBXYwsyn2tZMxptcr24jlv9OCwS623Gtxr+iQK8H2ysIQATZnT3HPow
6dhFNNZHE6xCoyRvWjaZKVq3+V6jXb7DNaJH9ShsapGACGzpncfyXH0bDAd7oMvEQWsY7SU0d4/y
og+ZiqKmjymyY2ZbLUiH3hjySIimltPlEMVD9AeRKzSZdnEn5AabpEjA0mTMJTAWysM1CgYOpeSf
xlSpIVIbbyw6mft80dW0h6AIW2NOtKQQ8bPTJ5mnqjpNdg1Y4EQJNSM4TWu23L0vb9BYpRU+sGzF
7E2EW1g+XGh2fFYNK33dbi8lTfNVJQTUOKBeh9sRxDsiYZHv0zX28t2GeS4Y1m4CuNaQkPoY3ait
bxO57m0oZ3YZ1FzlLLacBHYYYiZP8UoCZyTBdVQ7FU5DlrMtDkG/WoFnfGRvCX8EoGIMB8T/1SXD
cKM7NjRYmJeYyb6zgCDPpFliuYu1wKr07RmSrlv2OBmS9CuGtZkNRtssCj9nMZkru1NzNLHLNxYz
hcMeEVgxGsldz6BAaedx+YaPi+24mP6qYYkf6Ysv32MWEAsBOSUAjQimU6EnbnrucpmsoWiuFl5g
5qN5m4MpWYvy5hhvrbMCjoV3X02yKbDuGk53AOEx8SLD/1qOHWGVrN2hDx0c+xuxcODUAoeGcT5o
NgQDF1Y//iJdtu+kVeWynsDZeZreFzvAqirjFT06uhOL/DeXbxzNTdVW/EVE4X8kHb0ZiTrZjOgn
2nIPVtB0nYhBooIhu3+/MJfyLzWGrgp8gFLPg51gNs4SrNMB6VV/V5BDk9kd2tl8ozZ9AcOzN/sj
derI86hVJ86SAdEKECFEFUFyfcbEQY3wTeOPxplhk2eXce3sI3flzjVxw18ENg2AcGeVbGP2wVDm
eDg8+NlO4Kr3eBpf/TkdiEarl/I3vPBS9yvMa/yAmeT+gjeox22VqZWuqvR6/2aYnzrK2JB8TzlO
clwl6VtBJQIEY/4iPg2snnsJaQc+mF8RfrCvzoIbbNVtvgcBaklDDsw8of3Z70k+QLdU36cLn/KE
rgKX0KdQEHpZSbIIUc+2Dmw6skjvSLGnYyfdxN5gzIllRPd7neMBPy8WIF6T4a8Rky9Z7bB/BsgZ
sr4nR8Y5lzlkx134nDpVPF+CqAe7QoztyoTdIGhu02+zvm97CpNA6f1LcAz7Fo4A1VDv+ochVnUK
NQT5ti64ewVtpzWR4LtyGy9rHa0KaRKmLYncqCGKWbQRzhZuBHdVVWJdrjAJkqlyCP6rj1gMRqvJ
ao+5Z9pkL8yYIFG0sN27eJKqb1g2G0DlQZhgmdex98FbobnSQ4CZu3/+al01ifH6ODv61zZqNJ0r
nrORPI7hZd7JnxzU+/NBYyg02ku95jyrj9KLaUYnzhkRSfRsA+wYfVoW3mpqufz7n8yuVOIs8p9E
wKNdQlAZAH7gyv4vccXFqQE8qVmCdaBH4+0ZH2RDiOuFnze+U4iMwf6h3jd9ep100xOjaficbbGU
zcI6WYioTaDZPJotBqtXtIQk/E/8G925vRrLM6RTNecO1+ouqFqnAw3ukzg4yw6Xgc8AN5JqWqO7
whlCsMGOss8zHr8NqjqYilRLmP/t94tW5Ls1SnaGT//jBDpkT/pZwArs9eilrDXq6V/G9HzRmyXV
M/7p/WoxZUERu2xALcx2hI/si4wleoLgbj3XuyBXrPn373oxh5sjY2pMpsBozIa992dFvw8qsNSn
gl4Y2gXiM293nAW4vvtt7K2xaukmlpHbo34p6pMJ4nlADuw8HB9yzwSMvuS3RfEUZ0kwWxsZoOrR
TJcDzzcxpwHscCSsZGgrOaPdO+QKg6ZLFT4UyISwyOr3w/CgNs8EYh2lMNsAlCAStv/5Oc6RVrJa
EDdfF2gHREcPkaxysceRnKbxBlxD/5zvA0t/HF9H5ccdWv6HDnrJKbRZdFp3NAjEDQSk5zA/Xy2Z
BNZXXBPszgpkVQ4lcmTfwslVDXa8lpigudfPlrF5MEQPE27LWrEd9+O8utak3dqpxePghhkUK1rE
h7NGJTZW8ZbXzyhVE+5muiclLOO9lLPFCqZSPJHxt3o4SXNdVaEm25XI/qTABYhMjkaHk9YTJQZa
fOopOH1podUWM88dX3McR2/PEVYQNG99WZVKXSIXNQUQFsiYYOcNAEyamR2S69FAeag5crn5R5Nn
T5jGg/GoYgiY2d0uMTYicfkVeSIpeCwppGRa4Nuui3ea1v6Nh7hdY4DU19rvsgAZToYHSSVY8dQh
VIEkraCPbzcfH3zLPOkCMOGEYlnZqzQXQA63RWt+s7dh+Ca3PGQ9gMBe8sMa7PiUBswlzQ4F6Lrb
V7SOgUD//G4s3aLbv2fkc6MNzp9DsutpXN2FuBctX8eLPnT0H4FUSXNQVwawgsF3WMUPOes1Hh6j
PypEmJzsyvXcI+U8AHgd6NP+/QlX95XbFmE+QZWICRm9e2FPzi/FaK/D6rTBmV0khJPFiECe1saB
q+hZQ3jb/NAQqRSVGmiOqUMdwzpKUcasKg+oexqTVi2ljlMNtT2O9winO9VUuyV2UBRnlnB5RlD3
toBhFt7TmNTIbTBGVZS40pZ+jBuU0e0mg6Ay3frHJ4V1kw91EngVR0e7v+nJTSVOhAmSgS71Cdp/
d6haxKqyUBl+/i9icxSkbwA8Qq7TYq/CNZtaEUxYmros6wV3erhgjhu/SE9q2RqQ+nJuXz+YShWT
5chYTxWmomhHU1a8zW22DSRnd3m4/NdSpuoLF0hxKoIT91ty6ZiE8A2QSgUw6iVBTv3sVxhccj0K
kh8dKaqvmse9+voyu3Cyxz7iJ25031Od1LKaPwBvSnB3FRmKqq/aRL3mb8EYfVL/IExn7aGXwv4y
LbP+a7z+HkMpsM0LDcoFn8irE3Z0vRyLVbz5RqjfMfb3CHxZ4pkGBbGpikmzm9ChZ4WA1affMSII
BVQYTuNgik/wD8MX99nZyFK2uRySaZ94mCdHvccIhv5NKR//3VgyXb5wKGhyhFYT5hqsf2Mh5ml9
79+xm+adg3JJrnC/WxjKrgewVV8IaC3fI5C3bJrtP8fKoyimuNL/L2AaM59NdHNdMFAPZsTOdpnh
lUVPWd6F671IJAJShKV9bhGR1QCYx4Uf1SRqfRlLMmm8j0kYeaSJOh6eI9rol3BKTWgOqEeJwFQ4
jJHCIAxeKaG3tuhs+UuqDe7waXQp7RBo5IcC1xl+WxPz+qq/eBql9fmd4egoLzeo5lItfAayoTmN
NTTHPvratdeQbhHX0mBu4QtOEIuw2ENtZT9HfiawJppSOyfZrrbLuIldDT/76cIZdWe0+YRM+Idy
zooaLHOO8seZMVlI4WgxJM81rPSV5jfFCEI3D/O/FVi+EtbfKf1gcRMM72cFtXjhrDfZ7VESSHah
2c5gwwkYwekzNsi0+Nnc7sK+h0TD4vsvZLoTOR/qZiHzhztkI57oahkVlcv+ZL/N9AfAimDFH6um
eTuXhktpD9LsH6WZNppsrVyWVDQPqg7PtAkPi4piy0L9LKfLPugpKs9QMPhz+S6VIellHmrZwjv2
i6WAOlP/7h4O4SG58Hesqti3WmPuFN+lJWgEBA0j7Oh9R+fyOTH7V5D/ZjR/w5GBpiokGdzdHN5I
Nh/P1pfpp0kOUtdG8o7JKtK+GEQNMxRuOmIIGM7f7sK5gMqzonoh2TdvSmg/ff6eiUC/nGEiacH+
ASKWGSoSd168FIeiBejvfjhSovU6lmCrbOhg41HCXap7JeI7dwPCelbck1DfyVi0qoRXebhswtlJ
Jbb9+iRFSpjzkX8MApQIQuDXec4mYrQ56OtwJ6IezmYd+NPraVr58t7ZMdWigXZXngy0UglNjyJA
dvw+fnCFx5rxOKoGs8d5dAfD71wEV/v4OlU1/47vNNh0ZFvpaJembZgrlhIAmlAur1bSYeJLakS2
Ucz/nkLWAwjUVNHylWnclzkv/O/p9HJCiN2hckMT4ADmpFYgIBWFVdZO8Os61jkl3FS1kaSkSvYQ
mU6GizdmNj/XMzvOg0z9L81zX1kUF9S4APjJutYVArY7n9wFrAzc/wxtSkeWDv+RUpHjog9qOSYN
JQ5LjzP5yQmgBXily6hTrCCdlPCHLEgjBVOgWAL+jkF9/IyDsDPoeYpsEKN3tdX+Zi5OlnC2KMgT
TdZq5hMi3BE6/wXxh5W7+WEKI9/c7sS+xknCyBS2n3RHKqsBCAdoHWBKrg/jHf7Lu00HbTDeRaq4
piuq9HU5o77y4T2WVq+igKShnWB+zWzt6A/4yCUjyj0G3xTd36T/YfuooR+cLFgtXPHyP7KGpHeb
1qgXBJmxMDSQJciztRgz71+qLQTxaeYlC4+tOQYoLEYtssL/wavEXPenJZbvgapE+AeXMpiCok/k
GdCtzswcId7doQb2RMdJsGdCj3vqF9O5m7kMGvNKjDPAzNdJsNFWj+Kpx0fSkUH2jmnDSPUwNl3d
7dT9YUtvc0Wyz4sg7djH7Ai4zdoRDoiQPQdgB63wzPYrrU8aNJDArucNiXW2gFOb7P8AV7Dck1Nh
iwBMKsMtTnFg6hVWqbaSV3oP4FuqcOOS2i6LMKs6wrzxRzK2XoqEa6vz6ksn3AnosYQ/FUArMkq3
FoY2iDyAQQqhyEGY6AW8m3ajYWDwxS3642X87Ct1wbR0P+Yw+G69fsMpbZ7glUx0qVX8rD/URJDq
BvMOHp35+xIDA0+jN6j9HG9IUM88cfPtaaYsHSrj5SGgNzqNFCEo7iiRAknnMPHx8XEl89L6Y7Pv
koAFDYxQdePMtiDu2vw7giqZSPxfhubUsvO4wZiNRt+YdwlebcWYQS6HEPdDT3oS+nOhKVljwNFL
8V1uEijPJ3koON2Wdut8BcoKsptTERA5rvwe89/Ai68IpqN8okisDQQMYOIIuCXDGTJKfKpSSPR+
54znCvPEsXgsyk7Vd5XvUooNXbWc02PTOvZAg9IYdWkJAnD5mJUK4ajeM0ypRwb9NTc4X48MNLQi
nyZAWO8jUsysLpB6WUwQoTPsS5KE//uNCRJJmKAkBQ7yAiD+3O4WXp9axJTnUhzm2XajvvTFYnmK
clXQI6ADV+FY4AdHyMUPHiw7s2yqPsgt1BrovhdubWuCjXU+IKh/Z4T+eCA9X6A5iKXX3OL/ngH1
56EnCWINg447YcEVYyQMahTV1v+el0riz90yFQCwyge8YTGw//mkNwC6GgRBVyD7MzSYAZQOXJuA
E4PZLgiHoI/tJuPo4h94dbdQ/dq209Xr7o3Un5Tts2GuoUhLLaRhSQ6mxVDx2HMsLR0CPQd2OTqn
DYN154DA6lFA6g58KYd2x+n4JdIgW78Zd7Gwh7502Ldu6b0QQqUkP8uRQ7l/kw2rhjb/S1eu37pj
+UDiF2bpm6fxAz/9Wtws4iyE8G7aQno4MleevAzOkggbi4i3pNkE7/vY3no4AbBLMw3oA8Napzyt
SYyLDUMfbQpOmBy5EwXonKh7dpKsnLcwUkUSNbujmoPCt1RPTYRoB0OwVQMOq35aKyq4TTTK0O5P
rEoXO5PyIQ5+Am9ceFoUY+ovQ5fIrrQWbDlhKxz6OAC1FFR8xpPkbOklnC5wpWxgvYL1fbshiY2e
eywXtwVlN2wnYoZ/ufYmtCtP46WUn/WAVQt4AskEPcBpsbfpJDQhRQKKo8VrOhJd8wKgoki88286
Dkwd9OhKnDpdUdhuYlZ1+dmQWbnyK/jtrcGWPHb/+4tRNRQ8x8t9vGow7MBqUQYz6HVySS3uhUGe
MozPtsiukLLAz9aysrLf1kEObMyzapk0TN7TMA+bDARXAVPZUedAWfA+GRD/sA9oYMduApdYFp4Z
wE/r4rd2pAfxwrqtnfguIbIfUDpJVj3qfi/z9puxCJu+cpofsEjy0RM2LuzQMZsYU4RVXuk1RFUU
bO2+C0vP2gahqZOLwnrWBMoyErNmT3hEcpH3Jvjc7lTfHkq1cV0A1CjkkRomUR+mLdcHgSwyvPqF
Mp/xNhr5z0+QS9YqvFQQYczdpA3wI2acgpjHPkGs2Cn2g9MATjJeWsMuw6O3owhqDIML27KKJKy9
fXk25/A4zNjUQ8yuyUjKMQXEMRj1IeQrmK9Q/To3lvUY3ktu3A2l/KVzhheRvnoyS16jsn/EALaE
JfDr/2TcA9BuWTqlwuQSHSL8kbscJR3QByDn8qZWwLd223LGYezvrgrlvTigWKi8L96iQh6oaLbi
yyOJr5KoMdGa5Il/F1trBqw8MERUWBJIXRY6clMfQAk9iTd6mLf+r67mI+Rpx7o+Y3MIn6/A4n1T
6H4OsChDbkCpvDe9y7Ofrxb2yR3XZ8g7gyzHL/feaN/h/R3Ja7CyFCWrwbf43BAEjiU3BPtNyCj7
NzV/wTcE8Z9fN8FNAh0h6P2vtE5aDyAli+WSerCWucNSu0QVSDS+y86NVM1Q8nGBtEi7VnNbO76v
2YpbVni58VdcOPwndydV+oLR5Ur5ypiDFH8AQfep0qHnYbFiHQpUlOUpRtwb4axuWPYDPUzLtS14
702wCkAUaXQOxY+fBO8X6WvGYTbyvzR2yHwXzgOOJ81XnnP3NAerxG7MH8x2Ydc0DIZru1ikNjr+
DPgrszZFwsI1OHVdILnQbF2CS90dq8JmS72ismlpBZcTpIg8z1i7lYYcBJ+6X6J13Rw8LWTnsMak
BwA5GYh70cg/PghHI8+ppAr+S4wmQ0Fod87j+czE7xfJA2dPRlrPI6H0DgJwM/y6bxt1wEAloLK+
W0Xg04illQUDtxaT/c20QjIOO9fknIsQfDeE4bYxx5KZN6e2Z1JhPIb8hPBMY4CEJgD3p3nL/CFU
tnobr7hoY/14QzHTD7NsvHdICf1hEG5zQhIWXqwC/gAJ2eV3+8DeG9i/qhniX+M69cdH7xAZGZc6
aTgbB7i9qs2eMmPOw+Cg99BSIumDMeQDHXIJ5knIttkEuQjtkLo1bE2HlSv4NQ5wMGxfOuzUUFHt
amu8XN+8v1qLBfaoYCgfPlmD8E21vL8f7mubOthEWUmAJ9pOchKz4uLRMe1/MTB8hqtrRbKoiFQa
h6fPRi1XP3HWlnyQ/swXiMf1W0F6Lkexup2A/6L19LUcWyhkQufkTp2sYxFTmnaPm4CwuD4YPvS6
VENgjwpZzBjVpvkNxMw+zHXnwEpNU/Do8heu24Fd7RcM9ZQnCOmdR8A1TxYtoerObIwPAO3U9dbb
SKtJ37VeSFRF2YVFgTbA38l4suoHV1noqN6QVco+DDTvSC/DVS7bQYdetT/8f0flLa1VZf251ByI
7w0ipZyY8I7ZRIQzjIrFGIhH5LeAAdj6k/GVQ89GAmKkhoVN9xONxiVr2HEVzkJ30aDnW86UVRsw
7b73Q9UY4mLvql8Us7QQHjvGjOpm6MBB0hS47HMLgzy4ki8KLPIT0GoZfffvB1LMJJ5rr9W4Olyk
HKgzSLmWXJ9gigpCfJSHDbkmQcnmNkQaYwTFg8yk7lB9s0rFkwx861WMYfrMH8Kkt4LqUweEjSuI
QRLQlFfQli29ozrMGl74QfAk9is2fJQFvGj58L4Y1Ep1+LyWISrpNx8wirypoEUTN60RtYq9MKWl
nwb5/C5ZuV2hMLQIcIecdMG9GhrUyT/UoDpZ438MWZ5YfVXGTn5RzXmVh85OdJnm7JH+ysJjwSAh
vpQxgq6xNK48QjhhrUwbV8GazjA5tngCKNPNxB7+hBatKCPfWJus+2j1PPKDzvEBvllq2supWpKP
o3tqoW5d7X1UxiRSTfwVqt6Dc1VUuJwPozFj+C6K0a5CUTO50RaYmByko/s/NjhaykR3W1fundy8
+0mn0rpC1m1wJ5+vwO79JKl7JcIMdacfLSjbLv0hTsrQw5wGe4xwa6NnL451sxXBH7bi3GsWDqMZ
VHixBRwkcOl8g3xBRbco9dCIFJzXh0Wv21kvRxuuA6VSY1knLrSor3CsG5uOho71x6NgcWhMcHU9
cWoMv6x2PYl3uUHNR6oww6RkhdnCR45cbk9oUKqs87VIyJEK/7FXJmyQBPklUqMgx1b4XUK4VIuF
37oCv/a+/Ffo/b+cHZdxVGdeJTIJ35lOVJEDvIbmlqFZQutnJQ/F4mS8ayASMGz7rBLVa7KEP/yo
+/fDkSfg2DaODQ6nsHh04wm/M9ZviyDfuwnQ6tvHoN76UhvO58ZARAI+XEgxpzeLEgnYj1n8reOE
Pe6PPMyEdD/ODSHe/wUVUKTWZCHEtPSK5fFGRkDp+E0LyXPE+AmDPjyqVD/+nPIDiCVR84ILOtj4
ZegyKloxQjQvCOA2qacWVTiPQ8mlInM8YR/He8I9ed1BvYjHY85LNYPQ61SG1dBk4IV/sNIDOu1j
x80cgGeGlDSAIT3jsyMy57b6nBZV6QS9EbdGq3hTXnMoftZJQ2x2+JWgVyiF118PRYYDzSHDDOEZ
iipXN78F+uHPJQsReykBgutMOe8MefXCMun5lT0wvuRnZmEp3LcyLOUWTNMfVwt3mVjrBEguCgxv
WAZ7kP+82f03l3th/Jro05Eh19vealONR1NnDb90Zd+POnrg8zM2XED94HLIJAsjBWb5jTmw4crm
P54loMc0+Jupov13+mI5HbuQTR6rXc1jCKohE9R5GIBotufBPCb7/Fz3O7Mfx1q5/yWmLgSdUMdz
JneckDOE6RCgK+My556oXbfrZWAWsUn7LNfizfG5Wu20jLaLA1Ea8j08ru1Yws24MRdOO/udLZDQ
j/v8VG8THRjZLKtZbp3q+AS+KZvxyLFriOhz7jYMvjQ4G28BabKBu1/PByz54J/6VDyvOLEopGBx
pnk1UaKnMzK2VjSombbluztw5CYXPX6sVWRxhcgcivSXyn0OUAaFi0IiVrpJQBrlO4bRQe4JNNbS
r+E/PCD6+BSdHqo0tNzIe1QXWRYdjKxK50DtrDqGfB9NL0yfMLwsZqsE0Z2xrP8FAMPVUPH2F5Sb
CthWecZqOdcXMXIXbqLQa7aVUiqI6RfADfjlTf8U5HoawMjBnZDjUJueogM+MZwx8jUPaoyfFFFv
NtnWg+0wMSrhPZI724M3BsZosxHXjo29kHcdwr1hiSvhuNfCDVJJqpQB+LWyvMdAlDkwmzpNK68i
I0oTiX4+VWIlHjxfZ3ev4GialVj0x5Hqpycmqs1QPYpCNXNFcHj5DeKA5TPomGGsTwHYhl+Nun8z
8Nb/0xCvHmTykH9lXRZ2Y0yJ7c5bqTeUqjs4phgwARCGoKrQ8kNLZEiWwcSKjgayeVvP6m5zhwN5
Vj7y0jmtm75JMYGSBsalQ8BHsdEM6wjmA/Dm2KiT5aa5LWOuE4muqnMlhA2W2iM/ekkQaQmF5uvM
FDhXy2ZOwlWFLZqHzLO3rIUepn9e/GhoWXPqEb2VnRCILUxpAZVuSQOEw5x7rlgQs0GQtLBBz+eE
ShFOhUay2/AMJqsPYyyO836aYtu+CjoEjFPGGxBJxLuJA6b3QbQMRh+Q45j13X3DfKzH9KXKvVfl
ueAbak3SgGPJ/sJZoU7GBmIFu39uMfCmKrz3OqSaU8CcoTer+a1JpIcXl7YlhVLxhDZcGAjktXP5
UWrarMpoz5sf2IOJNwDvLlMiO0+TZAHRremcJwB1JvSYIxaLz2gPnQWydXwTIjVjAyN44ABsH77x
Ua/pMELI1v9kT0AUGx/DJyK5AM28ImlyxeQ+qngZTzNLZz6BHXCcejylnTbgfbe4cZgfi0J8iLDk
L9rHGwxXWTmhChVbL2sBxOkx+QzKM8vWEPRlGZr0RI1fTN3K6v4d7EZ/LCGmxC8qLBf186PtPu3P
grO345qyQxTTtSyUwLfnaR1b4My36GdfLy1CA73zAECoAg5p6sEEV42CSj0s8TDfwxyW6WaZnHc4
QJ5kpSdUKTd+eRL3r78uQUbBH4AkFw8HNVawcaCoRmRQBAguahvMq4gdHLz0KDkPMz9MBGru45EZ
MHwnBY9y4ruyoCVNCMUsulZvgdG4XCi0X+VywUAPHiwI4g9utA3rjSciV/4Yd4HgmbIVomTVQf8P
oUHNbsUZiJ/vDTh7aAJlAx9c4tJ2qcO6+ex7vwaVqD+qGFqb0ln1LyPF9K/fX4BCiSZM9EmG+72q
X1ThVNd9+yePD9Xw7GTK6mGai2tPeW2y8yx1jdH4VzatDAE8nhSM9DHnHOui47zE2YE5wEA/kMfb
MjKcMqirkKYZKOJrsVOQEQR9OWmGiPBLzXFd9GPXtORZTqXm8tI/PT65KdRdnN+CPa1Iczh2403K
RFf26r/cPa/CJWigpg+YGW98Y3vhylH59DEzh1R2xD0jm50SAnoauGaO8JRzGFLKQJAZf15PPOIN
EZvJ4oOQvZyka6B1SN/BMLr2ttmqnmHDQpUxdfq0gOZhpOG7fuibZ1L2rLnBfN/exGDKFjhbqUJI
6kB/XYiteuOttT7TiPsusfPml1txkFuRtJtU9BY4P0bNH/xtzFLXIl9KpfausiGKq74jdMvwDPpG
DcwrfAuT4JtPE2nukfWoqEqONY5Tdt/vZVpHyOMbdD3TigonMk/oKMuulQBtBGAegKhUEUEgmBfS
i6tlQUS2CjlFwPUnieoW2o/CUhcw70JclqvbWqtHSCRr7cSXN01FFwolVZXIWWLPsMFW191YGufp
UoZ2AgSCnxb+t3bAGeeXzudBiYYR7R/sxc8qxSzmVe3Ir4LlywOFiMMBEAa5srPgKd5BxSdNJvMr
IJI0eyNAxHw2P2XTIfeOGeLqkI3QFPfjyIHu7meWNHbi3WUX9yf0rvN8FmjLKBCBtvSiG675/tT1
HUslS8hZt4gJMJJrUc8rEgEpUFKTC3anheopHoBaW0iEgbxww7L00SPZAniMOdXt45zugUw0X3W8
ruYiG7mlch7GYghccS04lKOCpxOzopWa8OAnzHH2m2GSZf7y19WdEoXRCr9ZAVxIpXoQi5ql5hTc
9ogHVOWLWhCaYv3YrOz48hVYwIJwVK6uDLJUul6wQePqU/lPtkTZOSqlAUPD46rmIaiIL35+j7Yl
39XedkIMk+exmukR9JEiqeW9Q5/dlu6XJN+WatLc0tsf/AiVlD6xzLfYj+YnYwfaagyHCTqQRI5x
ibMegfzFoJMvoX+Ou0b+S33iGF3LDNrsvNrsj2bwnuQygIcGmGF8wYDIUq/mSt7LV3OZCVWX3zOZ
Fu7ob1lPcWjn2d922/xkNegMULFr+3eekYhLxgtUSgB+A4NAfkA0XQuJ3Rd1L9lnBDe9cIM3cPMt
rrBX4eOGPHg+y1oy9lEhMA5ydjwDwlzAXxFIvK5RslAS+8MWZk+Qqeb5HPXUmqTjpdtZdx2IGe10
foSQ0nHqCMPltqWeV21xar/m4LvBmm8YFdqzMc1WLKF6UU6PJ5znaiy1xUz+U6+kCn9+nNOhY1IA
+uGgZqOG4PufLZtPxWhOGhcfXInibhUebk2N+anAt5ASAHR45BZHSBIuZRflo5X0W4Vr/wu4j9fX
DWmD8t+SetWxhOB9bLVgq3W2LfssPoQ4uu4dCmG3Sbku4SO3L+57hO/9NOjfDncw0/D4CZ0FMmzl
sf+7YbbOmPgDsFHZmoIYPeLKWnMOZ9tr7a4rJkt6tN6FzcJSLqw+Xk63BYm37u55bUcMRhPz43PD
3mWyzHQc/Hh0F31ur2KJZD9/ov5wQ+6Vy30Si76ZPJLHWSJB/po7phhLnB8lc4pN7kCkhbb0MNts
8s05NaX2VRn1mituFIy72yWr3aiBBl32B2oq8vmpVi3KfNRMokxO0KFcVGinUjGsKoThXdYnCQVj
HQFtG3iISchK60y6PPyxwDoBSCZ6qrH9GJs+xZcwjK+XIw8glP6gD/3bqReL/ChxhXtfgn2MWze7
GuD8VuO03ddYf03ny76y+71frBL6SUJs/PQBcQfgKSyrmc1u10ixEk2yC/KR3kyLLprs3RE3lDrI
60I5K49pOeeQPf0vdfcliy0MSXh6uqwYTh56S0Bxj//6zhn0EP9Fsdhrl7UNXfxfTkSewddAkqRA
nvRCPq0Zdh2JGtaY5ubIgACDzjPH8itpzy823zwkzW1qVC0JVAGWI+DNoF9ArDw8LAsA8Ex+FsV3
F4z0vq22Nbi0RkntzAPOmTR+D073gq90jf7i7MBr2vaydKQAr1TQif7D9Y7JOfaqYxj3DbVkqs+X
kKpW5SwTeLtCSNnhYPbx/V4dINl8wF/0VWmmdZSZaMbpRjv6th2SBPBN1yKLbCTp3/blLED9rA96
R1/UWykcueqIjhlTZB0ZHCcIk2zDLipI/G2kYFyvFGaxZoWcOEHN0bV6BmHQ27K1RehKgdlZ1CHF
lyiWvOEEPUuW4nPdjJfWOrjrvfd2O3ADbFtbMs5jTro5vmZexLBps1b3Kph30wwJ+Ny7p7ZDvyhM
g24NOuOHuUazG+n60BWr7biNbDr6uCpI402K0AlKmpvYqT9FsHZXrXFdc5ihnBf7vRoytCU2i7Hz
WVlineaiZEDu0BNSrLtwU5widdrUGQyc8xrsgtFtAr4b3Gw8Lp0HrLcpGkBFbIpTx2hZyEZHbnwL
NS9qetqZfy6VkroK3A3hEgqtgvPCRkkrtOfhQg4/I0Nf3ICU9/0IkDBV+VKXVvuFqA3G0ncSUWDB
tuLUOsaSjJOMsw9XHQJU9r+MGYhLfBxqmr2qeSbMf5psx3XYjomJ+bpGOCzN/FvG960Jtgpvn1ac
BF3Br+qgxl1RnBmJhveEmMrqMNEL9+Sgis+OMZ84IJosZJ9vmr5wuv7iH1/lNZc1n6nQCrNonB8L
FOwqN347OVmY9QrGnUgnb5D4zdQcG3Yb/qXUn1H1xPvuFFqqytS64G7isIY2yXNPtYWEhoy3/J5p
VV5CIOon/P1L+0nG4AHkgd40dfBhj7vHEICUG77+UGrWhbNmdW/FIsgon57jeSrIhJRlWD9IuSLj
lvbu4pPH4a/J4Vz3iIXBiOHABbyKAywyV5jwB7OjKEuNxb/MIaCN1f7EJ3kKdz7yvWVbIQySXa/k
v+3AO92Yqzy1HqvhC7hK77l9m7oIwUmvTKkLdzfi8EEXzfAqwgfl8DloIRVjlTtYcekg5QW+iY4M
XSXuAk1E568S8sRhtG6P09nIAmrBFZ7WnfmA6PdbBIv2JyStccrbutrlHA5DtZbkqwnShtMvMXe5
67mswmDwkND6qjHwT+myeJ2iZtnjHkE8NFIwgH7YAJNgNw/4c4WBFczMeVCv9gdrFMbzLgIL98ds
c331R1gEPV7LN18IKyRS0GDOgWdLToKDqyaV1s+/Jj3NTiI5dsQpajV2rL+d9dZzEAmzGKu2BqQN
UYtCHHQIiDss57avPFg5r0j+d7SMKiTY+wCbKfTw1JqR631Jv1kVQ5+jH612ZJ5eqHQ5sh7FVGnB
UY+7gRGx69vJ5a7wZfSMUSaodo39nasJBttabyJdp6ERYAZm9whlVhI+9eT1ZWLRwteZ3VHeyf7I
3TkhW5XCrsDJnhmyiXX/KZCm/Qfx6bUK9pxAWHwmtyhOVAi/JXEi+2ds8wsLxHsUbf1CHImcsOLH
GckY35fbpj3sR+QaArKbqD3iSfIXtnqqy3GQ2P1ZY+yq82au3cpRBhSCsMHN1QMM+1fsaREu3McO
BnNaGlxdIkxf9R5V/3rWaycCS1S8eOnd4s2XwD3+TrPba8aTsJYuSkoGhqj1b1FPaVYaVM49pT2t
yu8AMmV8825WLyDnXNzJ1ejSpyA0QBLk7HaRt7ipdo3b6X8cyB25volvLy6aPYWD1moZnGvC6rw9
v94iDj1pGloHU1QK4ax01scKpmz/8tkb+P//lvy7y5bUHE67vDM2STnipEU4AQHY4Cnp24yM+90d
C19e3cGk1nscXlHCxywdX1E6Rvylk+GFOg+14S4cqzsXv05Qs9dcdaDSLfxOBGYhneH4d/ymgJyK
P/wjb++aru3hnvFfueHJJncIZERJOIqMie6GOBmBNcmk3512xWXo3XfDNq6rsThtQ4mQ0ZS8U37Q
RrByLId7iyMV4kXviKSZjg5Ywl3f1YjQB4RnDchamHC36bLj9cTYjMwfBu+kdcc6+eBofRzFPIu9
iyzXniJCLVrBx9VB5qxTHrBGqrOmIMjAmaFPPENplWEhe4xDtc0LDZYZ67BKQANUBPhza1MC5thl
s14T6mnEmWtTvMHzpQzZvW/LZNe27OIUhtBQPHCBMgh5b45mKIbHHfgyQanCDQTjo4rFJ8MOuO7F
zsp0vgkVRlQBczrmFGS7CBhjqtfC/Wv3Ma5ECl7blplg22yEQVUcOS7O6XkLkJt/iWE8we/zv7fD
yarI/3D2TqRiTbBmiqBkyViQWtoIHhIkoNPZLO6Xh/8bPA2Hcos1ZDQfbK1dJn78DOHvQFBEmJ0y
OsaMITNyVz15jX++oM0IcieJq8Yf0mDoOf7LcN8ug1uZaFzLbmde9sMn+OgO4jyX/uuWV2OuY52K
6Hk+F6ZZUmq2vmbfcWbtKxnNxMcuNiZDI27No/6H2SZxiaDwQDW84scmofZqnvjPesA1T4H1JE6d
LLkhOspN33fvf/eGQ7TkiG/xWk9RpDIBj6M9CYWwLKZ0JISZb+AKR9hbYSX0wNRl9+1P0IeGzqlS
I/jDD1+CzzSn/bESxlx1OiMovxKMAb5nshhu7ZBG8/igXMVqnnLpZ71HBekzSF/NwitwN+Fq9Alf
Y1WSjC+TdVDbUkRqhZXq4hHFJBKbAYc8aMEjotPzNvL/eaQSNQySRcOatmImhGSlsRxNkRMUFvwS
V6SjKZXXAtwQGS3ngsRAv/gyII1oiconu/BGjKBHIUuLxsOlm3A7TqMw2oEaeVem2gGbwQqmoADg
1U+hKQ2Q2w24aMMpRJV3Xhe/D2rzNbYViAh9DW+fyEx45BMIS+GWSShTmiXsThn7WTlLFGJWwWY4
ltCyEGRLTXvT6HhF6V8xpCZodOeX2zOUm7XBgoRahMi7JNh1AG2m/siZSMEM4rklr+YJQ+kuWwAY
5RDWyKztZVC7Hx9pT7JGrGLX3IPpNNS/a+LYASe16YArBf9EdfM5bRfoIQ2aTU6a1V6qXBNxCCKE
CGZ/vRCCIu4aBb8w6xxE+4Vu4549BvsChVcH6ya03rQrdZdKHCh6MBUvgR2BTeJeCD9tzZZuOFSS
8Zhu0uzAVkv2gRjCUrXF3+GlXYwnuXcJA0367Gs1tbjhB1EBKoG0LlKz+dzYJb2bVuus18D57Vaz
Bekke/kLsKsTY0locPhsoNZc7/g+BpxqrJN26HFTBRhkNR7BlZiTP0y2+z9XKSqz6r+eyMu0gDkr
ljIlBE7nvMaifiVWmqs4NTPZKjcAKcZxEZptLEwJuwiVemTRAmJFQ9ak90/q0hrqUMcw+6s/+O/G
eiriBeBQHzAkxw0WrFyIUDklnManGQ4zIh5G4D4mgE3g3dGCT02HyY1wZ069QjTkwSdxKkJkeaGH
R+UZORF600uBx9QodAxwzCPv5bp64rJYGYUoqNpGov42xYZP7b/h7cTo1R5jSrvUk6Uaq2Uir0QE
ot3IY06bo2ZUoJsCoShpv9C1xNEsJ1fcKbk+io2aT9il6kN/daqhsKzFkCD+GIvP/Bn43ulBafTT
VHbz0FA46q/VDb4F0PhK1VzVhhkEMsvYWl16/PIj+QtjMtXwDZ0Kd/qde2GiZMDq2lCj7cPH5sd6
6/J9cDHrPb+0dB5CERl6cpuass9u9mRgtu3Gpn0pNPeeIilQBGawIoQ9+PYUWllbVIgUKRyrL9VU
Ldc+F5XoJgYUPiEl0DhzwBc+sf3BJ9GufhGYaJ3/CNPdl9/ms82bYuo23M48IZ6ousnu1yS8mVVs
dGb2oW+BwO7vJy2PTkUMa/dYNcmE33TTuLWzTXIdOumAQwqleJE3FfHv8jGoxFhDQWcTKg11aGM7
bS9mHtYqVA3Q+sngI508ZGR+qL7mow8piFluDlT1fhE3R0behn4lx94Tqdx0b4o4PXqPEPdRMOca
GOK3rcaKTcioIZO0BKTvmQErmDMLKcD0W15hLak2QwB8rU+qcmbcSVOf0Y59DQAKHcWp3gmThscO
2mTvYvy9ZgFdtPNRdu8jvk9sybsgmIxQnNLJKlPkXN1EqHwBfzIAhoh6RVWv+vYEA9Wb47ewZ5dG
LK/hdz0tPsQkQTLTO6UUc8WHExHlFMsbUrTD95BTKgVLO4jtHQ6s/wNEQCNb+mXTMctmU4tgWvgi
b/+j6o5+RUNCB7TC1qUXq46DdXo1JCF36q97m2NsqYFL0NPv+/Byo2NPL1S1x2ZigWRudkmiPOrP
VCt0ICat8+BL7WDdT7N848w3A8Jxm8FsYea3UHyrEbNhazU7SKzC3bC92vgsrSuWIkQdZo7IdokK
8NmuM/SvGPCsle9GnmvhK4g1YTy2NUO/F4ZyjKA4WWk2KmwQaMyYhzEmXOe3C6SZmj1FikHGpR9e
9BwdOeaUfXalIiDjQ4dg1wgEp+SPCweRHWyE0JRDxZJqdZ7n5BdHEeHF5Zh3JmkjednveZCRGfx2
foIiz1S1iiDCtLWmkqT8MG9zqGuGlfOkf+jm+czvfqm/1aIZHmrM8cBbsJWSa4h6Z7fgSDYqr1gB
FR1YjfEg8IBzW9A6OIw38ANRcZoUp++6igKkBGyFyYcazgic8tFtwey9CQpnPjPVcYtfobQ00l9I
Eo7hnDB0C4uXHWIxwS7xOpmlELu+ELZWEvPg1CkDHQocagzsOo3V8mrUQ2Uq04YsQQQbk2/fq6eg
WCDBC7/lMmfpuxA952xp0iFBPibF7TlA8iMWslIPIQpAPuhOAlDIkw6K3PjlnUasKd/xf5UWPHLG
yWv3GbDrgfXK9tI5O/JDLHLvWa4yDiNldqooP6DhINqefXyjIfW1Y4+3kY4kuq0CTg3ltiywUDY6
/F61wE+Qp8hxr6Q3S1YZ9vgp3nA15MRnlNxyMCk/TXVuE7O8Fm+iwpj09PJio8EEbyl5wDbHgcBW
zUQjU8no/xwlHcvtTmYxg4pAWBy1KLp96Sxm+TGekSU4asLs7VsVcmkI9ckE1JPwOZTCCtu5cztj
RdJjPTsmjKDvKy41izM7e34xlCZ44BsdtbLI9wzIlO6Z6akAC1vluFcEq9iaPPOsmVhXDcNH+aut
CFV1B1GCendYw6X7cuGWEYt6PU/BNJaL/Qb6xGsEDgaJpV3DPwKpPiBpQMBp5zyjsiJ1zMvrmeH/
tsyKZnoCaPK1f1bzXy2FIIac0b4pLs9Pt5k6jwzuHv2B/8dCwAi3N3kycEYnVH/jGyw2FWWnmomX
4gjHrnH+pC679T+wLV09TRdW5arnt5yDPjqq7rT1vo8eEFL54Rn5Zj1o9G6jUC9L4sPGxuQ5QeKQ
AWJZmkF5v5jlaHp1zthOx+OVdkiXBmE+HSohjDRQPm30Rg6aoLx1xGGEuSspDzVMv0Aub1OYfJl9
M30F/2Nws8YhoiKda6wqywPuatr2cJIltUVrvc+aC7NVGFaQTW3UYKBLx8vkfus8UsfVGRJa3B72
NDQ+PHYWc9V04MwqFFB6e/T95a5qYx784Y6NX2/K8qrDjN0jHAu2w3vPV4MmH5DqnZs9VDa6sQal
xaKpcQ7CEP6K78HxswSQANhT/EF2Azo7EPzLJsuDM+9v4FG5PKMm43oOEjsOU4JDMtHOSRbyVdAE
koBbFYN9DVZ/ZEjStSMeZm1xgrTzwkD90BE3VxL54ygcKplnBazwwjLw2gV/mKn4sUzVEQVKGluc
d4RrtTnYOPluohRU1bqdNP+MAicDOmS2AIVfAEc1/J645ezd0mki4H7cH+c7qu5yBLDRC6pY7cfx
mnzZULhpkCQRLk8cPuDvTWJ35j3LvUQznyX9Pg7mje5R29h40SMR9byYLVS74HMB7SYPvDJ4en6F
sfeHuyC7GNVSopfbXqn83mkAILYgHPTCFtFNsQfnh3RdfjzC843Stpm1Dsy0Fvrht8PFHfRq3Mia
6tztzPnQ/DmnrsHcJGZTr4KmK/sEvSi+a7y0moK50LywbPfK1F+kXy33VYG90oxVP8Jz30myorcT
N9u1YNgHvLMAtJ0IExH9cR4RJyWdLDMzVSs9BoQZr3fJ5Fe6RHv9HOJr3hREvvrZQC36pMjs3Bnn
w+YHhnTo+ybY9LoqJzdQTApEJaUlgt9XWQ5i26xQQZjj35P2ZVUzRNhTByQaeoDM5zNd5rcL6xhQ
yanUFZeZ55VCewTSopmAw4LTEfHhngY9Z5rsBptN8F4xxwWeAYAm6d6E4IAA4HRMMQvCe/YEOlWs
4lhiX7M0OJbbPjQaepwHijBmX2xRt1znRDzRJdh7TEACDWduHXxIZsMAHgJgKrsIzrGcljdN4DcV
OgN1PpTF/DomzPfBQjN34vqqsx2cTr6dIMg4dcRYVY0+2hKwqVNmPvi0DAZW9sB3ocbQotLO5DRm
UKH4zjP1NmYgEv4iRSb8rNpEx0ZHLOBuXBlAhB1qV6sAY+6fwWqNuRprveBTIgW2aYwR76Sc8jVm
grpXHAdbebR16jRya+RtqB1l7EA/QIxfp5lwpTfNj9+ey30ZxlRoHFeMBRUY30M6uhMwGInfaSXa
im/AMiETtASGTol11mO64wVxYvr7mSM37NfS7OzbvgSWpwrCZkO+yWxuLRaE5a0wSkBDL4jZbmo2
/3om/Vk3F837ERAVFjj0bxcbGoLan/p6vWlOHn3gi1nvJQob9bdzPmrd8ucDxdmWcN/+q9L68Rzz
B2kmt9HoxiDdJ6hVAkEotHZet/CSAblrqNVSthWHIVthSjnY0edkcNM6DJpC1hG/UMVt3ikXXnqx
YrMr/Ap5hzDpFMQ8HDv1fktYiQknvw27RIEKjmh/kAUzT4Pdmo1ZCrW4dhvExa+nmUSOlPKWWjf/
2QO0YYH+MlIYKY8igMa0g/SpCVt/vu7oblFwKYehWdmDjIVA21P3bRG1oCi2c9AJ6FPd9UP+zo06
hbMxkQjM6b83QHced7S9Qzu4plKhAxQxk5flxtMtzYeCzf0/YRiHvI7JK+//z8Krf101YLxLgyGl
XXbswMpweCNYsGraRq81M8SjKV4Ef6fmdR1ZHkwi7px68ER/ofhi6tPLFYNqdvNrL1Lnfagqjwi4
QJZg6wXNbsmiMgVK+RdgKY0NSLhlsjrX9dT9vq/X6V4I8nvceEHWlOdu9IUz72c9qJ+0rk7/sTX7
aiKFT78D+k2s/iOuPpPSpSl1vY55gA3MUC6TY2rGLMkZlQ7WksZto5f0U6Ho0t5tnOG7GLF/VQUn
0RGPv5TksIVx9AKg8OJI2zYOC3RwfMfz6GaYw+nDF/dV8MZrHhm7o2OEcXD0hjPSDdwG1j1+NDnF
EyVkMnKaAvjhVdcEksJSvoZQ1Sxup8du1x/6b04F1QWtw1i/M2dAkhZ8mTmCVT/wrwBYRWTm0sFa
Pke6eLC+bQwim+u507pCFRiC8DnMClACUBmZTiIGWG8STol8u7sPS23BXaQEIpm290AZJXu0+gTj
UmeuXMDeZUZQpnxdUFmcNp3JaBujvYBHSdeQ3P2X53rbbVG06jg5EF8ZkZiiptdH78Hnbwt/Ofrm
pzl4ZyI0XNntu6WvRkPe/SkehisoMhIR2gIDyPf9WU5imBr6eGsAAK1O3r0TbL0RATtkbc5HFDPV
XNZFTn3p2eehbfiegA/PHXJ+r8DaFUNtXN1CGlzuNawkYsVQYyhVKO1LI9C2M9jAETDlQSUQyRge
LSQukzdsLXavfkpkkMxpOWoA2oAch9pc1xtwSZm6g2ZGhGNoSJgrA9QldSDfIrD9HZXmSDJac7BW
DhMgeaYztF+epOXvrqaVFR9TAAy/yUxwZ4v+e74ox5uTzsOP9FPNKG1y3e/lD7p0LSgJ7DqMstxI
j3T5WbLVJfVyqayM3wSPQcTyPC4fIbMJw+DdbPNDt3LgbHtlnx9xCtOo7v/KZnVfDwUFwgmgscur
EUMC3mkQFo565ii1ulChDOeYLpSEtCGSeH6m9aZjD4V9Zetomgvli+JUq4wfb+aJkq072Icvqyla
02qenr7dM2BXAqqAZk/Ea5edctYYXnbsOw2TVgcRtiWhB0tiKUZnqvz7S/E6t7seiHqVgNXVjugu
5wNGbAOxWpfqWNX8O6qc1D310t3nNMEQ5QEv5oGSOXxbanbfmxyRvsjphMaNgrUOlmILbKCE8HM0
e3yvINuiK+DgSoJHF6VFA0uOy1u9Fy0Eczc02SyH+eY418EJTTSeA8fzACkyoSArHkjn8PjXTq7t
wYTfKqf2/RfH8GscEhAtg71+mjJ37y7gDRNpYYy7F/8E7+pNVsDEF93aNejMZNcrnZ8ka9fTC+T8
6xJ7pq4h8qEDP/wqdA8DjrwoCKd8Zm73GOnpEX1ezvG7ot43Q0uGIvW33yFmQuGuROX8zGRZHGvG
eXlHMHLuVtg9EKyMZ0JRcCWgBN0wPi3oHa7cN5XatQdDn920ess3UmVrM7E1Wx3didAJe1OKqrR0
XtTD4gQ4haL1bDbUhp5HW1P3wecYjP7cVVP3Z6K8ZRlySwtjTqU+lbtDPmvho+PGfwikOP0JnScc
OR94HDucdKuVQWzfWTcUeSgE03gtVfNgp8kA6hcFiQHPgibAq5wPwX7HjWVnVfUlHcYE04D8KECg
chygog62nzbIO8d/wLClH2NiyDWFbZDCdqbaPmbozAFZ+D8m6uuunrzvGptSt2R5jb2GRHpaEL//
k7K/fGf0PoYJUo9g70yBfD2LfYRDY5jXV1UKS9WzzMjKJN8Y5y8G2ggKuNzeqdiPT22DihjD9Ax0
Z/nNbS/o8QeOIjvlY4y3boUDmFt76Ne7IxHnLat9C1sFY8lOhXhZ6Hcqg/6WtzInipG81v3ygeKv
k1g7WxYx2D8vkr2+k3S3c9mYsM4bJEfErmHzuLmB9II2CF7flyboBx3ip5N0JjhO8E8tkDSWzLA/
eJLeUWnXJQ/kDCMW6gg/HOQK+ecHiOwYkf73XYoqdjnNSqinagqcnq4CL8waMyqoFLbu1ka+usXU
X8zMk/Pf37tJ4EW8WoVEGcrW7No8U0uPbz/wTWXZfvINQrBf3iu7iUgqhF3yJIWUSProR4UDn3+y
N8n2QC6efakVjmHRKzhX3Op87gN75xrAjFFLY1+OWXjkADR6MpT9iAFbWI2LRO9DzNPC/aJjeQgr
WuOjT09vJ1d729FymR+fVBFtvUbdEUqohKbm+orI88RCveoFFOMCm1kNMYbLIamY+yLkCBCwbOI+
pcEfcucYSoXwik7z1ag9fsR+uu1M5cq9nbqm0zqAevd4f8gTatr+VYFduWJwzRk/uaPRstZLz2kU
jDrUyYmwH/n2heBuwDSbkgIkYYxiRaPpW0K5EkxDAtHFzPDmhEFxfwYdj9S07YZDThEVD/K0BTak
cbr4lSwLDvSGH3LG0NMPC+gOW+MyJs9gzSilDvK9dsXUjRzqrPhnAo+QJd9GA6Yhkx7znR4512YW
ezUeSMXQVb4jg6siOO/TMOLS24WO7S7vStXsyQdyRR+DDYFjZYbZtIIG1xf/tXrVfZ6nkkwXy1sK
flcW18+kn+P0w5MvrEKJ914x2UX9QKum/c0XDJ6kMdMZEUrj6yt+VNaI4six0dLN0UPoJqUiaM9z
ZLnr7FaeyOELQUJSpMrjqaY8rxUiQShmZ3IyHU/Ws6yFqu/MDmnCc7JDloJeu3ECW/HA254LrwS+
40lWS3ChQyCSOxkq+ptqfjhAmqQhKg/qiUD0O3Zhq4Ej8Ub+99imp70USz8fHmGMkXWBbUrgPbI2
XS8S32q3cSOcpBVFOMw4MYAk77gXhQ35em/ennFx1lL5ykJSHnbAvIbIMjkw6NpieI+r3kLSC16x
bohAo6bfScCgfxUwinJcooSVlVCKldtLcPFZ+hJKMWbdHxhnmM6lJCDTN2NkLAZlGAELqd0Hz284
Vzh8/F0+4+jEDDJvwNJx5fYopujD+5FY2mDRhbp9PXmW7gU/+7vj+9w1fTtiA3qrzhK4zrvelGqB
JDyeZFu2a5q7lhK3QIEJBEbNAZ5LyCT/+U5IiChmZisyMdcmfzdOgZmz/+J96WMCV/7Bq6YNDvTc
/tZt10+fyS5/o66McmnIE8YRXF8ZaaLkDDXqde4Oz8uc/EIr6cxJlo+yzfpnZg6aNbA0k8JWPBZc
2/pafp+VR4ddkoLUJlKKr99LNv0GpPsH6sZ5QX0I2SS85cEDPM89Ho8wTFreMck+sbq8GKvYDuXR
DQs2NbdYH77ocFUHtpDeIqmdBHmkFad4ZoX5Z7nefLDRt6oJHCY2xwqVB5P3/zsOwrFmNXJbGFJ9
01o1Xj3ruvA8VSj77SedcYwXT8zbYc6LE+qRVYkwjZSEKjN6wExJ4+y8JFRRYqO2DaDRi0/E5kWi
Oxh9u9dUg+NXYrpXWZg+NwL3ISVYLCHvvooYNlIrEznPzM2DdsHNjHPh1SKUzLnasvJRT7esB/rl
E5jr9grfds164wIjJ5PAzeWDHQdLP3SFQGZlrk+sK0f2e9drRPyU91x0z+K2fA5nQdPpLqo6g3EV
JOan/TwaDeu8q/wHAhFnDky+XKgMbxQKsZ1LRWK43q4sz0gDwFTig3gFKZPgi7QCIEAE0gd6cjKZ
hF5aZKL5JN780KravDXPwiMl9k4ttAOjjXXPIh2NtjLCII/eexgTFYDVxyL40yy18Faz3d9gM4i1
AXM5Ixgf4dCVJFufouiE+qqagAuSaFOQ+xmUaYoTc1iptfVCq+wlJtg+WWRKczdUMp4Kz5uBi11z
SFwy5iE8KuGwbK4SxXH2itXr+BksjpCrTSDwVTzPpQIQTnMBVF3yKgnGdelwJs5LH2GLtR9mHG9S
Olb4AA/3fAggIoG184uO9oR9nkbnjzOQDF3Ipx8Nc+T9A0k1K/wIkLd2ur4pocfAYcjaWE5gRWZy
KTPzmPi28OwTSIgPn0LkM0nynivWuM6b0bDwWE9lHadMHPB6NcHzu9QbNVkjmoTWyogjg/cmtSgJ
OIEPS1Bj8kElZQKH6gT8MG52h7jj/8jLse0O9eYuC1Rm69hOIxLq3lc1a9xzwTdFzUwBkwc80ZM1
W5es53RdBC4xIc+bqh7KUUHBolXKRCEhUufYLdxETRzsZ3rAXygA/vXcyKLp3CSDdNlPRh0UVHok
pEudsnyRlIyGqpXf80BBTGalm0fzTtVTDv/wMs22Ofk3YDy8CXTNx+aZTChJYHfEZpZBByAAjqvW
Bzmzhu+2H6PcjTxUt9f7hVBhl1PvDCi0NTgk5FsMOHh/F/SDlJHL4Njz8I/JDZHOMhapw+Sa1/WZ
KkXmWEMlL6Yp8tDI8ZXCI7uiQTpELeHscXTtFUBdaFeYRCypa/LSGmZKDWA9ilnivbubIYNYanbg
wIZJ+1PWidIy90RDpyEPBJscFFvd0NpeSUWpMIh6AQbjVles3ugyOvT0oD1JHgOGWa+AmO2/+Oro
vyly3yCiccAZ7ji5PKhycJGdtFOmxI2CeaNN4+7+aAZFm40uqUhv5JcRd+OIoGsmUeh4nzBylgCE
zCiLWf8GpXVIHkjeDV5SWzTQ8GKCTQQsBfPbqWreuxfayjp22tV3eyuSBKc6K3X/9FEWxvdt4Mx8
7xHb0zQNjhdVc1Qn5i0zHZtghAqaSdpUPpIo9cPzptMlkfaF17SuBKZ30YhbjIJQ8ekhX1TDTAdJ
5lw7pRzhzauHvRxTVs7/V36wEBXrxBOFIH9KJ0/zriDZoCJU1+ryvb3q/n2+q289Vjv9EaNg2UkR
2lQjjyA5SDvB2hSsndS4XlbVYTFqgExLdL/zvFjINHwmgnZSIRgQKZsONX6KE1tMuRT6Day0u4Gb
/9cAw4IsCsUyG5Xz+x2aOQ325XnlR+t6koqCs3IzdFjdsVZtOf7yNn59GvfkCkk78QF2duIY8QQR
VY1YnHEwunv3Y5uKaF9iisS8sQNmRGdZ/CXVzHD1Gt+WvCimAMqjV6/nzG2PEXZOXdHcP9ZSeG+H
XZi7ioP0vbMLWTMUx9Jmf6qZ1UAla1Eu1mxNGY5Aq9vhTPAMOBd49H0ilknD99IFRGDicb2owaLi
j/De46RDl6KulfIRoVfojQUxqLol6O+py3BDnhEKyCAgi3oPoeOeP0BU+zG0qMnFuUCK0yMkks/p
gthhArEDdYQbirOgNfZ3HKh2NCvCQhhFsiDDqNkhHN/XiQHPncJfZ7y23w0qh6gVmI/3bJ28wc95
co/N1ZWA/BHG5DjWgYGdm1tU+3pxTA0a/dDQ6wMVFVP7wKmBcNN6QBQfZquntP0hp2J9hgDlEr00
43VupyX3UCyUqRhhNLyZUXIBRbepgZII39SFDmiWjtBNDkDY11BtVdVAf36SwEv5IyNb0Pb3Ps9N
c9Ohkt/TJEBwFJkWzvZQMEGIgr8oL1ptU8yA7U3LpRoAwDTTrg0/RF/9TQ7PxgbCYGcnzQJpk9x1
RYHQJ6qDQ6CE8f/RdhvKTN/+wcg2gHEmlWJwRdZ5cy24GEl8h2WlyOckDVmXMqT0+++xrrQvczlD
9kX+CexxXwwWU2DKerUCIy77lu/gglldENUu3/Q6knFEXSSKw8WvlsM3BDg5oOAY2D2fJYL47mKx
BGOIorpP9B/sLY6Pwy7Lwl9KJWUR9kezAGutC5ARjbno9wwjaCa23bWx8/8dAQimxcslx2v+FsVp
hzRPkMStKmJtaiehklmiooo8cMo6H1bvbmU4Bvh0DrqCcy9097yV0Wo3coTg2E2FRhtos2umEPv/
wSjusdt/85vSYnQlqsPSAtB5jq+lpCVxvlJVGBwO2rnF4CintUVsfA4lwuPbxuIm5iMkykgAZ5uv
O4XsdEv63TzdpWuoKuXf9Y+W8YIp9ppD1cFHacuN7N1V4TvOUSysSnRZfUtI6BCOitw9xfEkCSoU
uZ3ybczmI1N9mokRAjOD3mN8nugFIidQ+EcR5ZXsAWTcK7zTbCL5gYLFLZQaAiue2/e+oUmzJWRy
/xqfQPo3A47lkKTrsgwzaW2ZAz6zXFA8ArbNu0HDZAtyu3stLRrJq67ulbfvpv0gD2RiUI0p3tL8
8UXIu3XVLUHlJYHAsfOJHme1eTu+xwgNt13JZCScig560Y3XwPMYx3mzyBoHLCKhqHXivdrGM4C5
dxSWopnxlYR3AhaM5GKRlYY5h+ZmvtO3kuVgUtirSAwkhQ4sLGv8ebqUmWAp2Z3B9/XfDrt04Sjb
pjCb6wHS2/DeB1s2hzrPMmmwrCkrJj/+yrV2e+mRdW17VP0lbfZBDrdIlH7WN4JJlRqEkn1vTnd0
YSme8TxtJ6amcSzyZhC8UBaGajk1oWyqU6bbygUj9M5sCfZ8/fth8iKm20zECw9+o2t0JuU2Txab
dYDa6GySexs+SpE6NRXd18DhztOpxDnv7jIRQ6d/7sgSKKAk9nOU0IWlS2EbtKElp7pYgvCCaksH
uacRtZLfFMqTdVa0pfjVbUHbF+5HKmX5vq8nDWGf46VVqQqrv/bOY4NiFrFfmd1ASdU20ddLMJFk
+3yrwErm7gM8YEZLcMIbDlbufSrE7ish6q5lcXYNtHFlvQgkqLRtCYKSgASUDQZsOJF7s+DjdHGE
8ORobBCUFIZUOmHXmkhT2koQ2NZyimiPC3S/gSp0g4pEsNGhU9L2fuSndjLiWNOtWpqgyb0M/ZWh
Lx+NfMKTMxRvc1UuYAe0GIYAFgr1f8vWfwU4aRuYM4+KXlStcmtX4Kazpulw/W9oqy2MhHa5LdKa
JgWmqYXPu6pKdemCj2jriAv8nGsJICfqCy1EXV5l+2tDR7ToWBl/+a54RecItMOJ7yWolLbyJMD1
oKcknGCRMbCLcRNwzMHMqaRztM9hi/K6lf4M/c5GHfn9ng0Z9bhJY4zydWUHawo/erj228rdbK7o
Qn06FrMcNAEDJTVEpJG2WiZmBa1pMxV/YLMLkzbJZuD5MHBsc4Iz7hZr86c/TPyRgMisBB3xHeRC
cYLPSEbCRwwutyGcFdvfgPJYyuc/YtSp30xlduHj3JuBjaCP+P5/8v3knHQo/6OTAJwxTHiXIRX9
SI6n3M5yvzyATjU/EiIY8VMGf46y+4k+iLLI9Zf3waQg1dzi8Su8ILoBaF7ALDpJZIUvdHFzJ8T2
qOuLTGB8MMhNY/y7whLWhM7i8SOqDs+wOF5EC+OlxShEKIEWGEZYJ0JDhvQmxA6XeStMYYuWeo0C
+/w9kzT5oQPoxv5lpGqZi3VGFBoGA7uqBfdH0B8u+dP2HEMfHmYGA9gaajffI2OQG/pinmhOMjYw
tCoSFvFCNRjeWSSZf9uNXvW8UcX4Lm0LyNZCFJ8+Oy7oQZYDmaS7rpfpCcignDHnRcoJTJ1vrdCb
6DXYkdWWCrikvYbCG2cT1IElxrmWkxNX5obYnl+BC3oR+w8PFCpTOJE0zsMggDknrXqnX1tKXAyj
uTjEW+GdEg58oEBtcErjo7lEFXsU7tYe5CGlJWhrzaeC0Hed/qPM1azuzAilo9HZqPkmdz5KT2mb
7BpzHvpNctUmAwqpCP6lYGKtynxhevzgLJWZ3/ImZRG8zENROQQmIKk5DUgWykMIFP6YTF0tJzwW
i642rVO04pA9ZbfJraV4jw81MFanp4JVP5s7hXGu1LVQ4ZMKDrwAux+quCwZaekJp8KjY8Ts92G9
dfR/yd1ujf6REQPeOgu6datld4S8Rc4rTMaptOK1eGZvyNc+D5fayQ6tWnPzGT1ue3o8iX7MuVYK
QrR7k7PE/ayS3Xz/XANhhKC1avmqkf/OJuVjN0qSmZG4n6UN3DPeCOItGh5lXVoneTZKnQgvrNxD
eXC4LlmQotZxKIFI9U104vX8WlkCWr8G+LLXKg6Do95RnWHhYtRD9mnKr1CC7C46Nf3Gf4R/8iAW
OzbmBcs3Z9w0EFaIGsvcwiKoMLcADILvbMcnGGzkLWBBDZQ8HWI/pvYe82L9hqhu8hQ2Da9ODw8X
x8O5GfUX+2fVm83OYqtu7MG7EVBYcykzII19PKE1kE7jBer3JeJZ9lcvxePxDmxAYaMmJEzAFk+y
03UOPIzKqdsa9bGAbTfj3spaJqC+Xorlp/mGctZm4z4399e3jNZeXpTW30znezf4EVHpdKWQUbMm
wLL/ylwcqpOcLVSHxtX2ho727YxWb50uYcM5vQ+W3lRXAqfnB3o8UvJoidbszq5uZDjri16iFeEy
AOmtBSfjmMl45lqy2k118DgfSzVrJp16ZJrhMXA+mDI72j+7Z+wFmPzFAHVl2nH+V6n/Ie6vfTqA
21VIFFZAsOD5NN/+p7NgfOxj4ky5YWjr+rW9q+QJgEDkw3cPES8g/w0RMfimKVPJo6ILwpoT2PN/
0gg3TAGg2zUf3fdwYYdVcCnXzsvHD4rXnFhOZNbss+EgJ2Qo7supqYCflE764TBqqkclEUGNTk1m
+BTgBN2L/VD4oyZL1NRjo92gzXeu8d1x1La8AlNB4xOpRDqYJcV9C+oIRoq69bsFowiGdnBwmV0P
NuFK0ay7XhNDL63uzSSv+NzNI7CBZhxtxB2dg81C3bk3A9mxa5dTLGGlsjk9+kNfceQrDGVjqMI9
M1vODuZ+IfVBScp9Nfo6m2JPD6BzvP3SGxsaZCMba9WNNhakDrNDwnoYm25g+aBUb/DMy9hyRaUV
ifwSRQTq56jSx/KktEzbPdFS5QjMHoOMPFXy7x4NquzT4FtNgZwWeCarBPYU3Fe2+r3XaxvpNNX2
9SsFM2XWBowT9W6AIQDq2JZ8NhCwcAf1z2gtTriSU2gqSP6HFk78Lc0asXnSzpvETE9Kw7P7gyVW
tYvcs6l4a+9OAqbrCaLbbgrDQucip+u6fbaS4+21a5QlY1ozU9nzlUkWHMz396IsZkwqIrwhkTrg
o1Am8+ZPPypDStYEmhaF2HOm3WLf3pCG/C2TELRHjmOLKJ77XsMk3hJb1BKGDk8YvXqaZu0bUBXq
fvfzfbUXHDgUin1byosqwkcW0WjSx9EZqtBPptF2fpePrp5Qg+KdYwPg+vKIbtEmCl2y5huExeeU
uTeb645MYIGqUvZrjfDDUQ9ibXk8zg48MKT+TbF9HSp9RHgOEWCxEMsmH0Sq2Egzv5uLhjtig0qp
PwD8cG/BL6SmGhLyYoZrblmFv7Xkk8rzK3KWhthkcmjLy/hYPjAPF4bsKPpeZ+VJYaFYvzR3M24M
3WhRtSKdifHGWtVcu44tPyilH5T32XLVjyZgILDNMyQ1QT30CHjnnpcdAHmI+vWk3PThBln0u4Pz
i90Xi7BAhW9qJ5seb6KujEQlAx8nDynJgtZn/tMHFVBYLFvIkpRGvOtcQKg63xGCIo53jordf4Ib
K68BUSyW888aGZFfc2WijAjxguoPK8FQn3AK489q7Vqdpni1l3E7YbImz295n2TxaBh7b8aXzaql
JCF2EQUsTcU4aaH+8olqYUjAq/pQlcMgTb9PvsuU3e4NilL3JnKl30Z450KlYwT95KURi0C4oFv4
JnzE+QxfxZcuTw2bfdGNjLm+oHnEzFDppBsFmkPwOYaI7PeSU8ygQtoAXQR21hdat981Tc4T/b0v
+9ibQvmeI6YZmcZsHPwR8ieATstNhOE26HVXPYEJuFjSbrzU/GgXyYuB305JltRA2Bf8tNV2Ire1
NTt33Rs00AeQ7vD43heNtEmTXt7n+KcofAcKO23JbwL7hQByHYp3VOy1Zm+8wKZhjf28fmyrhrGB
sXzfPExYQvAUeeG2xSgYNqYOj0ObbQlka927vdkHvgncVrSsr+JK/wdgjXUW1KQnTuiQkrdlke44
O1v8z2ssug7oEv9S1qmhpGEx92/kwxioZbgfibeT/zcFk3WcUMH7ZFuLAuhAcRkBlZ4g7nwjS02V
NVOQcsdTRkyOaQsDdgAibXAhF0RqCxtI60jLXlre0UxYPM0y9Szyd88JivI8Yy8HxCDs07Bz4120
Xtq4mZ6jfHSelBilzVm7djBWWCEZKbjv/ivBPv6yxPIEW7cXZjFsehDLSXq7jYT5ztWcbWUdVJu5
hTK1pn/xRuFBnIad52RGJ/qaAqL9XS7OUumkvEDCbkRFSOkGUJfq3cvtE0wD+z8E1wcYfAiyorG/
TiDo7ldy0RKak+vE/av997aX7ZOHfVKDZoO/Ci7ANWoRfR9Ypv1SKR6wJMu3uQ/+7kJtnoihoqKi
tUFj0G+cV64rvr5jj6hKLtCfZf8j4n13r1CNyD9dc1/R6Cl6RIbHlZ2BW/0q6lOX8asEQuxr2+Ru
I+aEc10wXcDDpnpQ8/4FIjsb7qHkqByDZfq+SSOO7VvpzxhxRGaD6GCO5nl/Nm3Swe7vOE2oFE0D
KKwguugFAn2GfB3pvMsjj5kFZ1KcDMg+PIxdxVF6UrhzAwog9u4ziTKaftMO0xoxaW+mhC8rznUd
FxhtJuh0d91npI7mnIk8dt8GomPSaDUNV+Yk+2oj3Mtp7T41SOSE7gri7pyEcVY+zuXXnMnXeJgV
AUE8i4rCoptHVAOmtITjzQKUGVyoqQK7E1QWk53b8NlvVpuOLpTAMABmIdYanjTndIUVXGf+QJmY
7anJH7y1po4aWKxdDewm/n9C7r8RGPnVCxK9LibNFomriDPE4+ivi1lxdLnKmeApGDQ8yd1JM6zk
7BJugLzF8OM22mVlhKaneDKYyw7Hi2TFcsJpq/DXpWstIdi3b0bXHF9SPGNnd3aZeOUc+OMH0Z6g
cjV9TT2pUG/KYGX5JNKMHa0xPPZOiX7Qlnx0Fof5ZgfN3nxCApt4yt+wGVdI9tRyJJQxa0dYuAUr
WuysueeC5bT036wAwSTWDk8BbacXhddHXnqNbqh4dTDADrKG7fN2XWO9xCKq0pyi0IvXB2EUI/fU
uutj3N+SbZmGKV4Nq0XPdPrbG0BeHwg2D9SSatE6YgtZW88VQ1AoWhGChu1dhxCH6WJPUIfHc8P6
tXEoNVHdlPtE5HLgzfESg0S+EK9fcRayi+ZNwOIqgEF6RvOWx1qCmHbGy8Pz4EQS97TDrXiOYhNB
NJxK+fr09ka9NXq1LSP+k1AIJTTIHLTknMaB5rTtwqfAAjH1lYp4N+qXfPzwpKb8bgANT/hBXUMv
EHONTVq9SZc64UPr0n8UN2wY7+4bK+zwnvUyj0BepGwxafCJ7SEPnaqq0QX5T7n10ZlCalqcYdWb
Wqm+i2XtizVTjKrcNqBOMkH7xBmN/bLZH7luLnPTWjgobD5ik/WhlmjyOHlwDo/ero3X2VFx9L8h
CGEBM2UMpt2sfFfUW++9brLsWw2x4nQ6DQSa75QJ6RSdx/i3jC0q3aDOWg7aX3DYoWtLr9KmnSyP
QtdUaSpyiqVtixIbXbAUJAmVjw23WbERnE7Fd++GreNbDGswtZpSvk04Bns1wt2hPchflzL481om
SuONYEggo9J+rIDutbTEYFEQQPQlHY3kjUgb8gTmxMnXzDK6h2UR5AdzE7VxxtpmUS2mH++Ykayz
DyGR2ucpK+5HuEht+1Yjh9cJN5BA8KJ5JrvNtMIxmRiT/wXLL2FmkQG4nLbZQxDP19iX7RyUifya
wSMxbNepUajZDMqTiNkBmPZx6k65XRtk35GYascidT83q64yWLImXP2mtBXvFAeg1v2NemMXUVcs
97aAuSDp1SipqcVQeQ3/I35tTo4J7dHhpLeUh/tEpA7oUGuqIu9ky2H/sszWF46n8V0P/vz+Wii5
lX+C7Zdo04nVIGak0K5Ye8DP3bmkfHuQtoHWOhzXHrEbGPYxAGI9VaT8eKIXm4aamqXANjUr2NcC
kfBYsTRFIL6mlVasNf/ONGrDW0N2M5ZaqjRiYHpBjWAdXvcYttUZFNzk9h2sQRb0IVRD/DWeZ2Ib
DDtg7Up2m2I4pNkUeXBBgcpWX7X1mM/YE8sXpmphl90ulbLv14A4ITp1TzP9ddluMJm/nPxrD3Gs
vrk2P3mSnuYsji5I3iUka5Z1hIEXrOVlYwSyI76M9f/TR6tz7RxKK0DLDrIQSMiymjnlgFSvQ1w/
vUKOVGVH1zs3tq+FJCDmHX70NL6CS88MXDRou7XgFz3fn0F/7hv711L+WlYrWjgpxGhE8YzRQ8wk
/zL9bej0pHoK6479vViGvRVYUUAjKPxnXwDuBWxZr6ePRr3/LeCglJWWuIjhSn3wzErvRyI9jnBf
JbQl7yIiymnXSUGSJoon0vrBCZn0cgnYOHQ2EJmGhYdebLq0Xj2okBnA5xKdbgG0E3HSWWKQSt4m
ptahyN7KChiXOlp2+iR6reitmqef85olcFu618JJrXlt/AktIUAeHVAyNDdIJ3VYFOWYHk/n0+9p
PbDzGNLqLe1ZnlqaE1cgeQVOCt9MW3b3xhQY0AOnhdfOPmB9PsTkR27t7/16+stcCC359M6tgWQ9
p5hZwMp0jTimkWRoFZBJcodK4HdpPOfQ1E9uCjagoUoK/I7nGRK+KyVADzNXzZg/iYe1iXhzt9yb
OSSC7sGC3GxvJmVF8rDXRCnWSRmtEESIZl047GMJIhUIXgb2llcOQYpSct8koV4cUjcHTZnNQ/II
rOSQacb7PP+nCyCqcF/ilzgoaadifJz22WA5RjV8PQ3EOhYUtCgN33eA7naL83ZzlPeFjFfY/wET
GBOdtZesXDsOWoN1ko1QPTBC6vfFe6U6HHYJLClJ3DJIbLNxvoTVCsIv2b+vWAWPckhWimp6t40W
f1OhPl8au8imhi5tdooBffU0uOFsUd1gRPdIdBuALmRlHw+rDqBeyPCQHE4I03BXyhR2NNDJe9Yq
P3iw0x4Pr19iVhgrI4cBIRL88/XAekAn3FiYwJf+5dtsPgivQySDrbtSJVa1Mz/ZZ+3hRoBq1CZJ
jf2ZMbg2NQb9emxK8HM7MQeLOM8e3lA8d8bxKAQZaY2XOYPVrSNXy6CMbRC/n9Uk9ImGNGkXmDiy
T1ekiJQWju6+F0jhUb4SomIOKCAM/x3GnNVSuSrjSvUI7ilZZhKR9eJszwt03TLBOg6jhXf19nZd
lfmrlCH0hOww34Z7Iyvty/gbX2R1L38lHWPdsuJYseJmwTNJhK+oZ5NWssxNdJ3BIj40TJExftSf
ClTqaBco9YtOplyoXCb2JylRbKHBdzupbWGd7IlmUJ0M0hNeHlUzMYXPFJUoFE1YditvoenGmKkZ
asV4vNee33c49dg5t3MEHwFbPPSGBXdqKkmHpTzKMdDUFLWep0xr/miM43drmfcvbYtPo/NccXvb
ohTIst6fM0K8BrZk4iLmGoovktHzX18+ZmUMvFcTSEcSxB6k2SAtO+A0bW1b0oJ1KykZvIfAIcbJ
hihE/G1AlrN4UxgAnj0+bna757BB4Vm2u7wRtT/Zcz5QH1roFFMiP9HIho4WH3Cf7QBEEI4VYlpk
vaNFtwbwuE5mLni3SUdIkBrZl8dEXHFiSDIdwhWIqIw5IDvMIBz6ig4oKcLjOv6xsycfmUr9RaQt
rOkIisfcKqPbpsuibEEA5qkYllf84yi/8jBSRzx8/lvhIGfyK96zQAw01O4CTp7+VL2vR3ba7jf9
A9Qo8KYfKyfMoEYG5MVeV7swzl40EMbAdkG8wFYCiCkAZZw/3OfGJgOHZIAjLoZ2d0PvD/uwyz4O
5p/IS9T+Rn+Fwooh/00LxEKptyRsTrl73sQXrSiHCeLkejeu+J3sSPLfF9wdJAzC/u9zFhPpIqX4
VW9Vy3wKRMot90SAMa4AJaxEDBKYZkY1LDxNJpguoxs/eezEwZJgWMpJcVtrf1inBARdz6qVPejP
w7aeyL6qAEt5h0ssBRTe/NWf4mN7fgQyUCkhUdR2Ee76NLpuxNIqGYvaj0TcdoEaP9gDAaBlSTGZ
4mh63BLD8bCJLqv1VSul41zXIZTDJEQPVqGj+wJwS8O1clMhWZ5QGXsYvS0xJ8g1fjQZjPfNlyJS
UN1+JAn/Xm5E4JOnQrV6bpGRuHO6Ke3A2PttOG0zLTCdWONWlCIr7trwmcc/5xbvjBmo+VIFbree
bXITgxsQTgVsIKbry/tNCfDM7L/fl+tyLtVIlAJ9cqSE8F/hiqzCPkef+YgZIFWZevv6j1QBRiFK
pDkGCKUYbVkgx+mTcR4z3MFEobbehqk+DPbQhlTvj2Gn6ZoCDkPRVy69GUqWe9Uxec7W/O/CqDhl
w9NO/ou4woQt+JLjDBWeYYqWfuOgMntihkkYGbbVckEV7BM7rzekbR7YXuxFhJIiurNhMoOiOi1p
Cb5eP31QVnNHBY44G9RwnPBMnw6GfQw8gvNvxp25nwncPUTDMOWg1Q5PVA/FYeWm+WFqyorbuafk
rblydpcaz+kdVcMRMI3Lp8jD3G2aFllRXyVPFovyaOVfr0/UY64Ietef41xSbolj0pv9uhld4JZD
m/usledsEXhjkDapb2KlTRXsSCvjW3yf2i5wTobDxZkLxFM8KK9I/WScUVA2JJHCxB/z5kSobUlj
LrswMXD9829y9NzG/7ZtDGZZmD58bi8n6FjuZSYf+TLKBPVMMd3VNd3Q6sQVZFeguP/5C41+9DuH
eLr21yrGzACZUjszkhQl7xlxpCmEK/jEIkesqfbu+azg0SMGVxQcwAJJnkwdWHAKXAoiChxzQHYU
8W6KQEAkWdyo1U2pN6KaMYYf4Aaq7atAHLwjV7EBaj/lfeV9D/FNolwlsj6IDqqAp2j0VV6z6NDN
1FVNFIHdHp1DIk8OS06hCFOy30xvxXYPh7PRr3UmUr3lT2SR6VXr9KjJXGfEoqfeSWotiRHdks1J
W+d3eNJPRspS/25nPsPhQnz56S+ulH1HnV4pkjrehVBLj0e1Eq39Tqieq+vJokL7zIXXqkft6DL0
0EYxuuFhs+KoAML18FG+0rJsxFhK1trjUVgGLVmaRbz82y9UmZh0S6z/bNuhSCTCk+lcC/faeuMM
ukbzId9fu92/dTpeBqjmzbYhUJgsGmUnJuewACZVTt4dj7gFONv0WU6bQDRB+wIdyfusYFBMqtPC
zyv24cp7y8KdBnqLxzeGkda1M1XwOjoDy2QQHXD1O1WHEMPec+p2SWdhObhPtI/ITbDYoNwg8Z+Y
T7UZ29Fyx288pO0EoCe/SfyYj3hukYoJUXuRx6DPN3ZnOySA2n87Y647wLro8DW8lZTmzA0owFlA
oUp2WNX/UG9dKtzmI7GFknwJ87ch94WmYphUecte5589JUqd1yveR51ITmC9HKS06ibxWX+AF0yS
tvgiFgIH4IxU+w8+RFOjG3vVF1wEpFwHYqS8l3us7YSevb/uFZHZTUz8sgUG1Jqw9kqNnlOVD9Ia
Lkk5N8avW2ec7L6jN5Et/1Lq0MA6wdqYisJvFsbW4cQp4tgidgs5P/pZNyjn5aTezU03bw2qUMRV
sz3g3vm45/naOOaJYSmw4zJFvlJn+g8MOeF0zn72gg0UTEhyNS7Ae/lx6dYYdQqbsgx2nToXiJrS
0CayitZ62sSYEmur/VJQM0S5BW8vdbFTpzdScayvLMEZMzlu9Ua+xtY1KyO+SlA1YgbiEm3kqvul
CXfyARybgcREzMpXSmAMXyWJKVV+mcRysCK78gSzPc3Y8CPvrr3Q7zKsVQI6YEWeAcA1EY5GgMnW
IsTtL7a6Pe4Ap+EATDRm1MAKFHfJ3yv+Uh0ViMZv1ukAAt9vDTShTTDVioWrx2n7Y+5vSZb8MZh8
8GxZDOkBTVLrORf2gMuJJK5MxRdnECF6946xpFLTZncwAHvm7EdmzFAHnavH9Iw4aFNngbdUs+pN
qg95UP5iAwRUtRMpFxcWGuw+5Q9x6hp0pIuEWfHr6RoVdgPubhJVCSsy4yohZGwcfgA1VF9m/zGa
WIft1zCqjYXty4w1G+ZePt3MoV0SGoLZ28UAdTu1Kzpyca1WA8XPoRb/V5LRybaCcNc0tZ7EKdcK
3yhqJZFBAy+mQz3KLTGFm7oT4hQLFgEU7uTAYL5FcxIDGae3euPG2Dgw7AEZFkntaEUwhfLJJs2/
HkcZhgBGhERNP9IK0skinQVyMaC+928cg4JLy3YTQ49K2aY35ZWv4NNJkH+HayS6bDzd9szOs8/3
jxyXpTlLB4HIc2gHtPzWdj69lH/KPsJsO5xxNHUTuweZfpzW75Z58tzPqDGpyC/7r0eFUejwQ/Rm
+928ZceD7xhGwiZNe7lFAisB2ZzBmNIzZ4QvguPnyFc0cVM8qzjNdJliBD6QjBdI7C5WZatxlCdq
3ToXWn3IZj30epPjyGpIQKuBNvPRhrIAj765xZXjB1E8suIrbgpzKacxewHO0/q78A8orvvXJeLM
lIanO+VE6LsBk5BJcSrz85ianFoscL31IUv5sbTvzSzmaRoDp+FO8sDgqSijEiZcu/hfLq4Idlof
ocpw+qHLsFaY3gRA6CEoI4xX5wwtf6tBudgMxqta2MimuzE2eU89EEa0v/MP3jiiHyEJqlCjLkVC
SUH/djQFxncScTeSG26UE8JwmlwwooM+ZOgT+4BgqEwMdyM2t4A61lBddnGxMAvqvABAM6POcObf
2dQQPJ82gkO5lAwgT3lSynfon4ZPpbspvjVQ8MXaVrYFDoKKIHFfwj9/M8dyJUPysOxU1Ll1hZ+6
Yuzdh1tUnVEqQn3CTCfWm1GwzHzNPkdhme0tTR3ba128Nw9o3/GkI/6SIx+o/DYLKcCtX8pFZXZI
TIpcBm8gOVuXtQbSKkHAMpBZ+0FMA33eDS8EqiIX8YAnvGhF54FN7AiCrNBTWBxgL56CYMkPAevI
RdzSbFuryM3x0QlXdkSU3D+aY71QOOIyrxK1JZAydab0eFpRLmKsSbOu1NbgNfZdilmD1LEAEHj5
bKcvnZQsHo+77JPKtzlrgjW98qTZMjhun61eWHW2rHHDWVIZUWhHJ0Oq0F16t4zQfaQroj8OlKmD
zCxdG3QWxyBF9bgxcjSy/0FJZW9jiUzs3XdO0RiltKG9+RIB8xY6f2PwM6OWjSLC9ZpMlDV4s72E
6E5fKRtbwn/aVApiHCo8Pg8Ufa3Rgkcl1fA1dc+x2BjnG3CkdIiY9pkVTkIcSTBdm3YMw4FJQ4sd
70KU1Nz7Esej4td9hq3EBvvX/57e8KUgEAESDfiNZ0QVad/FyOcTcV33WrGKxd4JiBiJf/b81ELv
jgC5WlBEMMbKZVqAcwVch4qXzPJlfgb27QRafo652iQ3ORDtf3B530vuqYL0W49+KQbrEIOF6ejM
pzzUxkvXK8SmoPpM1KONM6mikH1hGgkm+JUdiMsOLfS0LtFulO7ZlgLV8KF4x0IkMhh+FVOlU8S3
SeVCkh/lYbvEU3oKBjrBF0CzXkfB+bnjk3+OEoBKmpCAAzMmsd3s3UmfOs/WKLBLTQpthXXvHlUF
m/HQ46roZs17T0adrdVMNG2lhmRy56EbmuJ5eHUUsgaLd2naikahXIv9JVvBkfQdm+6JQi8cDVLL
2cjBCSx78avM1XABFCfFx+sYDUGbWCkBI2naZvl90Wteai9K6xeOOdVb/ro5fLgauikhs/0A6GiS
JLWgXWBynkn1Qx1bVPMRnGEjB7h6ZcNTctCHZwhURCVA+zG/pJ5KVh6kbpkGqJGUUKk66RwP7PA8
y3Nn/9AZ6cY3KGOgXZyD8m8zep06wsf1oCPoeX9rFdV/nvxutp3xDlvCQ6dgDY6/+frtRIEbJbtV
9efC2AlXdfuZeJb66ElAcNfO4s99kCE1wjVxqvWJFkZp9FWft+HIWxxpl+AxTYF7To3/nrL0hHf6
6um9Ii5xecUg0Nr0Aos7m3m0DESK3oMdPD035LaJUuQOaeBcXAhxiq0Jn0hhjB2Y8KK4sFA84WKz
iETGc1J0aQ6U5RWoeA8HPYrF/AUsh97TEGaKPtxOQ4NN7R4ZrmW72DtOtzyiPAf3MNsCQeCnTG2a
kRlnz6nDNIJsxjzV0yxBGJvKfYjWp1KDYO45kfc59v3h53biWW4hhILcnlCCcPxNAo1BT7ctYSQv
pm6Q2b9Jo8Y8jZEoTJVChA/O5lIMwybWs0SHPdD2YJ6JQiErbl64uCXPjtL0Cw9C/XuSx6Yjfy6Z
MZ3QxhRixlGzxusKCAyGFh6NaeFvwmEsnbWEez8tOJ7GrkvtQKjS266q6mC60t5dPDYjGT047Zq/
1QK0mElbhwL8SyTohXnoA4E7kGIdfGrMH18zscbw/2VxpD9gR/JAM24vsfZZ2ybQGkbo0H+fM7IY
C2bGp36HJOLUQDVHBQf7spmXEM5LNK2/fN09XIgePklnHa+nEes62WMA2YkHRxBpMIjnkEWyaMMV
lJZzRn3tT1Pjo1xgefW9oYXfXUdWdbe2itmudNyTFkDaMWkhNRGwPSHRDTKovxHZ5OsQ50z3ndkV
2vBhU3jsD6MoKCGMLmsNPrXdhBkOehSBmh/dO6S515jj9sGXyI7rR1gfbG6j//YOl16GAu36nWAo
nGcgctTS4sPpaIQX91a/HcxTX7eOzvVwWOHVJXxvTkL8hFkwnvSab8tzZT64aStEqWir06ZtgdF9
M0+yvJ2fBP1IfB3NgkYcl8E6mBVFL8KyFCfiSm+A+XcOB2PWN0cfGfDkTmBsQuu79ZucRTadwMJm
Tl93lPAUzi9kMEMdTffK5tZjpiSobyD/vf1Uxv9j5/+Iij9lz4Ww2jiUQGvrMcg1JJnI43cxnSad
RdgMJtGr0uIIiS8vr0Ot5kA58hQOsI8P3dBojW9IaiOWUxCUzdzk7rUUvwtjaL2glKouvRAHTMvg
nxp4PSo+l1mteTAqFKZD8b4oMQl6P/TAsQQB6dyZ7kkaYP6YAv6ffklgD9K2vZI00VJ4EOnw8ulU
t/wZb178qmhfS+iz1EX5Oouf5uUdotRB79yt/ds5sVnka2qN5s+8T9vSW1c39z45iSTE8zWWzxf1
JvGQ5GJnys0j3izrZRPlU8dubbThcwaE4nY4FdgTUbHzbnf//IxLX5nYZaQQCkzPSHK8QAI1WxJQ
jM/sCjyjuAVWcxkVDfIerWMj5pqGKuJjbQBEzJy51DRC6sgoGvXELAfYWfW2feZGdiVFXBHfGvii
79qhTG+ahWEpOfk5KDfEibVGUac1WyB/fT2pDAt9jfjcByLcqu70hryZ/exM//WyQoPTKTQf62U2
seFco12Hh+4lsTG5IRGOhtDT33X6la1zQDiXUSDSvozxZqmhOquBoi9eXo2DcREhG7niq2wgXcL0
CzSBUNgM9OL3CKVccxOgDTvkdvwYDkcE7u2rUQow2XAmTfS/IfNsFmwHYC/DfPdKRsaaeGXVyhK4
97X0517OhplQ1JL0PgNxDr74Sei7fs9n7IKKotC8dUcwkYczvIufs/Rmh2X4v5fvYGw4i778M0rU
YQqzQNuRLUyg02Aj2bX26L0EC8VxFwmJl1kOIEvMHXXPbkSYOZDT481Ej4TGAtdd/i9JrnrnvhIq
rtbpsQW/Spaoqr6frRg3Xc2uZoytFfnwFaNCznZrILYYIlQvDbQVbDirfc+MchdHJcmCtOvMRslb
TGQ8mk3SZdfkKeDOHsxLaHlTQf4ZtpR28KeXI2X7mYBj59XxADb5oiWejQO7Rpxm+4okX/dNtG7r
Q1zknHsDq56iJhxHOF5kG0ZNDbD/RuuDlPVCCvjjSva5restSG/lWOzNPmJYLnDqZ83TZoACjYV1
zTb/ANfpdkcxVZPRqlCucKALBx0pRrTj2PhcpbtpGHdkPsde1O0h/MRe2ARhjVgz8TaisADDNHh3
bRGf2pJafTv4F1Bt6IrefKYraky+0SKg+C/BK/IFJiBvQbSZu6gkmpbieKA48ofavXJG+jFMgSky
V7O7dQ2EcNOpYxiPLWXOyl24iu+bWxsu0rAu+cX9AiJQA8cFqTfnoUupJ4IiYsc6nIJ5Afg550Hn
HZlWxRwBZvXB4m44uhIqynbz3rv9DhZhMxxhihCcj8I4fq2MMeasnLAtRMoJnzSYVr1577ZxjMQk
KmUdIMJIsajemfs5Kd+yfl9tQm5JLQFEo1xijBy3pULsvCn9+logFo5Q/cCcX3FnZFCI3P4XD4jt
0vladOrw9iheYSvI02eFDlkzoURitnOdYAqyBdUSNXj4EyZlJJjJVJJa/Ep067KK3lNfRo3Jq42f
6C62xcL+Ew3SZUbho66LQ9i3yISUeiPNCZdgvignji73GMT1kkeMh1AnAzqN9FxkTveoSkmfRBTs
fhvsa2didLsZ9pAwOicppq4/t0vdlYYv8Q1nA9uBVoX0Zz+Sm7U+0J3Ds3qya5ml2tJjLxDU71eq
72wq7M8HQ9cRymLXhMDsGKQZSSgRekxslMIsMuYtA1RdStAZeg98l0lPXuRy4WTt3qNOAHXkm0Gl
I6++fixNH/R+efklUmm0xpFQnP6hlgbrTiyjGW9bbMPl5KNdUYkIhgh6CPxCRaHvN0uyTknP2C6K
EWCaJBntunpzgzIiWNGDR8uidc/z+txvjZxQ/kCPm4tf0Asymp7GNWH4k/VZpLzIE9WOiJAeei6R
7PeWW5pVNPbcTdCLxAcOgp0uoBEJt3FhAg7eMwEj30ctTh4ak74J/JBdyEO/JNPXO0/8g5LKM+oc
Agr7rpCAzl5kryn5LrGnN4+QKlOFWABjuq3Bqq5C8qrHt7wJ6s3A6ouGTnBEjeyExES4JXqLuS2D
Fh6veLGSVl0L8RhygC1W4+PqFD6idHU61mz4Nebyi6WUl2n679sjIGUdR+ZyZGi4+cWdGptYQzdy
CTGErokgguFnbonwzk6A1Ek2c1pzFq0WElAI/y5TgPcVGUXcjOnRI203fQ1W36gDmX8PXzY4cg2i
7qZ2qKBiC1JqlJb/6TkrDBDBLll2NE7Ycrod9jfKjeq9XfsMjw9iBiwcHJ13WT67Z4XH+Ko9hIN1
vHB76Udoym57CiUQ3zrTgPOOalRKEFUheJhyB3REEzanXkmmEhPVOw4h4hMpeET/uQkZR+dCaDI8
dQH99oVYPGFVeOdsVFPVnJWKvZ42JVR+BJcWprEGI34Vuw7WyH6jVKtNyAQKDR/KQx4Ob1FxMR6r
hQAJK6fKAmkacfA29dCnRpx3+GwvtIDbGp+Gx/RFbmzD1TYGjTeKxWs5wwbJIvxHPpUPA+72Q69Z
ldPcHDlYUHt75Flavw9QBKobF/QODOinhziioLSTIT1MZGw43UhG99eHcFc1jrdPRqm4OF6wbc5+
LVNBIGKVVais7X8yrNxPoI6D1YkgjongfZ+emxkxeIe5KqWVw2h8Sqb43bkV54oHTIVDhoGOCIiP
nuv5WYLasVm6H9C4iTNHgBsjCF/w9DZjC5J1ETvZ3csyPBwiItu2Z/BREGf+PRCdM67mfBnaMeQO
NPC2Rgb2X5aPYLHYhMwhgEYj/dLokpjVTmyBTc/SHsTWkQWNRK8tJGxXUmlZPpMwW2Hrrl6kv5ZC
oNhN+UZ+kxJ3nshJ15ongFlNC+0d6e1BR300yOsVkhyPFAazogj6a/ku/xGUiFNK8N8Cj7lYecdk
1dBk3Skv8uK/OTWx2K3c7X1CQMvgYoSEH8GDpMONu1C5VrWR1EFkuQtg+4TlWIdCFyhgMH7jHCQy
LHNzhMaBvZtDHa2urhZPzGimFxq4gFDDJhVoAF7oiQJM3U/n7AwVIpFdrnsVLG9y+95ZjdKQuDVB
o6jTA7BXvTMeNpEaauVqa+Ol14DvZLwmTUguwWQ4czU9CQrYHw3lX2mfHyXbXMHXZjgmK0olvmjn
ukMRi6h1BSJY9q4IRjYUA8nIpfqs25vaWS+cn5oG+Z9dyxdw7wANAkfomIyQy+2qn1hMslsrj8vV
ai9YAOrmQqjd4MTvJjA63XdktL5BkIFOJ4YaVUS9mX9StcMkKyYWPo2iVmpAIu0pG2HtA84jkwGA
pvXWWusPQTBNIfcm+CQwWpKKH6oc5NvULavFfooyijhCuQC54RhgFAzxb5gZesLvHgzE//gg3ny3
LQ03B2+xZCJ5pBDeIiGvKpAb90xC1t/y4Nmyg1iFO6iOFegg+KoXXxF1XBLA+zJLpSRzVy56zHXP
kpGL+mO6z9/ruUSybxmXCTNQSVpLnRckf+gwK1it1Hkov09Nzi4ZSdzEAeTLD0vG1j4JriK632Ub
QGLulHMEqmOYFSDcCcASCZuKFm6s+/WZRnvUGKWeipmlBE73IZrZ6CXpkwb2glAb5ThAdcmKNzaC
tSFoWCWdqElFgA4oW+KnsRVLHXz2pjhSytgEZgYJpgjbf5Y37T2JCOze2lfSzXMjMlkkOjszQ9Bk
6Na0k9f1WP6IRmmXIsQsG1sEic+nTLN373KEa9pixEuBhSnu5rtWw7e6XqXJ46rC1tN8m58DlYiG
a2SO/FW8Qs5XIA8U692TMKOS+0gHjWgDyKSHdczZBjbg44ZJV61no/Fv4oLGi3bnNVuE4Kkbm0aQ
6EV7IxX8TCsq1Wt4zFMj8KIkdBzgBOUsxPTulFuJXRWVDsYC9YJGQ6qXclUJHoq2LyPKt9TN+mTX
HVc1k1Qv0Kt19EvAc1UNNbt8C2qXehJrB7BoJc24RfMHiaE2T3ORORKC0j+PcAzNzQUW4yX/L+fy
SNAMg2J/Z5HnqA/+gS5v6JbXDWo7wLMgh+DHQV0LXMKhXZ1uJ6LwDu4gHhQ7UvsAEMvNNnmqmWNB
2DpUH/y5XPkqxGQYUCwRPQqf6loNIZmnN1qUMDXI/Q574ZNtPFXfAdoZKz59C8+MLAWLX6ls9j1a
hrcc4CUgSE3k81LHf3eHSf7BvkpE+u2i4DCecnNy86W+IUMOgIN4bwcKLTPDU66HAwUfzS1VyNCc
r2Ysz51kJcpas6iQA23snKRRBVXdGGApdQFr4K7fvCuKS8wbQEopqlaJI5kPArrlk+F1JTvAJqrg
jmI/TdkzItPgYCFaa9FapVW9LSWtIEcFf5EruSxnt1XLzlCZZmv+WH/e8xwpCVHIG9+HhpFWngjS
+MkBk62uou0IKoDmbySQTbJzbQhH09jyp/locUHzyWQECWvffjZcfUULPJa5iUpMEX2UmoSkzI5J
+sHjlT8Pa3PmihCmOAZFd1l65NHEI1RqFU00KQjaSDSRRQNZuxLrwVIybNf2DuolF/n84pW/7pan
JDtujsHJGOipSNdEqgrb90lDHFrwlY2CeMiiN99fXnJ74Rzv107CMVyPuLZX73tLk8NtOv462kfz
+EkkRuVXi6PD5V191ICiFsgvcteeax/Mitz4g19KjdIXO/PqnUFXyxNTAI+j8h+yj1GKCRpX4nsN
MxRImiq3Af3RVC/vQwdRUDBAdIMaqouRFuQTd8uSEhsz7gACicoztw48hH0PH2yTV6ZaEWThFzI9
xM4xsZ3fZyMt9SVpyMomIF9/zBXWr9tWngsNymSJ/nODbby6tai+EZ4qS580fpoKx0p0GMf80T0t
BdCbcU0etxcBBV+9ZHYnLuAqu/LzS73HNzVujwqP0+SZ79XOgOMPiV9PgbFLercUCGT+JWyUFIh/
/G42LSYYtZ68M3ELvoqf3BlttJxfi3VJEEhWeiYLKYeRbZmDIipFdqpqEqF7K9WoLo+fX6GBy1hG
oZ4PbiW3IDBkr0HVjujXNntLdcf82S+jiVgnBcCFbpVbiGcI/xa+asN6z+xwhY+uiUOaIfseYfAc
dVcxgd4UCCERSLqt6IY2/DvxtTQsw5nYsqv5KMDPbKgNh1VSXH7uy+3JOcN31XCNEEk5LuFh8LMx
tN1Ytf4/p4HN/D1M+2+2buubGH2GOQHlTgTGV4IEfzu1i1+KskGzVCsIFtpn7AnjTT/PQ7MMOAND
kEu2ZthntW1wqkrNNvjcFh1/D+Kb0WUruza5Rqcf5wDK89gAnDi8/fkFtR57qlKEI6sf9yaGYZ7M
tkvjzsmZ7bkA6Jicd2nXOs3Axn5NKbq+0CjqwEsup6gvV7oS3epTDME4TDzONsfl9Dfnnqr/b1kw
3QoTRdMxa3nTui6q4VAYbhm64eapR+dT2SYolvgu3RoWVzp2abnFSE261xOLIDfP52HFA3Zw02vW
fJOaNBD4XsCL3p073H8hNDt4c88v6KeGeO77230KVc3zVTskgr/zZzboyk9Xu1X+lKWY4cxIRznB
tsWAfbsZjhzvW67hZkFnHEp99S3dfT/qLSkzgRtjYKiqCYHdvKuc7C8j0FjDzNCebp2h1eK8wZwK
87f3NCyL3wTL7SkpeIXFz6BzmnXVclI9q3RlikDPQzzsSWpbFTxLAsJnA5AIUHQlE77GT+xtnRVG
Jeb6sqJu4/xWACzZuRUiVqZs4j/9e610EWRmxoCQVVm/Ky7WnoJkfQ2F61mTditypNn2+gqZwiUM
k/Em9uKu3l2rOqbJ3tScqvbEbvF3QK9eyyyBptbsPOaa5OL4BW3ztAoFdzuP9B6fzvvnlHfAdFwg
8mtZrKZr+MmPLZWK3+3WYaLjCSZB37X0tL7qMX3j88ufinXun8uldC/b8fLFzqSDRKfvgpnHGfai
I2lM7ztwYO3dOdiViHo8GgPFJHcV8n83Y74scKjVh4IbonRNHBJBXZL/DZiwXirqF6jRa7NYoom0
fQVZF7qe1a70gEzfZhi2ETsosN8Me2oCWrM82BYWA7x0WSOPs3iq5jcoSFYkpUAoowZuaEnFiVvI
taAQKBC7XuMORbyvkzzxuRwOraKv4j8yPah5aRqzOpTMF6nnHA7cbvhFRBO3SX3of8lu77mBNajm
pNs0BaVuS3eDDoH5q0ZJCjJuASIRpE9uARsI6Tf+B+CXMJVEgOCQcaLGTwUS6L2niqmbncMgjvxF
82LqzheuX4pdmc87YgRQccMclOt0rbWcA/x/g2p2ymU+HBDFWQ5+F35JNc1kMrXaVffQa33FYtXW
AzZRSIABDM17FxmNVdiZuF/77A6jMdU9PWwmp3nmyDRFYS/eZtyqLtZLF5DPxq2SDI25ZpArnKhT
DQLd3gsrp2YIO2WxWCTrtDtE0mK/k5ar4qTJ37ZkFs08QLpYDSc4iihwVDqrnVA7zeUMseuUsi+x
aZZO0FRz3cQDqw0nGI99AQOEjiwC0jrIKrY5ofhuBZI1mIv+bio18Uf/RqnbUJwzp6yk+EexE8mw
LFH7kChUB8r2bnMjqHbEsbawtJr8pm1nOOimyJKB9sxyGnbeA2BtyxB/oov3xnx6nvMSpOrqcVwJ
bRFr8nEf4IQB62QdzvqTjPqY3HaJRt+64maTgdcQNq5iQryhE1DpGikyuo2CbgJKJ3UUtRH9rxgr
Q0QRW6ljY0x9w42vNvVPlc7lsEqU3xAZNOAmnxfbW3VlxiOut5La+31GZlLiEtjYX5ME6giYzc8p
/WPGS+yyybwlJVwKf5fLCIM18r9GcwSfQl0EAuqJn5SEm7cQWDdbnSl6W2xDDlA2Ko7p+VsCfpfc
JAFz+i1uiHWAhtwN09b2JI5HmjNSGK/GJdoJNg2UQZolwvPtwxS1fyrUdcAPbBMGwznpV1H6NrIe
LxzVip7yUrrqPbFSRl4/omEHHTvVE1M/XLpzvjHGhUc0R0mW9oWA4qOjbg4n0GktRfqueS/lh7hR
UFxEvujca+qJbYv/zHU5hof1kbHuEEZxJbVxx96TLGsfpSkOU0tiF9nYNFIg0DpeRw9IoeyEPrtd
dZweyXzgqvZ96a3ipt6HREMpjcY5Wz+uMGanFEZpk5yOFGIc3HCLCTHagakL+vBVTcBbfUtTh3Zu
lNkicwXJuC3r4K2pgjeYx/Oq9S59Jh58zCbWDmit9Zt7tc9N+PYanDPFy+CtAO3Q9yFedNscEurM
+hrzeL1T2myEfCFLOZbdF6+Dl6J53E+dgNym8ZimMXbI2sAxfu/XlMLPlCuvGV2WUo9o26iB+eMc
ttMPdzuTDWbvMBbQ3YzhlnQmC2cacncB1wG9QZfY/vFsOIVvMUmTpbTZ2z+ROskJxRWfJsmxiCi4
AYAW5neIMIlOmUdsRRhF3khFtAkRC2T78JMGDnXyNztEI6hCKzROKoN6tDwCx76+31e6v8DH20Rq
u0V4InmWfTTyKEHCafKtL7syUEdFxjFpGaHnSCjN3Z0SpDxblidaEmg0HCZ+e0EmG7vGFBP5JFkI
GhtFc37bVugjFhlgrctwyPloUjf2LTlex11yvQWq6hkEwAJlwFMx9JEUoIfDXfo3igCo/tcIPMk6
0fmCpogyDYq+nl7DKUJLwf5XRS728iSsnjb8BJzjX1n1iBbSl2XzO00wHkAm1s/TjDSL3pUZSB7C
BIU/ZgLGCJ8Ocj0kVLqjZwAWBDZmY71RlTvCCd2BDr9DTM5G6Wh1iAZIEq4aKLKjWLrx3rS+9IFI
HQcVyVr3XSW7pjvCQaIZZjWbge4TMEJu3i4BN4BQvrPDPsY9p9gJPMsYV85yDuqjxF9idJVkwAnr
wMLomcqoFHpm2c2lstsBII+N+d1qoguxJJt5nwkBDZv+jsjnRwt03iBotP1ZqO7a19jQO9K1f/Ck
Xrzk5c7QO8q3Y50cMlnHWt7cAZ1oLBwIUJ4l5RrBBjyarFRdMhcJ6muy107is5dNilmrTTBAcFHn
83h9b5V3gOdpOY9grAD4EoiloQL+/t8m0c2GKokyfVASZ6EBjf1rBFhhWoBQawc7fihnzKOD41pJ
QOLFA0Q3n58awezUJ+hlCJstHLk+xkm6jP+NKvBiKX/GRvGmPCIFJqguJML860GXEpqQ/nwZIXJB
6O2CGDI3JeR8CFja85TEqq8L8fC0/fJWNJZ4AQEYXhYiN38zEvDjcJcGAHj4VCKMQj+PFc7J0JHB
PvMYreISOOLLYOfjNtIifHEKjKeEmoqCnLCrRRTH+ngQFwq2mm0nfxGU6Nmw1dWIA/JKwHMJoc/f
UHpwwv3NCdkGjyqbfyFpoGRhPFVw1MVlClOszst2IBhCWJ0uZL/omdyV0sVLG2/0LKILCkMs+nSZ
yLUo79TWqzKIZ3BmVdWLQMnxLnPqWTd1/VlrqAZGisebbfiSaCNmT6bIX++oGcIzhVa0VAZ+q1kq
iHphHgT34vc6hMXfrc+Xz53335uUMrgpV3co1oZ6pkKNx278Ejue61MelmeZix0f2+tINWDczZsS
4sFCcLJX3mErIVBKS/JTZn92nWVueZ4P5J/UPVOooTn9+s4mSUxjl0hFvEkJ8FWLWLuPgJI94ZtI
RdvnGA7IOsljbNV8Ot7/FLlBie2f5ydb2pZoo90sgQDoAz4lyQLtGpW4qhYmULW7QJAYELTfzHlW
fr/ULQBYqgtmr/87InpmUaBNvG9VSK2fU3Pdgv2cGYp5s4zwbsECaDKEIzi7SEnz+6cozj4cxN7H
jhCamwKjiZNH/f9+SCtVk7srT35FacwVOXZm0GFUxj07sNdv53e2omWlvhEzBPegC16580w4Pcu0
8zMVIvxBGlR5pVgh668mo7930pJLeIUAC5M9WouXoQi5ROO7Yyy4UzNUkvImcy+e9dFUqM7On4AN
BHLNqgbMq8ZXWni0tYQE3vVI3uWA2rskNY8SAeeZf9/GtWH5cRXzPz7hIeur6eI+ET7LIjxxSzEE
UgbJ17i1Cuz/Yj6n2DGJ2fv4eWSey2TYUgEezUaCB0cQLmYJaqzQMg5xXiUq+MNRtTkHTsVi2eR8
u/yYHYRtgMhqom7BXoDWGgp4wnLgUHEybNj7C4kDFcVyx0LpzygaOlX1OwXdChPIvGP1rXLz7mP+
34NTlnFI6q3iWXi0hCFftWBZusmxYQPOkxM8xaPI1zgtyTItYYC7m+oqO9v6/rSiUjkEDig2uoyW
3US0KOhV6DI7g8G1FUzHSIdweAMWBxu8qXMQxxstX7RL14Jgl5X8QLD4XimsUnAZGBO5NZlUhkvm
3tnGmDB+t5B0GvqTR72nWXiWQ0oWss6QQMABiFbNnOBev8meLMs/lelwE5BXX19/sQq1tAx25Xsq
UfEH4Q1kKnD2s3BO4gc9V5dKPaimV6RCu6dsDPR45612Ap++TWAhsqWaxEmJklkkcZ4vWfoKSDj6
o/HUeUc07kGGbZfl7mitjWkizNDZHgtdvKKb22IqkvRIn+gx9DrozRax5/+MhHngDc5rFYu+m7tq
mVW2lKzzLjJ+exfQLnAwCCaWJhDJMsCcPLzShJ8QB4zEXWcykGQMqm5jBoIOSkcrEkFy69UwNIkv
0+WcKgBEhBkqD1TP3fcVvUp8SSnKT0YdsTWvvFZKIrbD0q6XbK4Z4LvkIQbh9tfRz7h2SFfzQ/UE
aBuBKvEhEYfz9vcSjurtxovZI9roNreVBHn5IqSddGh0hTlbPLpy0mTppo0uyTm2hvtrCku/9wz9
tgvLv+lsnizLIT6xdgdsuQ48fPrzGyDyqt2eaRHeXUJBaNzsPOLyapNiI1BzXZ2J2rlElTossX4t
ihpEV5DuK8lHnBxe+7le7UOa9G8WrPdgiLp8pJJfWz2pvN40GCX64PTERrSpZl+nlwXrCCMPoCSr
LFrhdXnNawmQ6w3Vk0FJo8FM+BOWBt1h9VBimj2J91V49gognCfMwdAVDMJS6AOIOGeb6LBO8xtF
GUZmZVrPDnlTGU2KgsntmMFw+ITV8JCpAnXPH4CQMOxnynUTaWE8usPbFg56r5AU2K2lOidN1Sqo
eatTLD6rVe2JD7rIOSKxMEhEwculqw/QpKahurgHtskpEwi0+yP+JrNQAH5Eo36wL5nkyBWGdCI/
DmVySCgz0aFzgW0y1FdFOP103fov74AFeo+11VLh+7Yb9OF25lZkFAo3/X4ie8qVrTu/59xLjbhf
ALV5PSJCNXBcOCQwzh3zwYngBCRAbmvhFdAeqBi/bSrU32n9PJ7nb0qV2FXVQEbBgNJN8GPvZ8NW
bWRBkkhDYlSKgOagqg8eLoAEaGWuwX0TEbGhOMFlcJQ/uGHBPf1zUimTItEvb4imE0EVrU4WY9lt
T7LM1ZAKMXKvXtZSgfaIijJphSSW3TSRDfJ5ncTvrfY9mOZoCeUq+icxr94jKn5zhUwbyc5ahCgJ
gTHaEizL/nkWEqor3862rOdwuSWR/Qj6XS0L5EDfxzcbv30VYJh929+rCYLxGctdEHfdYsUmrp8w
wXfuguHbBQ+vxUMBjGKEY4Mv1v0emFNMom6e+Ziba6LJuWHU4px8rhf95jtJiPPODmekK9Ti7Mlm
WbRiiLDdz1Bn+z6JvpKatIFAtX/lH1WLmrkwlt2O7KbvWuR8eJN8Nzc8fU7spqGynW2Dub+RHRaZ
OQZykIjI0+cE+0CYtX1LgVLBFdH8J9WCiFTzuNY7+HbzQ0jdOR7LmMM8DSf4VaFPRcf/aABV+LFk
6CY9zlpPSVzEVsrzdwdalNGcx4Sw0UzuUyx4NJkOuMMziTp9VUV5CeMCrIgMY6hGwaRbUIOI9wo0
bhSrPMEwTbREd8Eqkw79KexzD3LSMjJBku1sm5TbUJfOX8nSOp6BTia/9ZSoNSb9PuBuBzoyQEd2
ioLRuCZIsz8HHpKtKyblM+UABeoJD5KFXUi1zV/4FpthkPS9F9KsTxrGSLbA6u/2yvI8lpHt5d6L
kEe2koUXW2UNSh82ZIY3MuFFA6CVBlwPKy4Ng75NClDVCSsuGUU1hb/xzyGFa2heuPRjzCKSuZYB
KftaUysVEJOG55B5VX1HzDdw2gAH2ZIb1M9efX4zKziT7Z0NqsJEwAPNwc43Y7BFCExjYv0Zk76v
f63uN6dPUxuwMLZO/ORRIxqmE40OFACS4oNH6oTQU1G6D43beUkGSTfOrAFe6uh9ne5CzrRjwWmQ
HFR/SaeWEAVNG90uLQ0vdp/Mpr9QW7P22J7CdlSg3mqbZQSSqGmipHopkhgLGYmfnveAdcEYr3M+
F5loO7orwY4Qt+JhNHulOt9yovDYdnXEY9P5g2FxWQ77RvRmDmFOaWMlmP9GDtBeiKI6xr+/EBFC
qQClt+lhgc4xx/gLtQCGbw3+VkgJ8hNZRIneLoFCrP0PO/ReTZA7nVZjrTen/xKd+i6G/fU+U9Wt
wz+TAh3jFL08iB5l+eMl6WaH/Vz60f6HL4n6RoaSOm1iwCfq1JxPpkSVPKbqJE5bMGS3Cef8VN/3
TTm3n4Fewyv++ZEuEiWEf/PFZnyRHji4vv/x8eC0AdE+foKYesmzFrCYOGX0uUGWuCHZQiHUIV9e
61fbIwVhPxvbgv5lvJlly/L7QYLtgnmjfvCEV3KiDRhR9zIjpepVEUCRmgbfysaCS/vShAaG4J51
L/dRxFdfoXfA6a5pnq2f6scialD3A41ZJ0p1xv/ol+UZPXKqRiqa7c/UY75FBZtcfeKmYxHF969h
N16laaXLgsx2WGFolX0kA9/ql+rMPJcqJwSS8FCTtw22gtMUxh6E+AWdNyjoS2G4lWVPS2Z+s/Bw
A3B3KqvolL4yyRMAjAEJBn7OM0BxKC3OaYVtH913+I8rs+g7qW9Spmwr705LDJNqa3erWU9PHe9R
m8xm4U6b/1ugDcAM5dsxrl5aPsI2FDh2czXEovilQt3YbGMryGsDU6MZxX/yTiCCX/N+kLWQwnEf
JezNMKz2FDFRBBBz7ZVW6vob5is1Tax/wjDZ8ko8fWCM/z2tYDatxTNtnpATN3EMCVixh1KURJz1
+LBC8lUv9wPc/ycOuZWbpBlHppYhBB4mBK9ew4jyWaq+riSBj8b7GcuM7bShswxGuer47+IFhGdi
brit8nBOlP+Kkae7uBCNNvEuG3jRpwvATJ9GlAY/duCRu8wkKYjPSNbDqkfY1bYuDlSjuBq1Gk2h
3TM7VdmMtLYUcjlr2f2Ido9bYdA9Rfb30/0Szd8V0qSsfuPCqau2f9hId4bdueC9JsSukkJVKIEw
xZPyxiQufu6SLvdMs0Td0gC9BSv8rFsnFg9G0S9pkrym/wSKPi6HmGJijXc6oor5dzL/v2T5x7fA
1bnQDucyW1bfSDW/udj6iZJMOqhpZIL9ozTU08ZReFsInTfkrDNMjixEXaGsV+KebOdSTI/sivMp
RQN4VjnAL4O8QU5PXLHwol4Zg/qqyf0HO8lggAlf5U7VxLyZAh3B2cO9AiycpiQ/pSstoM6k99k0
6iPIMYkZ7rRSQJK3HszzSg82NCY+mSBgUzZjgBEyILc+/jSEkvLYGkBB36d+h8+LAsWPHFRhutS8
qmsEAH1fj9gIbwBoi3c+hXQGLRGwRejp5prq2HLiOgtnwU1B8Q/ypNHLQBpWYxWzHjUs0KPbltmP
27yUsMk6BWmwLkhtJFGEqYNvfg2s45MlTae0xCAuc+wbWlKwi3LnHd+rvRHKAQTyTauEXshm4WHA
5hYdc/qXhmmqED7U8TkiB4FjBoA+4eGPwrBSF834qakix1Ns95k30D0TQFMl73v0U4i+9X0zVfJP
c1c013cCjlCMSLQXvY18EzQe1Fbf9IZJjXmqDVteK2qUtQ9jv0bsykPWtv1zjQeI350SpaVCbTuy
4xYW8j5rnZ8HQN6X0y8KVeltykWn6kRyCUYuxQRhuUCdEAP1yrotO+UR1o6AmGyKPC5v3zXjusVA
pavJQYjQp50Ig8o1CM1tF6dneITxZilSGfHDNOvBOWRJ/atPO6wS8Le4F9PAVbjMUNFj0XZGFpi9
yULlQ525b+3latJMRMsjsfitn44gEOX5Bvaa/pN54Q2QZT8FwRd8KSjyMccWaC+BlcpBiK3EaErQ
PrVuDtHF/Y/u/AsfdcVHAjIm600hntF4Krox4eSGYx6TSf7dyxQZ3o37Wy3W8zclTE687FCGAzAy
lUCO/Wnsx8gVc6H4qycaWPpfjNtq1JjO8EGnn9ntgNgXIf+cdXsXrLm9eSWBWfAogw2gnmhoRf+h
w4JpSRmvPrcEpLatAXAXJlxJJxpi9cWSeVfpM4X+HWd8hJmRTPsXus1v4VhbkHvhwUrblcaXCtww
6kvUrhGoWIvXKpMojJv517NHlfsDIGFKeH+aRU1DGSfiHmYmxah0WFSIuNzJsrH/ywObJ7G0/yGk
SFAvidQNkh0bmTg2XWWmTXd7vFtl/zBnKI6ZBP7mfVhOYjzzmrXK5uVFkIShWJDZuxre91+yT7X4
mfKFc9IskKt/Vr4Z/z8SYjT5WiVjj0OlsKSrOmm+sMbs8N7NvxJdvP98vduzHmluY56GI8QLk89m
+zJNCIkguYL5mvk3j3gsZ12+NNqLQHYIur9ZxpifMtp0fWRHYC9wFTInzk7q56iOKUpv3TfYog47
wjarN8lw6BI0IyMZxayGpZ82pBYDhzs6l8JZNYuc6CrrIIm6CpRz8O/uQ7MMekffYN4ukjCBixYx
R25hNIBKYEODw2sNIs1ltLbfJelEfW1Uaf+0pyrNtJjOuoXr0Ho4RTdFULYHqEHphogcJpoRPSKj
H9vbvfLVRnnLr3jYSVX8cPpmDY0SeY+kWVWtixwFanJn9ximzMCq5zByK2QdU5ptMf1iDfQwy5WP
uBHQR3HmSrx78UEvIJVs95voRBe9ZD9gRBs+yk2Qa5PdNzlOBhjb1AbPfOesMUgO2ubX98bjuuJK
OrSQYX9qPREdXyYNIGYU1UJaWmMIyFzL1e5ZnTpnB2rW3Ky3rdpNU65VmDIlVvz8pqaazkQyf5SE
6rn7kTbIhWQPEUmFN9swehxTqF/8ERThZf9tiUS/x/p1OTADPiyddfJxNxN0bS06Zyrce823O4ah
GIISQWQkJp61UpV8ILOkWR9lp9RFhesAjshjxvJNBjRsJA3sYJaKzlwFxYyzvG2KaHAUFH80mfDy
agdaRJvlzYJc8r7B+bSJwg4mCmSHbZl43NmR/AjgdTUW5gH6cmva/0CXAWs3XT1qK+zWjKMl10sR
TfgE46NgdaLxwETy5roeqrNfOpJ4+Kz+BaLLa1jUqdBOXo2cQ+4YgakiGPmu78VJTwis5PhPX7jG
gO0iIh9vQc3x1RWLdbCviQgxiKj6bprIrLXC2WmNkPgCbdT7YLIxAjbcvU3S+PzFkmYYSgqUqg1v
lYCi/c7j8TbRDC+g8gyWgiOEZ13ySsP28LzHHPwPSlko1quyhyb73Jx0gLAN3Pdb0Nl3u+cgKomT
Ivj5Bxkc4JQNESIRMEWfRF+EnL2WXwcpfnDbzVPLuj8AuTbgsvFUatbzNyMkvrZjFeFwALXTbvs1
4Me5BZqOnRsz6l1ruSbzwZrWK+T35Am5FOusNp2P3TG0dYT40Y4hkvU4U5DeXJUEdG6yIJ3OCqYZ
9KrcoGcJubnd5YtIwRigRb6DNV8/22XRH4yE4NNPuhZ3qls/b1p6ygkTMxPYGCKuTHeTy3YMBvsZ
E/g+1xk8w2WJK+KMpmLz/k6PA5SpqxpBkstml48dt8oGC6dMHlF+hicDaGrX4FUDitZFSGjByeaH
AYiUhV5o4dtvdNULVF8weaIcs8VRsE376Aj8U5o9fFsUjTl6aTvH02rmItiZfIQ00GHIUD1xLiMt
fG5LFciMxHs6GxGRFqDN95dua18+kH1cSHL3FhUNZKqz3quNON0IzvVVlt3JynpEnrG6G8ZrUWTG
PwcnWGC4OIefMCG1dJpGpNhwudKVcWtk5S7/BQUwdg50c3+qENGIj7rDxOWMo3lXKXCzTNBYjNzU
PIRs1vycbIhIytTPievsofD8UCrxASvjSdsFyHKXLZ1ejQR3ua9u6oPxhx31Ph5wFMOBe0mXsOxo
0jxJDmaKm9Ph7Zvwgoc0AOhH1PB8Gp0HzMVAM5WoEYkQO4jRzO3+HQj8sjC9DLG+Tf8LyGoF4TWV
Tt5FrvcUVDfTEk2EV4hON9yQu7U7u92rZlKFdpr9bH5PvZ5GRK4KCDighc1LCfmXj8TqfY6vzwR+
mxKF2p/6VLCJ0ZqRzjAZs/1M6M7MlSAWwnChkIkiiDl35l38ZI8kKMKvYOhwwcxVV5FaZR25IDGW
NtbyjAnGG0R+CV7dm17z7L/Ct+V5wiEQY9eP2IdylrVL2Q7Xag4QW6kbOfOhLwBgfnUylTL9W4mM
g5UWYZvPdHvZiWzp0moI+QyOfANJocJRAq4d3HpduF5No1GFNWQf71mVQsLKd/DVLyEWHHioucmu
QapKMNvMPYuGwWOlE9jBCTOgLMKmI+WcsNqnFBTdc6eCa+CXVOfAlHFisIIbnzKqnSLPUHIuadQ8
EvR/H9j/RQdDlBYcOlF2yqHQrQci3duSdmkciq3HTAsjgz48PowwHsBwmrIWnNIs7YBOBAv4WU31
rYzID+Ysx7tMjgJHUfAr11DerXKga5E3ADd1F+Wg5mW+Kt0Pu+u/8zlwlHUG3bSSvZvmv5R2JSQE
X6xRRO0hkpaF6URwF1REmWDmWJRJn8t+4H+TNtcSZqcl4PJS+Glvby/wA10WS5u+6kJr50UCNtIS
dlMFg+w5bv4RsAZAbiwFuns6v64+ql0riId7Nx4XNCx01msGVf5K6lMrN291++JPZHx/JN4y6U7g
AL6AvHJuc6ISQIsPcIVjbdPQa+B2PZOSKRr3auzRDzzgUaGxDS1Q2wHQrizNBEtPgFIj7RZb3Odv
MQgY7cILB5cWwdCIR8NhXFZDTMs8Ww41xSeh42SgvZeCzUzgJIinFTkn2+lRsNBAhY2z+huL+vVc
HjSITz9bPQiZv4kWz8On85nDKNpwG0PPt6LnkDm/3R4asbnUUuc3Zx84Y2sc1UYj37SV4p7HTtcq
0aTowwGTcINewNNWeV6EvNQDruvdkYfWWn8nagIacJRik2ah1jNaJCDPtfCre4MRYm364dQs9gQ/
T262xJGmDgNX8dFDgi+YicFdGffUQpsArqh7q+S91uSgCjWo6X2XbKJk7vJTUZdZ6SGkugOnx4zj
JVIUBidyNE4PfOLkyIOKHRQCcddPXOJWB0RgUVbeTkGF3fkj3XHdFMmmdUa/gMMhfm1G9RhCCCa5
tP+B5uKqnCR6Ttxman4U5fxg5cN6wZMx99a5m8zJj4bvvTIjwTt9garLfif3ADGnFjOC7Cgg39Cf
EX86v8gLeJ9d3duZyen+I3DJ97sQmCHgY72ShsATS+pjtZuUOS2KF1m6bBcCUxt8mWAEJwvwp2jk
9C3ZUaPVoXX2WTBJFlJJpATjQHDbtapbF1zYX9HnLq2Motqm++oTXmrQErY6otTOgABkGLI4rU7R
zT8ZB2UldSReho9+QkOxqUBo/vy5XE4SCFF8VCOjorbzlGM6dSiV79Qtg73w8pM96siXi76ZaQrN
qnHq6v0XTzLcCdx9LEwADzB0CEXW6I2BksQYqhDLcTVgFxqOARZq+xjYuVqVceAis7SuEEtcwYN/
dSxfgJLWoEr2CSZubgoDhEUYUM1YIdxgwHxf3WetVSh/uEtdNGO0cp23m3ZNey28PYbalBYvSE21
SeGfz56EU79ZOYlKfJ0Yd8SGpqZnwjyvLr0cq9hfWhZ9TuNYEr6NhUnukqcWosriD/eYpqeKtAL7
42Q4KudW4emF1icgGSlky0FkOtn3S17R2pkasS3OfdZjWplAm0BKnyIwvPCw8BO8Wg6KwMNT0XFC
19ioKwtC0lR82dBqYA9ktAjdAq9/zJB6mwnljHoVq1xpq8+tDqtm1zfAYu1eUXxZro55+ncHm/W6
0TqA5cMjhf1h2y+UjYxvjuIq4+7chW2JTQ3loa7vyqaGrNXfl45CTfORUzjT5tbxj6jWLQSjhTYG
0PPaazXhaKkVWbhG0TPX3hpj8S+YPe20iSBzNm7X/mcDS1XhIN1mzXiA8WCa1/3aBWJuTW7XoUHk
p8o8+gumVAw0TeLIKD5ihWwXfkSGyXd7fYuEIVUzsPpGo+2rmQsyv6Hp+syYMjf2SO9WKuUdUmRU
6DwSmGyZPD+5q+CgM9QjOT6VYwo7j4Kpi5MNjuyv0+BpfJVZ3NUDz1Hfh2q3HmKzI+4raSILxbaK
BaGenGlI6oYVpnrKTbFCO5MRPOpBoUE2nXaYc7htIEFnlJ5smBFRVJZrQk15kaLQwwR6LWNz/iHe
Ba26rguOsuOUWhLD1a6YmPrhbm84I7AoK98z4EBW2JHODgGbyacWjsYr3T7an9Q9tWBbJbI1S4rw
tmWvxQ6yU6H+WQECRUY3wasLNp3aWnLSuju60tYrEOBfZyBXPCiYsUBNH8EaT/BM1XXByB8hyM+6
lIl6YAItqfzSv2edsFkR9MZwwsd85wdVD7/MYnPuu0BUvF8MGi6Psw5W3MLC5+C2ozeJa4LRcbwp
poaPlk87K0yb/2X7twMTjOWbiRs6ckgh/URgOEfebhEto6eomQIqrH6/g4J+KNEVR33HGW2tz0WB
Sx4KaZrX+Fi45r6SyS7TJ1IQdM/rrfGs52gJhQg/ryistjOkb0GWYugOFS29UAXigHUblmc1FjuH
BtA8nr0qQiarrOzb8XAy3ltMabY0bAbQFzfuP8HpEEvbNcDtvq9rd2EtkbkSIFUXXPmwqyUS5KOk
nPuhWlaliq5IWaav01iHFtqxHY8v5/pIRE6DbOtDSfV0r8r7+/CGDu2i9XMf9ddMnG5vzi6b4Tjr
zaohpShb2hG8E9csfu2L9y6VbYJO7fq9uS8OEMNxxfXSksll+AZv5Plq3HTs/tTShpn5mFZSxwhT
Cdiz3KTPmBlkrrMwXCppIP2uW+aPUpDUpOcWF3qKRArw3HrCEEjz3tMXQ51H6jNql9K2ENGGY+TO
H908DyttAD1Ih9pYiq4adqFFBS6tRRPTjiEleuidD7V/Q/l5wmZMJBA+ijMdM2bqfYaX65HbJUbc
NtvMWuZ3ZvVaWxvQrN4Dtp47YIWUdNa+bcWDFQr9EyfnNBaY3elLpr4RmBGs1fY6OLwhJSIp+Vg+
F/M5d8zeaa/37lF9sDdh6R6V6Zwy+hge6zcGkVn9dAr60IYlmsV4Bkb3mBdZuTe8tYR8ZtvTQolM
b6QHg0vM3NB90aZ2Cc5gDoYcsVQD54bYB0qRsk+L6AzlQHhZCRycxNGI1qE+SPxQVKS1egSQiZVD
rFfybeV7e3AzWBGRskDLTREa321sDkjrD4tY0JB6+zzq05gDrC3p1mjLOencsbF4AY4XqRnrlkDk
G9zKI2ctCkffqjVPB3YXM4fCAhemZ4287xcyOHZazDcYGMMqqBRvA60D9t/zei5oftWhANz49+Hz
iE0G16Z5YvDamBSnvm6LeugZ6tZ5EOnTvQHPpvwAR8laVMvSiUEE8z9w03j61httL3aziv3JfMU6
YyOR5qxH7hB23P2qIEDchJGZi03NF3O6BeHrqH1EW9SAGSUWruUQ3Ho3MX+HsTDYoJ3Ulo7HjxUU
elTnP0H4U9i4Y+PtfJefHv/TF+3ATSJ7Wx8g+KMgMKkvBGEj5b4kqXlUopxSdxhnFaseIpDbVYBy
KtbdCBV934nT/QanUCzIFsqmgtm56xjTzOcfuoK8qfAArEFtaNHrfZ+31YwTYXl3D8BF2FxMIVPN
GD1jhIYZ/TitHUY/IezV3tCGO31OWoc/Mqmrz7+SdR2ichzE9klsrtDVEBGn8Uuw+QFma0mhXBSN
OljJew25JTJTPMZrSkJoZU8LAzq3Lvw8d+MtoOxsrrIKO1o7D9AZAY497QLDc7H53bZOnA203veJ
fvmbyMMP0dT16I7HdSBmxtPZH6F/JSpvlDn6bXgSMOW7ZqMtJpmPbdPbWNhlefq3iVbldXrErtUM
40Y6exEzSIH1wQEGwzVrEJxtjb4QUIoX8sfK7KbPtvl5uXdUYScz9d92yvTjIeF8LoFZR+l6C6a0
XcNnjj6TIcMCjIIss2Cp1AKCLOOq5S6FwATqR0byWPlYs9i9lPVOpGeAwVy9VSD/dR/1DMaxDgfg
xuh4tr9wqL119JyUWEUW5fx/uv0ooCRi07u7fiBYNIJkHTooLzd5/r5/pL6JZCWipbG/qvZWEAIH
0GO7Mpiz5AN6S+KG2dJWdjR8oMihwh9DYkgnT0h+6f4PgY4sepGUxSL40s5uvALUOf6NpbcUYi8p
WQPaoheALzgNDBJGmPP0pSw43Csnt8YbfBOAS+Yxn1nFKyigQlN+PyWlv8a00uRiNhztZ8gQXvgm
iUQJsx/vyM6mJAJfICSDcvq1RhFodSAEeqOYbjqoyU49Gdo/sIPMUy543IKy/erXHmtwFxaCPQY3
nTZetkf5c/xdIV6SzO97OlX/3DOY+r6CZ7KQ1oBAQNzODPk1ZFNHD+4gb0PbTpiyZjrDWKZr/g4C
ig6xvM+u708TrubPI0LWyGpo/C4Cm7/w8OypZWLYd+vW0cXkISTmIZCOT7L2hcwzgfUMYlN6/9Ut
WSjT7IiAYs+RsEGS5XGgBXyLMYcYUoWReQtxuULz6Z9gnwqEZjYARBODRHP4BIeQwlR4PX2pSb6e
VhMWXXUGdxn0J+LQG4s0ARKl2GIYL/j22TDXXZd/JeKkmIV7S/LlEiIDVw8Zeq5TTdCeozRLC5Zw
yap3OtCbT+snZdweBsP84IjbzwZJOx98q7edN0GNSF+9VtjOme0iJVAqR/5OiJolsFH90P0lx8/G
XqTe6NMb5ixSwZ12k+3vuUuLyX7M3YaOi83/kr9asEWcbijaaTNYBg+SzfR7oDBs4+gdB51ZdXdQ
E6ucb9lQEW7T2CfcgT0NJmSNK//O7PIJFlO3CMyGVuRE12rnj7QCvGD0nT9zywsE7FpzUthltI/P
5dApA07D3mMKdblG5y2H/TBRY0K4AOzDRCrevVLcifgxD3nZYW3GKdbz8/OejzB3fpIn0ZBYukF7
vDyzOOUTfaf/8cl5+GgSaeKQ8+ml9489G7yajxHFXpGbNsHXZ2eloj0gve2R4RgJPO50fxy76x8j
NPuBH3G+V82wZaF1O+kjN6rVV79WOmVfZAnzk1Ni0/S7BN30qpGJaQghijOKyyxz2+4JU0NoVziK
8AwADKvYWkyw7opu/S9m7yqrES/30QFpCVx1NBcUVemwIRZRYBKnDvdMd75J6GFAW5/uBpOVJXyr
9cXGMifHs2/x6czKmNTwLznGMssRDYx7xj9cyDjG8xUcrSpPTZV2kip3dleZKWmwFWMWk6v2U57z
fB/d4ti3ha+RnwJEwMu9K7bh8Y5Rw+MkFUHjgMgsdjjv9WYYrwUzbYesqImW3+kPBBak5zkdZyhW
wGuoSNIi74rrafQh9v5ORl4QrZMbTgKQ2+dA2OTYu9Gl0+/yogmMuclifKpvKVzI6Cr0inJsvkE3
lZPx8Im0w9S8wqG0cmGjdwdXpSql1msG8qje53iGUSIxZCj9g7ISgctHj47e3nwIW25BopLFOrHo
eBFDXWU5w1/70u/Gf6sWfaBOW5C7or/048sQ9/v2dglj47hsi91mOZixRC/d6T2w6C3UNmBLPrpc
hgdewisa2BzcyhNsYZz0g1OKD7iIoOeCRy6KojCoBtJH+iWzlu3im/O6dZd4O3zNDsP7kn5Nyr6q
j1zm6w5AF2F6h8V5sZ75Tm+v21UpmsXJddLZCYFYkJ+EJXJfXg9RgbsoubXH3H3oySbkTai6sDxj
5QTLQ+352r3niNFHY1cJMOkiwoT5+FzwRZfsLrkdIOQXDLWXPa7Hwte1q1fwTxn5EDClDTMA4HCE
QnFuxOoiT9H2E1nlICYVIgcvNNRDi15xwJ8JKq+v4bW1Z0fH2DI1FKHt5bq9EppbyskHEhPWNw+N
PNGdKv2m5f+0Cg8amT3kuJjiSTtOReJvpitBQ6wZ2DgF5IXfGQbQKGOvEO0KDXLtw1G3EByYcLda
8rmGwLdcUMocy41Dqg2YE0NmJpOCzDze9uJ8ZRk6Cr98q2bX/vFrrMnY/4g81ozj4/vLt1buJ+Lc
3R7zyuwz/ttS7aurYeI1pBRmLJ/CPbguyIEHD96ymI3xeF8Dfr+vJzBr7LIrQReW3wNOKYiRm3Df
CE7fALcpzM3V3uZdHhLjIUtqR+2DWuBWd444GVxbUa0CbbY2FbzMfgsTvK8lDfqXZVwCK1ih0K7x
kqOKlIlYbVAVub6HjeYzMi9fQtR0FTypfJFWLBJUuuXllzWYKDIlNnM2YAzgO76tAdtTfGs/cfKx
HL+lANCd2dJFnH0GIQpUDmpUiQAloUv8SXLajvoLWtUoRS/0rXc0P8Ya/NhEVAfTnbN4BBN1RZI3
bfIQkgA4IyN1MS8qbDvUlf0HMwYzc9i1nSFzv//fViwOubd4ZR/OhvSE8WtrZboUrdME2ZC/eVVy
UZfysgsgAMyclGLpr6T7L2/XSXOHrNArcL2CoTVddP6VkNgR4NHcYUhgHp69GM8oU1DDj90cLK/s
cyG09NgXOJcFuidSJ7HDJocC/BBLSgHIYPhK2L4bEyqoQ3nP3tphLb8pCdACHiaSiOtEmVTx0DMi
tOBDrzYEwA+5jCl80B53mcoUFcK2jmI0K8tqudFNJvD7y0mC9DDGRKhRxIbIXjxMQahJel1XDU8E
0bh4Qr/ijscFMKrKeQ4/fAn9BTBCkTQ8MbeU8tI7xFiRIzgLjm5u0ESA8EtmSbjoPEoEI5nrPLNa
OyJbzkzVmBPq062hubIwmZhgpVkrYTDtit3UBDsb0vkdGJyVlB+DWN0tSPQypHQb7M2XiWwRNuIy
/Ec8+fgLHvLHe/PKsV7mF4+vPGMUytzk5o5CwRkO8cREXtK+639iBe+DwM6qv34gmIgzTwBf16Su
8HoNCZOvoJK89yeRpPZkm0mgDNQ8iIL9XePTHv4ugODvaDa9SXikU1uoErzBWXvonkmPXlrwZcpe
gVkhkehnVeU9dR6gMezhRVbzjrZKYlZYAoS8jUJayZHtWP/SSrdqxwBpWaUjJWZuS8ZI11GtM1MK
1I3gxk39PMpDCtvJOIUyl9b23X0Jdwp6i0Q27o+rB8RwO2Nqszd6pzFgimMVd32mtbqpZdDlZvZd
s2bhdKDSuV0iMoqg9QN/pKJ5VkC6dOKr8t27CcJGfFI51j8oDXn8DizgRD78UwSqMZxBWoCg/D7N
D4yKLa5x949w50Mwx3Gwh7UxdjkeEXkgK6yw34DarNBBQY1xXU6ydn4+WrRf26hMDn6jcmXTgcmV
uUyDXJgqZZSmR21xB5ZHhqUPI9CiUt7Jnsi+nIDPrdmsU6AKELTNhJj6yvWIjri/teF3g/msmg5d
v9S73TMsBg6PQv1Whe1ba8zod1sbB2lSDI4EBzH7fRCleC16zX9suiIfBbDU1dEILex34AXGRDwc
89YZn2lm/c+VTydp21PkW2rkjnBPjuSj7KJ9pcQpbTi4U8NU5khEsBXxjMzmprqqc+zXO0zcQvFk
Kik7tdXf7xCly2SaMwbmVEkhKKLukmjEUhy59biyGDDIAgLSDD3iHkddfiy2tBkIaRW6OspUZ8EI
x1IAOWVidY25fzG6f+XbK45xi9LYih6XbGws80CUoZpJSIyC/DO0dYt+0RI/EyNi9i3kwxOuanrd
he20Hp+wAEMUpKrSdOuBIWQGEfP+ZWHe2afVeNXdsHrde0LplF5VXwD/qPNAAjKaoYl4yCRR5BvS
Tuj6AOgH9XzKVFYpdWgU4jl9/1BkswIhnPIXb2t9hFc8DquySBVicghL/QIcJjj5pcj7yJykT8mu
mfFEvqhgX1F5qqIeSfV/OuniukCklnHpjhEsNqJY7RBq/6MxOwbdlrWavhhi5h4djocjtbKmzxVC
E66WS+gik8yyKkGjwBr9tN154qnQ7LeeLpyx4wpH3ly8Ph1gDNRMmjff9OJqGU+aasKiYHZ87kuk
aX4m8T84Z9eZejM2ycySs7LpyLPqP9HjzXjruwdOr7EsnW/g7HPwdp3WwyL1koKu7SQHTaZLOnmD
mvOP2k1c3JkPsyjbrkAYMqvPq22xTiLSO6pFjpzjeP2DoGxmm4WWyhNbGzLhLRbLMHsu78un/3xZ
nRUSx51KpCvJ8/uhE/5tgl4TIoK0K1hJZB1RCqAEKHCFpsDWi8ms9jN6skSyb4JQs2mon8HGgilO
gilbxyVAWqXV687bGpQQp1rQV/H19IGu/SRYDm6g8zls4c2cJ2htp/cn1J1YMUfWJP2Wsyifa0EH
38ZxlNlcPcK3lcZZ3Y4i+VQS/zLlqLgmwvOk6Nh1HhYgSNcAsGJ8Rgd2kYhErfjNKtjBeRodSKxL
D38aiwO2l67fVsbYbxZnXOTmjMQL3+C1ECfQ1NoK1nQo/Yx5Nalma92lJoo6veeU2cyeHt1fOG0v
9OLCQCxB/qs7R2rQy/f57XCPkPd2QUFHsF4mkCXYfzC/ZPI8IlEbN0/WZ2GdwW8QdV1ZKTmVt7NW
eJF+6ykoh5VQH2QGsVjxDOga6EluRJIgZp8HDWZY76zwru1OpDzf+uD2iwcu73DR0Bg+7Bhf3Ccj
gWSsiYuKsar3hdaFyDFeVDNmlDkFrRH0Tl+pR9mM3WyMj0czoitziB21VfcHfOUmxVc/HTCjTR3E
jL7W4eX3BfYXXfmWzHcUhTx5Ijfp0lWVLnR9O7LAk3vbzPdViegiZS6GgncHj0U8Ka+/gMSdACHN
H0gOwPCxoJuqPglkloCpk6QpZp8xBpeTJZwP04M24rQtFdZEJWb2jBTDhtPAsD20pme/+oQpNNjH
g0sTSd8hgjOu2VAQRbOEH+sGLxP3rnolD9gBZEqB4VDJOZG9nkAmhpB+E1slmH28GWsl/EkoqaT4
gtOwcJsCc5o0BsfoDlJKhL5S0YbnB8YFYqmoD+x2895ivxuiNvk6/Wj94/SF0srb7gPJgGWbAgMM
Ty9sfaoAxRM+j4GEWZdvn9hkAVUTOPjqt2p2l+AC1z+PW/1mhm137Cfpak1oxd2C4P07lzpKuSUm
gPx6rMubkwRLVTlV27HXG/tPP831yRtyrMNa46Wn/J05ZEvCSC0R7CmRNg+NhfclqN+79bRHUy/r
Lb91x5knhEC1xSzrCJxeyFHV/1y9LK1CinZTlK/OMyasJ+9ZwcPKB0tg1EIDdDFJuWnCgfZr18y5
MMcwc2ICrrDei7PdzCsqkz+GkDYFEEmjYGoDMRDF36CkkJdMqWpEquEQQfgGbpFU4AVIKc8bHkN6
r4lOzPkAyWRyb+P20rXjBXjhrQGmvoS5ggwJYLQHoIC+CqQSuq4AN9I0c7fz2emHftDPMTDsSzkd
mW0xdluABO3lprQjFBXgxVCtDY9ooyvqVrhslRMYfklDsBn9CNAOpKPZAhFsBZ6BfGyaJtWX6AVN
A1reUuozgoK2oU0k0uOgaiSFrp+mfb6SEDkpMvbBr7ItbO0f8u0Q4CG5NVWJT1TkQkGsyi7FYWgP
0dUYRYlrEP5WBnv5NKtkWh0b3sDpwS+W+4gUC1X5t26CfloDO5ApNMB+el5feje+9Cl5h10OjLmm
14JDTdSY6KQaOzsrgUJa+GhrKoHTXEZXE0ENhmGNLykYsiQuzZC0gUykK0tSfz95i9Qjt5IZjhli
atL3YIKKwkW0lw9h0T1rEW0lco2NVsEegQ34LLNJRM6kWdXbj+B04XP62vWxKfb+bVSMAKWyXkkP
Q9qL824vPEOW3d+y5IWagL85LPpOgeScumtQTgyijGaUdl8ZslF3JNrXG+Y7nUYTPmWOXuNPfvcT
lIACwJI1wNcbxlVKbpIK7dKFjgAIt7IEjSkbPC12dDT++J8BxI1SNuiD36nPbSjbwaS+FrdsxuFO
bTHNHMsOLU1VRNXyVNa0F2rByR9+pkuiWfwldri0UybuC9R2yZLt6iTmmO4xSa4cNMySJeoLgado
HpSGpnCJsNZubS0TI3vJ9ePRsUkKabCyyBK82K39etNyz2a/AhQwGykrkFSqEWrvK184ciKsvWD6
8Pn7x39y5NcYN2FPwpzBHeAeOMGEaRvHmBahn1WiQYsuAHZgwyhfqQbcXSELr1zzKKjXfMxEyOQU
BrfH3jbJkdO3ahele7UC8+thJYVRJT8gXkQ1N+frrLEILe1vhTP8JSI3IIyFqpyeelY6DZZWj1xs
8ihHmfICRfFOPwSD3uQ3/idtVW1pSCxD7KV9yPwNI4tzRLeYGFFoEpAu47SVAiFFBDuHxpLhwRyO
SEKQqwCSfbpi8bPq3AmZswsvhmAjmTYkXpUDaDj+6hDIFEs9AyE1wvyyGlVag/T6pL+zrTKEYUMJ
yLp2mNH27X2oKW3rBymArwk21gZnbrw5wAIickCdTo3SORyF0CS/+42tGvRQdFoteznnL6kspTO0
U1hIb7S/R2ZPRyOP+89MRSwyD1jeUJSPI+Uw0Bbe+HZ1+PPf4KN6lbzSgje2yOhmUs0hV9ALpOmo
xyqjffFBlnzAecQgIU1HQExMI/P1sPefnU8viIqsx4e4MrPxdlLevQvNtl8//b7/MMQJZHL7O4Ks
IfKjRg+gVQy+mLypCgoJ2TKi/XJjQk+ItoTmIG0dTJyWYrvaDlCNVaryl3sXutAojnbw/ZxxR4//
3zebODUtu1ak4h8IDFtQzoIDRBUw0SaohyOH4nYJ5o/NfjFLuA+6pnjBc/ni+lpWrNJUYM/XokcY
/5FszKLQWXYIUoB4QRyJHb6unH/R4iT5bKJPeUovOV1s9xoFPLHAPEL7w2DYUg0h0Cu8MVpU8M1H
M1V1QyrCWSXMY7fon2nNM5LYXe5U/C2PRuoZkg5WYpTrWcS9FS07nMS2ruo5u2bx7Wj6LlyX7veN
+/uoS0k+M0ni7SCUZ6jW40NZmJ+EzfWrFx4VQuLuXE+TzfRy6AXHJPkFnQywXG79VdqzmtJ4mp/Z
yHS6iQtIg/dwwtvkdg8s9PI23mI51ygMlRKhMF4WxWAtanKzyEvQqWbP9Xp1eSlv+ogDLIwTYTor
hKUiPlpY5H1koRSvs5yTatWIIXgCq+LjstCnfoi2WudvDzTH/SpDLE1xlC3VJieGHzLA4I0M5s7y
zieBaeslRBmlgWehRUPXF/W6NmR0mtv2I1rrE708fs+OHceFt6AgxQV4DxRrGFrkdP7gH8VMBy6j
xp/3WJ+9bgCEkNAXEtL6SjXMMt846DPvK9PJKKrXtsVKzC4XHH0alHoymfWQzQbJaVRLNSmJ9vQO
DRnzBOejbRnPpEE9kxCnA+kftivGqEmLuG1u2RJHpWDTWo0FngPE8vGkL8aiWBw0TNS1Kra6MH4O
v0a5iPiqKJd4rOAB+D904Zoz7S/EFSXkLgqcsS0dlU8pmOqeczO+uwmQSJFRc/wGdJ9+dONTmzsw
0oh/R+cQW43GwizQVb1758G/LmaXtEhhQD0fD0kl4iQ4Kp4/OZAVE/oXOqQvFEthdJ+/jK4+dSNL
UDR9wYwfw1UJ4z1gVfmvur+KcgvlOEytckAx/zRjEkEtWGi198VtcIQthcPZpcoNNPvm5G2+gkM6
gPjVny+R1hYPe1x0UObqcr+ZTOE44nXJDqXYIA2izTyt15kgnPiVMT/zCdjnUS1yUKmzEXa9H2T/
RwVONjj4AJ8/mS6+6EzvbZFkwrcmA+K2PhFVL3sSnWpjRRQSpHHi8nupIFkqn2YdnnXnwlLjFz/W
G05l1wwgvgsBqsnEfmWyC0Yp/t376F1InzsJv0ZlmhkGSLe/TM7orsDITihwRgAXSLXmbNQShmWR
d5dfBqbTbe1tlEzdBMq0VbztwTzE3hU7YnZsJxRNGFf918nawEsMKTWSqc/dfjodFdVGJcUyzSzf
jMvYAlmUcce6ykgQ3ETCymr72kO71xDfCVmb0EmuVQEzLwT847napZat6mXkSeUFJ5n3MNyxRBHN
QY0PYsX1rNaXvq9ONaA+ZpxOdIz9/YslpTUR1SUnHxEiMYGFZIY6tDz7e1TU7KVgMxr+We+yNbFx
PGfWeEVaFkamBk6kq1UA+cP9jcMOYaSDRZEl15cUapwBLv29h94MHF0bth8eRxpAlyAnQXjkm/Xv
T9jZlA5/qs12W07fpeP5d/lHap4FBR0UL7GroC3Xb+ojrq0JwNcJPbP5RStbF+w3fB2fbrgsWHLi
oEVBnkW6rEU9KPe6e+pXG0sunyEs/7s2QSX6DLQyISU92HvkIO0laXu4RinswLd1ressI1xn4JBy
fx81XsbHsCK9ZzgMV337J7CdGTglQ4j8mo2GtV0T8VTOnFATdcYuBq9O8Q4IJNjtRMuX1OgwibG8
PXhGqpobZD35w2u70Xlt6Jfi1v/JfToMUkJrpaQ2ymwCXVQURX2Rp+J88BlQG8zAL5lvlsl2mBjW
nJY91LmgUVfl5sRsASlOMca3L9EVFBodIFQ5qo/2FFQ7QViH9oR7n4BQiIgRU/J4sipXsnUUHuK8
rX147FcHsgzYZk+FiCfcecG8jcsU0oRNPU263wBCgdVccvRq1dRgcUGYg2q2noHlXEq7PJS1JmWO
BKlFjyWyWNlkleefXoN5oKTDvs7f+zwRxn1lrI/iMpnwTgJYcxL+X/YOCY235QYJfceBs98BHJD5
Xcilw3Pv9GjChHj+eYfktdWIflbibUR+vyMuNJxa73NAUcRap4p1X8gWEcWVEFhFEjZOJCDAmjdr
S8wqqt5lmT5WiyuncINk8OaRyNQzB7thD57tYyd1j7HG5IfXsAyPNBimGYE+OtnOJck4miezD+Mv
JGly6KGsgIfizsXHIbCMEko+bJT8nxq4VNZGgdpzledHjM9U1h4brDiTcfM+ePESOFjAe87ERgRf
9CHvZSBOeTlcFJ5tYVD2YBZIslKpr3bAiFXHWNLnany1UlXWfYFWUcfY9muJQnZBhsFkQNWJx5y7
4+lpQB4++22r5Gzz+D8CF7kja99wMCdyl1U8t8ybC9QH06WCIuGLeEOsdO+EBpTBTDpcSTSYu9Cy
SAMRrTf2OiVrxN83mf367pyfYDNXqMABDL0OolREB4KC66DPB9QiTSOLZ2t8ypQu5xkCRXiDYB2P
mwp/dubh76vqN4IRV+waUKd8AWfuUTTqDnESH8OzqCeU+voorn1k7wMzuYbM9+d2D5xRe+Dk+ZGX
eluc5r/zZHJRSmGZF7A87cXz8HDZsyoTeAxTnQvNYbBTOoSqnDbaRU9/uVqLOMnLbnK38N6nnj6B
ZWQ/fepXD9ZxhJ7nhEk+oF+lXMURJSPB/LLNCE5/OZgCINbWqLocWqHrM0psR2JUln/hoZJfg0VR
e1zFBYDjUV0rWSb1qx6qL3yNJ4ZIIqgyc5BsT6hugdg754PW1OZwX6ENq2r2BeqOIe7VmbD5fsoK
ugdT+ee+27iSL0KHJD0iFTxEfPufJA9XEyTOqDpVMlUwQkTw2NHGF+1iqNk9vaQrm+/s77nJ/AXc
+Tn4rcuEleroIwzeF4uSrOZRW3EoHx9hEOPnM+wBz6cZg8NmYK5/yAB3/0UjXMQXGki8rubTZzrK
tKu67ZdFc/wwpW+/VpMpwvGFTL1AfgNUpQmUjUcWTp56V5Cmu4jKpcarG/XUaVlAPAAmMSEkIOtN
lYlvK6bdC0ltswEprRQNQ9CtwxWevO2Gn+wunzjT6ninUoGA/Tb5Sf7uxP2q8B5xAo/17pJ67sTX
ihnIF4NOWkHLBosLuH9FeClvXgRNbSydJHjre3kf+3Gneaco5nVh9Tzt/nqpPVkwlWgYXSVTX9sL
OmiWXmiRxkllQTT6KrRHgDv5zkOQZrwURH139Ajmo2yVQrlURhmbeWgYVFmWHga86tJ8PAMCP/F1
9TAe/38lBuAfFOJ07YFviv+7WFBS9hryVFOSDRMAUVNO/QYebC8hYdE6OdTXGvkopJ5tZwmp4hC0
EV/PrulMgVc7dOpb/uBGJsZAb7RWbhHG/zQKLKT3WctlZWOKVRwtEDoT8WwBgpUHbVMkOqXtgr7v
6LnrwvwnG/B27LMej02S2ZK3HHkaRDzIPTNj2h8aRDPfSTUdmIBnjTr3e6ed0ekMER6dYwRAWteU
Sq14AACRNmOOAypcSZzYGzlKXmLEfAqc3VPwGNUwlM1vjT80XasK1fIQuOs9Uvc0zd7FXJ9E/XNi
62Dfti9k3UJ0EW90H84u6N0yBfDFvq0PAq1puhnq9KOWa0iZ19cXj/4t92fldztE6L2m7FVNv1bd
/3Ek0+3rb0S926kJ4K3TfEO8OHmRHBtzNsMlWxylg+mqcMIOAHYIrDIQrZwlaocYchT/9I1xoEHd
gYw4EcdiONgSS3R6vo0LskxNCdWvMrESnyFXW2qx7O7/kAFWYfifOQZSthK8N+b+p4uYDLCWdb75
PntDSbNImefUq9RKnndzjPomOKDwb5bo0aApF7fjSLRizTNaxH0KQLG9BCaWJWE0+IgotjHyJ26Z
YnYCXD+HCLXrrJ9UVb+1myG2FMP0LVV9hoenH0gFcwWq0NKC5r5cwaoxYI8jlTsAAfNhny7eXGsQ
4LLaduFGQYlDWUiK9PLPy6zs8odhT67raNX8WPYHExM2zqrX5wqBuoK53W5bZn5bempVfPJ+eQEZ
mNkyKW+jPc20LM3DJxVt2lAIn4P+eaMRZZJAmha5fxynqGWkhviydmCQkrSTVgWCzYDc+p7M0qp6
1LtbtQ4S+dWcOhr+TnG1mFmQuLFKSiwRoSmUogFHcd3tj2ASSyOYRY1DCVeah+/XrUFrpjVqRQeO
Xj+LbmGguEq6UfSlNLXLoOhgf/p9R1AVGkEOABmX/RaIBvdvBVkO0J6AcCQDU9FFu00kAXUt4evL
8bS/77yIhOvGkcsqBvPxR0PgFGUkSR9uNVxNS9HHFK6NNgqmmDsxoTCiqOQV6Ua5cmjauSh9VDYX
fLT9RQdm2gx8xcOrmNO6Pj9BWJvBdCHqpUlT/KWCwqtyl8/4pRHGrNKjxI/FTK8qO5C40kg1mJM7
2h+CvoVfF9hvQbCfrICWR2TkO4UumD0Cpc+o++cuQkXX1q2TREcQadTzGxYIuqCLykXbHMp+WIUT
6GwyRuxgsV4K7iBSLsQgV/wu892l/XT/o13f7MoCAz+GBw1abyKRGT2/IqzD9PSznED1QQTYtVfs
dDVlKuQQhq3BSiAcQT7uWv/0DcNjQAFk7xprFOfiUK+9/XWRBe6ApZdc9mtnnPuPxltU/JhHLbtH
8+rTjulXeUVeHb0FM5sSuMHgXoeoDloQ2Qo+sfjwd5IRpNdn0GYNcFRgwt6l99KY5nVU3O6oMV1x
wDHzBWI//RpwsJQp7k9LVyFBBK/TGZBd8HKWHD5m5AZak440XMp5dJ13sfFG/6v/in15YOiw+79P
Y/wXrYV5NeqdGPAXopdQ8xZc78Uru5vs2oqElScF+hppP0DrDXhiIavvv5yynYiqwvWipY4UncyT
UGcKzE4O6vdXWhm0XJW8TutQnKWHm/F32WQ2zSEcJEz6LkqBddVwocEGsSpYpVTE0FZYlo3plLJc
vRmLJwFWPR7gCdD8SOe+xPD0vKqWyldi4zludDJ6EsSB6D77Z5OAKoQxADfdCUlLcDY0rOYdYzTt
BrH3epqZiuBmFyEupuuhVn7BmnlwcxcuZySGE6VdnZygFh6NW6lGwlC3ZvRYJns/b2HLi4lp+SIr
Q5Qqj7MO3wazgrkEWhA4t0NPWsKFJ9MMcvZ2auRU+t+NbO86pvGPQwuLBOtqR5/rmYGvNKPAqaxv
VdvEIUkTGWYFqYWktu+uw1gNgJhGoVpYhA7Uq/pU9Yc/qV2BsEmQirwgOJPVmg9ZF5suYelgf+2Y
C2zN7kM0HyndztOY0s1IWVDrXdNS4uz6RPssFCn4UGeilNuEIzVYjv2ECDrJzveidbrFbMM2rF4a
arNp1oqhUYVlCHD7s87HX8SKdesV1gmFkAJ+CKZ6he2XRt1okCeMN65JXS53Z9K9D3YeibixMTIo
z5myaSDYxYspR7iQxF6r+KwA5vJUAbn9BXyOuuil4fNGXh7k5g9P87kwu8D+sdC4fYoZAdd9PFrq
3fnRFPMsQ0UIRmjVEBtNszE24gwF7DjNj1/2al5hkVgPFajjygI+9oelNt3UNqokx1m8MW5RcgBY
mEtp8UZR/CCizkQIF/0DCwiFZmGbVsGfsiuW60mctkUc0TbVQzmHTsVX5/EkMcSTKfNdq2uVamK+
o0mwoSoFG+zqxRf5lPLcmjasfnizcV9vEPJTi9Kplndt17skkDwlZN9wCnJLqmSdCEuoA/BVj7ov
zMgVlz3vCb02CfnbyiS+BDbiT78Mc4YMIgoailtzi1E11NX7D6brKrMh+rTZLwiWAR0R7qlzg1GU
mYZe2ymjmv6MjEsyTuibEuO3quOWFCy4hIyghk4MQaBxFnLfmiyylrLleJiJhp/rwnPqYYMwwZ1c
ybuVkpe9zsC6Iedp5wLICVvF/l9sSwLFrACZ80R+knhF16/NkxTuDzohkOP36J2rtpyoSjXiMcR4
YgEYWVe5MYQebs2WIbsIKKZh8gQaTmwovy+dkEJaKSxf7SrNJtReT1BbGaJqPh4Nv7uwjYmQw9YA
57j6Nhhck4+vHDCJIu2g8z98PuvS8UE6V2icGNZU2xri/VJWq8sIz2Ju9lUncFMUiYnCOJZv0aHF
TsMMZX0Fl+V0zlCRgL3YdceOb2SKXJQlM+x/m7Ak1JL/C+jJqDeeYaKEg66OpfkEryBniq/6eRWh
OTg7saSHq7krTbAoD8upGzSHktlwkC7418t40FIHYG/bdgr4xNR21s2S2yOC645Mg/+Gr55iQqyl
w9J+y1u9bBJaXQdgRLRD3e/BayiALh6jd9zwVrufCRRRbv6v6fSZcOFFub3aHD+p4oMgOAvSMjkp
xJN7CboBTwhRO55zPkSjC9obDhzicuOP4O3hsrdyQbu1tRppvKYlq6CAk6DDJH9YmmxqEtedljIS
SPo16+kxUTY8owNgCW4eFOU41wtifmcP4xH39YrFMHVLwqpu+BXkOvf1braXrqnNzWbg8e21SzYn
6Ti7+x8i0H1z9p5mNyoJC6bKhnREmLp+8XAJa2IlTfWmEFuW4c2rf3KQDg/+GxWjgbGlQj8rPp02
UwbvzSwWUA/1UUNmXXIoT/kDVtaCs4rg7/LysuwlAd/X+v+DIwK5jBQ3juMYbUZAAxx3EYSdSLnV
kSCiOX7sv8r5OIU90rWqqFTxF4++luBWKG46XF8fkN6z9Cxi2PnamRWIdjE/u9/w1jASWQbwKHkU
Ld1z/F/YlmUDJL5J+8FoZZJ0dUovl3GjL4NPFqEwywqGOX9v8z7lIB9c38h6QFSit/xakxtiBaav
YLaY+ThfzVZRWHDrFTWZo9+B80ovUFW7WMbPN/ImHN02Y9emx/cfUQq5lj8nNFZjUq9vcPCXDKBe
B72phkCn73wohS4XIPXKmqfQ5LVAHhReSMjqsOFzTRHeDcLh6cDsejwR4L17ujwMuHuk58JATnIY
UoOpy+HD7Zxw+cyp3A5i367iJJayh3ctYG+bKFDNervsPmokqFxRXPNOqmieT5QwllwOQkT4lhWq
xKDXq9Bjm/w5qM1XMjb66CDALigGpUfLX0d2RFw4QXG9jU7TBmkh9YG9EF3qqNvTWd6/REtIBmtu
ykxG+VWk2Fzpv7wySdgQU3kOJHIoa2TdnSnAUr3xTqYhD7MQRQmP8OZqpU+dRzHlL2BxYxspJIG9
B79IJ++QH/3v1PRtxng2+tyqOch7boBwtJL/C7M04mBJwGhlaRzLKc5ZXuSoRlHmufqI25/QsGEF
a6qVFaTmI9F9RVxJVElcxWEgkwF+RBtMrmHmGDlmAKXlBIiXbWxsyo2fHHw5vqVWAlMkB9e5urgB
MV0FrJzKs4UtOgMu4M9nKX3Ll0A9fXKSJnmaGz0yfdUCfPRKDyLK0BHz9G7s0NAkJiQEugCouGxv
ync98Zj9IZv5WYLLNfDdKreYBD6O8Fj8wLWZMQMyzOkXhnrPTeMQ0dnUTNs/qvQEbasgPyAswyHZ
W5Cf+ahGuawApFgdxgjJURNb4C4Jf9AZAgAsjqm3f9+LDL0+W2PUZHiLDmmNcoC3AIgaO5lE/aq1
yGH03SMOEaGacQM95SseeHr6UgzvtXxBqwBlXkweCrR3F9IZybXuRupmavitUGPZIK/63n7Amphh
mfaSij4tx2AlTkrhllW5h+uv1T2hh5g4rbeB1CNl5uPBb3J4iPr+/3vYpxXpiIICxgWcDYr5Ifr+
HPCgHTm++5waXzS15lRHjxk7xDC8ozTh01LaJQquF5c/BvSfjYrRSTbGLxPrFlyr0HADuvNwMRMt
oc8Ge00A2FzUGwcLd9/Vle3/hl4bSj9S06ZEcS7Q4zDPXN9tPBCc/J9aX7vFCH0jnk7Nv4cdPNdT
2NtRZgZn9e+lnQGMIB803vnTXgqek7ZZIGzzDTf6ZmJgbyJ+OBYWx2aQhcMCLZuBpd3Vwd46WQ2i
DkK90ynL9gTk3jUVV/NYlNCAvbI5PwQdHzaxksGwwGHylXQZPcX2m8plTL2EqcImGy/oVKu6cJU4
LQ4sHl5HDFJ7bksc+fNWWIxSbwsbV/LZ+pzotBjlrbgsI4+OK1nXu3noHkO7KY3wIu8B/AcL4zPS
i7G7mLQyM+4TVBxzBLQ7QXqTFfz2DTvARYzwHxyJdg6q2c6ioKT4l88VOvD0jPFJDnVLx4OkSvef
UyMGGMIstn/qMptXE5mTrMkB8BRf9YtYu85kbP62h7Ed1gz6mbMWtp9ySxGxzY52h8znPUreLgKz
gUoOS+F6L3uO4WHbj4Sxum/TV+C5VRvUj/Cs4Y6HTt3V3bzDj4DLQqNYBkrx8oP5y4RlwLQhA/t2
8ayPLG0xe98jr3g5Vyr6yhwHbtnM8PXssOGgqUQdXouCFE1ACnB2nwZlbKieLG6opP7mzWGfYfgu
EgEDdWOGf0oWo8wKQijwAT2rvISxYGW3vQMayVHNcrDsQh2GxphZEeePJTpvXB83YWpsai56rOtZ
/K4V1Jpufkz+1ZyJXyiSrp48EAaaLMN/LxgfWx/833cbEht7KXD+vtBlfwKO5OxTdAXlbV00BdHB
PabkQJL3kMPT12R4JT1fPemBTtYD45JXN5B771lOOwDkIotdUAdJKKyGNfluBF+TjG7tMo+gX0e0
/skDAaCUbk6Tdmpu47ZtvOsVtve6IZVfF8uw0qCx2Uw6GfbpIUOfbm2Vg6oe1e7UKYGzFT/N8LTp
P+r3nr6xKuOrni2XHtnJAawnBV+2iPcXWurR6sfc8Qn5sXOyD3tFOaE7dM9C4eyAMfX3yNVwC7v2
Q01VCMyshNt6p3Ly1oiG2BN5W3CjfR22PYJpIIpWlXZSs4HuKp4vYnhtdIhhOqkqva2m0xgOcFfO
uptEFNncq8SNBNIwWD86VQ64womCxQi/jP130wDhVqpPfCFu1CgpUWY8prggT4huWlsPFhxelvGb
A/jzTu0oLB+nwsIbz8T6R+1yMRPM9/BMZIXtCVWcfAy1nTkXHMepCfBoJ0rzrVJZJpoUTJr8vWeC
z/eYwCy4nLAqbwSb2WZDaw6UZ/xnH3gI4Qd1ff85oEe2+P2N6fnIssFr6OIbeBD20awrsiX5Qbbw
EVJc/XbxO3EK25SbeHbIBWbwep3oHIXpNcbZTCTIy2kElwyutuehM2vePtu9KcaUyDCJYqbKK9oU
xb7LFSf3v7P8UZCXMS0yo8uAd2kX2dcxVS0ehvJs8fqemUpdfkm2K953C450K0L+2CPFY1qD8QZJ
Xmm3udq4O+6eReoAL7JEpXu1gFks6uH9jGwbtE1ZAgmM8aSuN8/OGAUiUfaa2Vg0hi8voi428z1g
BRcyj8T7mdmvBiLns9VF+BQaTsPshi2Xn9kEutBvFnrt15ThBKMOnVNSLfOwAQILLoB7PNjBShnO
c2WB3dkLnVp1s9QX623pDGx/sOF4V6ldO9UTxNrvE+Z8cBi0RpYB3bZ5iAfTpTPVu9xxJKkt2l9/
NjNolTujqlPHcNH+/a82WZM4H7L3LVmzQOYGR8AipETLoZiKpktR5dmk/eZ9OgfeYUxovfQEkyuQ
izAKXl++y3VTYltg46yA/xASenHD4dyFxMCEknsc3GubYbucoFixcshPr5jKIdgPlF6GkI228MkY
DpC5N6+MIoblvcRglEWJWcvTK03mEFiH/sw7dRGqrBpVYrT5yb1YwoxO7rGIcrSSJoX7ePCRdVVc
/tLeOx5fYUY2W9ZJW5smo7oHUM1P/83ZnQiDHWK3226yx2GvHANT+vWip/FV8jIuihbOaz2OvkHK
AHdnKV4NdFYs5QQSZmTiKAMMP7d5bAwP2uHbDv+p1UmqUGYJFtuu6VN7xhdLyrMRtHDBNHHuTKlI
ez40PKDgAIfmHc15OaXsE2ANt7lq3YIdeHB18POpnYaY+OGgIkYbpNifh3KN63QGGpJ/s+KdcvR7
DGUvLcraBcBMBFYej3OXUoIt1kLuOHgRsFfWTNpWO6d6ZH1hiPfqYzGyfubCDV2CCPsaASv6XUjV
C0+FVJjhjEbKzBnVi14htyFei2SfhZT8k8QZ/I1q/8VAiimP7R1Y4bQZF/yWRx6A7IdsgiyVYndx
gYdf54bWwkCMExIF3Vu5M8HlsFEOrxO3bek1/WGnBcr+HA4IZppfoZZ5Rk2LHREsuc5Jwe5OdMBT
CFV/ulakHgtbvAOO6m/ai915BabvEzkQkPQmYuw4JhVCEJZadY6aPlXUP03PMvLM8xYeyaeEaFca
O7z5hU1D+S7JPaMuYO5nVa6AIpALQSapVbVNhIbWEELoKQ5Oh98dMKK+GBYrxTrr7j4yDVhlrxfE
ZWdKtGukJwe+21wHrruuaXk0GU4rAMBXfqOPlyCFr7i7nto5qmWHiwuo8atWPyH7BA82Flbh6TEJ
0Sljl9/J7jZlXPr/i32kMRe78gJ2DHRs8O6yAka9Zct3/ju0S2jD0xXq/6qQygPVImydEFCDRnF6
jUjB2e9GHvt3Mwmp65k9XyW8GfOEiRr7rRTX37Qh5j3WFbVJ7DKpt/Er7RBxcCErJ1KzUxaPs7FE
MbmIgBmgqD/u6afcMz3ZZDo5nw5ygfUvodHXtX4UYkHkPsXyMMLbFMA+cNYsf43Q7hhzIUsP85kJ
Ju1JmcTxGFAJ0e11BBcgvwWbOdmTLPq+8t33c21uUq7h0IGK8943N9X/r+uenc1998lygDzyLY5Z
33LAEmjMtKTaKthRw/4euFvBhEukZsNoHR8JEh+AA0p5a93pghJC3+OykFDDL3UMxmXUmWxrW4xy
m2I5k6FYbumoHaNJA6pkpZq5r0L9fSV2vl4PkmMCdjKDpiijJumYj6SiVPV0H5txFfEYdusuA9MR
gRA6ITpqA9b+z3YwLCETmLnGTDarrRSyxvDa2FmBmLXxhlumVqVvgbfdNr8D3TMqr3clexsuKRp/
ZIbAC7Hg7/EWSuVY+oDXNN4+1N2/D7dOT90R1884aq4i6NFFI90AKWP1YhkoxzBw3FasGy2OkVy5
0eQMRvofekRUlhf495PeBhaHepnSqnsI2enKEp8GG0mguiSP5hJwQ+cHoTZZ02W4VQmR0g3BQwXw
jsJn/EkfpTw0oyKGmtT52PBQ6WfpaaazkIEq5xxHMQKVNz3pgDs8dhAXDOLm81Umtg5XyppJVqPH
B2jReiJo6vCtbJe4OfUMpHgNTsBZApzoPNQaCYPvWMupKMjYGg2EdzQMcq9QTg3CSp16yLMTyIUr
Pr/ySihqKvIrt6+YDcn4rhh1+/Zm01BrY4aD0C5aW7FOiXehrTMnM3rjp4uf+IJifqJ8TKlkEzwH
dus/TYRY4/iPOPpSQLJRi1Qt/V09BRHUKCYZx7itulOre46ZEf61ZcsGEl1T+jq7MekwXTd7l+cD
lxG11ZyfHCVah3pAk3egg9RfA0qLw1Wz+1DJrRC0QG5eR+rlvb+x8eBrct7+puJLAG7EAc4g9tls
aovdZNhJk4yeGNUuv8wpVuswkpiwktPcsYIEF+slWcQ118NhLMEzQjGPsuygyJckK79m7kONDt0y
XCU7R3ov1YiPqxWkH3cIf20fW6mRVLNJhF/815mbRCbqxQmCOVVikJZEzknMNzG1D+DnnWrmVvhE
jy07gKAm1xvgTMCCmf6Nm/GAZA/2cLevs0sohg2RcX4bA2uy6TGoUYN5LUDc2zxpnk1bH3kRwctO
xaZDN4SF1YjS5p9Xxa9x6P3YWyqtll2BAIo9Uy4GVyFZoQ6ci9adLr1ON61gxwQ83LeeSsl27L8U
dcGPrzYXjTaOXS7Ys+d0gxmMbwaAcii168uDkt6c4zEuRGtOov97Q8YH6lMp82flLUldczbCfZw4
LcH4m2Wz2wnT9mUYNMxyAAMUVniRE28sgmb4o6iaXCv1/tJBzf+nMdwlaZek3j99zbf4khXfwloK
+fvMPyHukJ4kaG6Qfi223OU2VVX9lcD1vbsHPzL/jZ90DKbQYuIGYRyeYjMzp3Y2KQMJbYlwihl2
VsIruvZUZLkuJ5CKfZkqksiITslfYRVNxtG+6TJ0lQo0csUb0LYyFPLG3mFfSeu6n70M3B4j96QO
r1XAr552j98LdLUpZYBEq/g2pz1TOKp8qEoGvYq0Ab0pxX68Qqj28j8q2EEIj2+JuQEx8R0vTA2J
nDtUJHGvPigCl0korn6cziV8k08TK+KzYL38hAbrBn5w0UHDbupDl0jCt9hUt9HPPNLXQ4zaVM0N
vGAdYkFwQwNzvpWplMEu4iBUqzw1n0MxFhGBxc4tviQOaASnbCWfXlnjJq1pua5STXhLQlcxDlvb
aQc6yz4/ZN1KV898FVg7QwggayST7x1oe4k4rNoHfNtVX5ZeTW3EUVsXIucoCKpBjJuNCm4+OwuU
nrLJJih4WR+f42sAecnvQad4euowKzAdna/Cntdfq95+VzXFKMcCZKLp6ugTw/ahw41iFwoiDGSF
7VRcsaZ59nQfQHRKnsrhF9GNScdW47JvYKBEAwDPA/RAdXB/7Cx+nicVK59Irh6daV74NFMpKjOm
twd5XurRKcUnXbUuk98WVXEkBRsucFAFbm2AuLGzysMAhA4PD0av1yhSHDwBNMdvheo4wYkDSHmp
BnKBupgFZJ9o7j/4cpxPPALe28a/WJ83PDIiV8PU0pYhfOPyqVzzNmXQnuhil3BG/2REgHDxbYRX
Nwyqw0WxjOn7wHe0mNLloHO1b9RLzxcpI96JxFyhWwfNVLofNFa37RkGi6Qm2p0ywdIaSZWkyRIX
SOFXveDEMs7kNeAr5OPFNfMubBJV85gYNGERV8Xwpj0VMbP98hC2sAdeFuyqCD6oK5LuDU6Uv0KV
Sg8JQw39/G1nAdYFC+25fAL5Ph3Od+Tdrjtrf3el7U1eCo6n1qfnIxbbWSMauEkIpd2YalHLfNXd
fKtZ4al1mYXEcqXMt+hge394vvGYR/i+Yhmy0XmtOBAeN7yFmzlqp6GVS/ZkrSccQpshQZy2CzDm
Zw16RNhu42UlY9uGFnKaM8zQetZc/8Lh5IRYdyVbCpYzCkZeXNIjNJu5uMWlKJhwMCIPxkUwWtDT
ifgLXglVDDJgCbG9YQ63zHYqvwvLLro809nxy4KFkD+9yQF9MCib2EQ/OY7m7IeecJAAQIlvlWcn
JG4Q4OtXvxD/aCqQpRP+KMLI7/X1fJWo0Tzajhdqx3FfV0nMbN5zAUs2o8dAzgOPuf47oOdJFCtU
olTYlrDaARvImhvwkgTIg7l73PcXkIJNIYf0ZiaPSsjn5kNTZHOodzMQl1xCy3dP0DKLeQ4helqJ
bUsVSpLceT1YdcpgxVqYXVte0cCGlfKnlKM8SMQEYnSzcWz2bpu1NSsgDt83H5uLKHvbc1Q2oX1w
MSkX2Dux7KuSYuLV36eu2GmL4Ow314isMyPt8oMeE6DzyyxvJf8V6xCEmQyf6/8jrSJYxnThUBzX
nasArcMgw5Q1sOwq0Y1nhQ0VC9Z5ATqCXVHpwNJ5/FsisEFVr0WC5dtHzj5iZFavM9mnvX28kviD
kUbJRfb9WpebkwEFbQ0npWxTrK3WM8lMa2Z6VdLdcLSeGGrWUVNFHVbDR0AyZMlpVV+QRyDkoZDl
wTMTVUc1zhCNdWgxSLtw1Wx0MpAitB9Im2QPb2V9U0jUVpaOLEi39zFInXze7GD4IDG9gpk7ep6u
Al55dRRWX29qcSGqBuncW4WqgfLpxpGcuRtg0yCOEM6cRZgkk+rHx0v+Egh8ZTKrESC+AB49DRT/
+3HZ1icEwC/2kDa6/fal/oYFVU+DaMtDrgEWEslMcWStBzaZj68DcLSdKJJCg9g/0gy2F5O5y7wo
p6mc1pf5igxT6bLpLZsyiEEsJ9OioEK2DJTbGI++P4ImyB2sfoIjoH7a7t8w0jFnkawqKIFM7fQ6
xVXLepSn98spQg/tvcS/SIwdU75RKgbbP3pXspGCWSXtsyZh5z0oagd4aSE29zIPpw/yc57KPZCz
5bwaA6UFMDEFAR5ZSUfVU8OcT01kdrsbo0KpFvKsF7KgvmWjWp6tuA7M90I+4luttEriLVSA6rwB
Ck4OpHd+VxBgQ5tSFqgqvSfHQAdPvNeyChFhKkrpPkJqBwINL4wZCLjUF68obve7SrBoUK+zpuMw
N+ED6iH8aAaRafr9dWa5Wuh96uNba8vQEVormccXOFmZcrEOcNqycZzlfdQWicDdi00N4RQ4Bw6q
rO9FFuaLW4DmxXJMngm0ZAfVSG5yt+YVyFbguIkdw+CQV4XmiGHRpHggzNl2wnmQI1rS2vQKXE3/
EbkHA3akeVdsK+jWB1IFGxgXAI28VsfGmuQfknSL2QLTL68DO5cjgneXRHP+1l7sX7bfq1EVWM6J
hU73S40tC78uQgJ4ag1VVyLpU9PwqlnmfE/jv8zKFjVVO6E5Rdc4BaSb9+0tFNK2ttLOOKf6itIy
08qEGfb9qd/Ul2nXFIWj1hOmfAZfXlZ9kfL25vtjAN6sAPWA5SuAFJhMxqgazjQVrDxwgiPEoFwD
oGQf86zFBIjsSd2N0da5ScxLg6KLOdUdE+c1tI+zyxcK2H2lnGEL/LMx+BxCRaQLRkoOIx3H7Ddy
on5sVXsWXouzeN2RZZtre/rgBV7Rj7T+PTY4eiJ9JaCrQPrfDiZVWalPIL8XM6K1loKSMca7Lf3P
v2ZlbJMKuXgFaCBaSCkpq1wBS2Qz8ErrFK9p/HtP6lD35ZeOw1WxpYdHw/mQZ4dwj6rwyjgJacDn
Z0EGQbXRPO4uW/bjsetDgWliCsBv3HlryoBRYeHqf1eVBTY1Eryi/GJwdvHwJlBkc1JK6iqdUt1O
ZHj1B/t3q+hioJ0x9jYWckyp8UqWQGxtOixSc4d0/Bni8TwNu4XvqZm6KIzwC7ayIZdr1IeBtDxU
JyO6XkWTsDuocQ+padg58A1cgX4SRIsHzGQrlkzOB4jWt+yd+lxYCXkkCkb2lWuda7wV2HsGhH2w
9zNkgGD7b0gozRPW6mbXe9NNFjSXDiWAdTtcSwuKyyAzLgTyf4Q6+1CKBNufFN6wi1nXrrhddwbk
bbh8h5Fwbv4PVDzNncj19KG/FZIFgRwkkB9dt3O2g9Lz44rFBU+NGksiclu8ARChiWuL1DZ3TWXb
24G8CEI2hXJDm8dCN4yiFyr4IQVqUNMQqw36SxO5zDhRry6xJYTF+HNw/51EpFa0p5otPyQXYpqh
LqkJjReGDXsbQSLWVo32Pjiy5jD9flmh6j5eQM+5T46OsJjkgL7YCGOAsPQt4qW/B7WAUOScXC+F
d3EbRO0mFAQqJPvrfDyb3SSDsBKSF3IJf/r4a/6qvNgjTrkezMn1Gs86WkqFPUw/BHJGFbCgZYy5
ewG09vmsKAdGMwU29vhHriuzEIi6fur2xHKarxNSFlF698qEJYmx01YNZCv+iA36ZR1VB3AHQ6xN
j0L9WFIW8QJY5wReDs2O6EMZ2cIpPknBwDI4mJSxjA+X6XDH6dFw0OhOwB+K86s6SPH+CGmKaCYY
Hg4LJMu8US+Po5kiGPR6MHEknuMEFOJGPkLhJy214AmGdv1Uq8YDGZ60e/6Y78m9R/1G7b1fdeFx
5ro6bhkoFAJ2ZMhtsl+Vjhq5r9AJ8EzBY/RVlgnKwOVrijthT1bm2UKu3T+qRbrz51KBzYkRkU4E
Qex0b7I5AJaUBk7UUHHx3vB0sJv8z42nJr3pvKSU8XU8+p3zIWB8i7AJLyj3KAyfaHhtR8Z/xbDH
vmsPrF4l5XEaizGkDsL7W+enMNvvzx7XOzxbK4YjldfcSyidjhsDVSif6M27pO7PbFsbWBuFR3UJ
U+fGEpvOLMJfE+kQ5LRxVZ1qO3XIfoSSFHsUawyUPhblMrNDhVko3F7H5CN41Df/Z+7RWlqy/zZy
GvmKPFIYmz5Rx5fCIfUQZ3pJuxkJEwHOWKVLhAz++3523bpB6X8m5wj6XWXEf0WLJBiDyKDv0cWP
G/KyFeJL6XEOlj8uO1aw4rg5ggheDRwmvnOw0wOq8cOOxczWCwgvAFInGC3dOM4DhlibRHGJs5EE
fP5KgKQpeabcPQSCtTa1iWvr/cqm425jLgbeeL94ddPBVBytYsfVy94EoFH4s5TSNYaO8hSzb4O3
2i4qiO/eshodftfC0+cY/ahELY9a+HJAjgAhgXe/eCI1AHgznSHhCoBZECGuSx5sWnJOdsBX3GKP
JBO2+LsnKe3lXz/iLCrwmhqVraCHzDNWMFo9xqpzhfQ+NCh2jcxVVR+w7INxh/EkeU1ymvhf0bOR
/T6DtucDf/YFq4R8HACMpdvA97ia6afH4sDlFfG1mBbdvhpzmNrS7S/r5gMzJG02OeDVkzsEi+v9
XtqFMpRzVknGggbeMzk/LWt3VR7tHu/yJVmA7jVxy7MwgxnwHdOPCziXmx4609QOugWhop+SdV/I
WFaeiKqC5UuYdcr4A8wTsoTrY7NpI0PDi+NagBPwtNgg+6p7tcZsaK3fLM5EFg+npDe1UhrsLwNm
fbXfR+8VjnCrIJle8E1L55ZysuhVACs8TR7aLUdwrwHwg15RONsDSs+ZpPed+PY+k4ZiGzl3BZqy
KqGoh3/O/B05h0KDS2xu9fX35HOP4SLecivDJBuHGyGKpj7gTSumoP3/JXaZzK6H51UzMgk6F5BU
Z0UpW1lUx+CdcuoHmH+BK02iHrzFG2gx0p3UDepr/t/5G/EQVKPw+gYCWJ4ybTUIjS2o8B3VfI+u
9VhA4HWelKiNKACJhaj+DgDrQFtszrR+Hk0JirNF5fSSwbak205/aUBHN1Steed1wMGv4+fyzP6v
Vw2WpzhXqicWThgrunmjUq28+dp4o+hPL10ANLYIJVpz7w9+a2syT59KpDGFJnfI3CMEToklALKx
bUSmpeN735vr4BQ9jEiZyZJdr5LklyasdYVDFOd2AfwC8rbCFN+xaaIZmRH6mlwXR5wfUZXkbSd+
4eDObM3bSZYqWCfPZ7pyb9xKDSdO0bSLEqt/9EEtfm52SkNU8ihG4k+bctQV+2mJkMpZ0UxNhncS
9gMRpfYyKyEOjFaH4cqd+oQyheB7FEcBjJ9WSSw+m0GdiDv3RLyqnl8lc3TvpodXIS/S8CMIJv83
Kw8/iBRlC+RkXPfbY40qHva/miW5al2ucF6nAJ3y17XdVXIsxXMCsdDpQ0Var60Vke9CcT9stjeL
wzJ4bOxDEPo3K+7ZW0XmUTBQiAVCv3AGXZ8Yh7s1Vm+aGlpVjAC19/8ZP2RBHd8+pNxHxq4mODCE
WOjryN5QcZbJD+FzLic37pJP3z6MZKgLUEns1QmBug7qUarHEZbzPvX9HZWK8rQ0PTYlN8TG4xq5
iwCh9bG8jYF1cw4a19T+MFp6JmO2xmXzW2kx1XgoRW8wkU+E7fOaK3uPQSgKKHboqC2lwd7OPB8Y
JpEDAj10ai4MYwo1XkA2b5s8tB6ucb1CpsxsQAdzBs7fwHYKgXqPPT4jfoPJGTNQYAZVd19DhNQ3
zq0Qp5a/v55eDXEk2+zPOGGIxLmNK9SDYriBC3mLYRIy9UNhIJ9x74asApr3htzTLSm+EhgjHgdV
0PulB0osrXjJZhIU2l6Mp3Q8a2JRq/+1nKhREPHuxo+XO0MpaHp8bkX7CTXDBiodKJMgabm2iEVU
152wn38t4rjpb/R3Vp+wU3ntbgzC0kJ0Hg6cQaWxY2AjSlHKiM6sj1/0XhxLdU02qknlKtk4iPhh
0iUZwwv3jpTOswjyQ3nJaUzr2WkcjqRaqAOunGBuLRAXT0moeZ2tr313E2plZV4ynSKr/9Ne2bgX
saknz8z4iqOg6TUAmNjyV7PlO0UHTZtgFnwovlb/0eb5NOOyk2Q6YgUpbl7D8bRy1ugoPFYQZgVu
kM8BZk1BBtqe4ZuOugerlfnKwPYcFCbBc5fdYUeKdpqkXGFJpKNB6agBWMx6DqLwNJ5JG710esto
gjJ4ArzWbxhEdHaGm37bUlhY06uJoPfIhrn+BJdzSJvlf8ClR2ujeCjLySWJiNTKPdgVZSs3iLEs
P2pDMfEVNSs3kxkaJAemm5FzeGKsPywWBy8NEAS97CG6chfipoMAYXMLLhRiut9nz0UrtOmn+Rcq
6gm7Djuwv0N1eHjtr34fKJ6eryPK9hu6B1KsSNcfQKpuIrMS74t7U8aDrfJI90NvXiuK9wEtG2hA
JpvOq2BFC5w3fZla2xU7kJC/6uUDisE8k0tlqvkMXaOPFo4zRiOtF2WxQLzY0G7U28/7Je0Eg2ZK
bZA8ofejAXsM8mhKiYUtrLrQuHbAQxIJTgz+KyI9qn1s+mBfKe7fwaoa44Ra4fE6Pn1q/XuTyq3Q
xRpTfMsjLTVsDar9evmt73MmBDjwINX/2Ttus+Psns2qmUV80bxQYZmUbNndFjbYqg2ITFl+4bCj
M8QWJEAuvjLEd2hPPiQMcbuq4R4t9XhtRs3vMB3RCvraYXvg3czOzfpA1PHwTbEDA65kULj6A0a8
E/5EbdVKW/I24zlDjwqhJ5yhl70ZHSpeYW2e7fqcO8oBxWm3YNQeDHRBjVq6i5XaTdVJuoUS1Yzs
eFUJ0/LwXjiSrkfFOY/mhXtOMLn2b/bSSH373TFVwGxN6rriKp1z5USL+5PnQgATifRgDMyKF7n2
BiEXFGVe4qx8c0ItzD0sftWwWHnE3S/egLrVApvoCT+NSB/rGu9W00OBa4OtMCaPP4Emd74mhtk5
vY5lFn69JAS47euRJNY6mrPr5ZVw7RvgpQjpqZWDMXXOj9oFCpUMcZZNUUqLmOwPTuo1/EnpD6Pb
3u9AXhR4iGTUitOUxc4T6/eQz1uGudT8foJkD3P5RKa8E5+h5IAnInrcQCvr4mc4LAUqT3oAddEn
Pp/tgysQS1Ly6cqqMgLtn9sux8iuu1n0N2S1RSD78He2udHwWCbOdg3n4N9OsS43jia4jKHHoE7z
xY0l5/NHxY4HeZRgIVZnIVwcOphvjM3dlrg+Rfxseb/GijqYhuse0b+lyYhURG0G8o50HBaIi4/g
gFGk9rT3A0RbawNsrKEmhfP3xDQ5FaiKbYtzHSLoa6oiD+l+SLWCzISFtfoMSofbdi1e3tXIgNtd
8eRL8/JCpaZa54M7Dzmu/MiVCu2V4/MaVF45UOeF2qTSrZu1rnRpxG3O+2lEtZZAKMg0ouxe1RSj
A+k2sFfdItnlobar1eKSmMxnpDI2BCR0KLPOz1J8IiiNnAPk2sar+H2BbsY+KV+9Td9eEna9nY/X
E/58FO5kP6H7ydKWPHy7BfGRxbvgRAptypjAkgJStedfFdph9NGN2ymqsTF0Vc2/ATmgRMg8sx0t
9ZpuC/aqXLGz8Qvgv5CYn7lqQye42ekLR0iZnhyqc3V57MfTelgbQREZEmTtkauIOSRETtvE+FJD
nIBFN2+6MGodO8Jte4b6StKZCuBiQZCHizqMfJsHiA9E8VXlUmGnoBJ4vDkSenjeosTR2i06LwdI
il0LXXtp0xsDEHJVUt4mskDcN3bpfFzHTFLrduyOCaYCm8COWs9vo0EmFQJAas+0Mse2NCOCy/1O
2NFVo0DxOvvUf77QzS9TKGTin8UkJtDuo74R+74II6bfjrVWJNRxqVjxFgkXweSyFSgCltQFP1On
k/gHgirZm/qCGQkmr3VVOKMXiniOlnnDFwacjUAuf7ufuKKEnN2Ke38RwKQhLK/tRJ7Sd4XxwXci
8wRjlZraVwzjTEvLtSPKcSGZtcFpQ8ZAMt3NX2gkY4dlfIsJSYcKzQaywhonYCQ0q4vPVFXIwV4n
VfOpfJxuuIJ7SYzzbquDx6hdnn88Rzgly3cF2A6TGXUHLqWkAHJWYw21Y8uIzZQ6zZHUThtZKJCo
rTY1lQCBQtxkDS9fN/RPAgwKON4IIG0Nr5RtB1ij8gQ+lDm2fFt2cr3dHSvXv47MCwxFuohlONyn
0Z8od4lUayI+uo+WbWo0G/+R6n241tkuVxfFL0qqvGprSpw82/N4aXn0ab7ES6/syXqJWuZ+78jb
iN87pYhDtDGI+I74acDNlMJ4oe4cqK4kT0ShDn40v86TvL2cdnB/1bSBSifOhlOie4pL5Xs7PrGq
EsqgkjVMU4KD7kehNwisYKnJQmSaCNZEp87rLR2uOs6TzzhePWfp6BMMbNLYqw51PtlIDDKdyD9g
gm7iXmpSfwE8tT9kURUJSLiD3p+Z5LNm3EsGGTngJUVQvrmCDHn06LWiJ4GpD8tBmROu7d9VXPtX
LzI8ckcyc0NF/KM8mbkfUuZT9XniBuFak5p7dvQOV54G4PVkvBDfLGVjRhZuWllQmNno5S7jVNCe
ciYUH1cPZ5byEJ3feR+XgZb44jRRzizZ8or+gGMLPsjDLBeQrhDnoRnYVx9QYEeu6Mi+Ci5WwhNv
UVHmyOLleDfhJGIAU9DLOGjCyp5PQFZNkZ0N/nGbr6dT6Ue1lQWUfxZSdN0qg5G30nd2ezLZoH8x
jnPcjromxr9NhZWVaxL+YXcE9N28OxWxIfjI5uvVEdCtXFwsa68ndnM0JBODDFmM8uY4ySNOQPiO
iK49wyIlu1qdRaoLsI22fHHnOMzskomKnfoS+KiJzDLf/xLKjIx07F0yVKKULpcQAMDigpejPzR1
+tXV6GxiB+79TdT+cgh4NmCPJewtrdByMCssMZvKiIkhCT3LElFYbE37Xieo3QVsyFduXBo5biqG
b0x3SXFg+n6JWvWkiTjaNEAsAhrTvFj6+2ulmrka4yhOOX3vm3Bwp6phjpO4ZzvieRiwE5ouFquy
Fu+rtkJWEOFOBWPx29N5xwXd8YEIZjM7/991W9ZeS1U8V9FywBru3WI2+Veh1IyBsSqbM97zg2YD
UhJddBcex34ibsuZhNQEyWgc1nTSHi+wVuzFLWgf1FZEp1usMUDElU3TyQGDWu466uY8RsW5M1Oh
cGhouChfCqMvekPzq9gN1zZdTmCU6oFwDDw27u2N8inhsYls2yr9Gy5NLJxrlfCw1SNQR7q45wLl
+ioJ5rCB/Vehtyj/OzIuZD2AliNHNKRhoF4hgwxPwRZmsGpPsI3Wy3o7ko7RnvhJRd+2JXqMHSzn
PCZS4KkbjXNEjuWSfqyPUHUtpV8fOOXUmfSLijf5xpFYo7pFGM1UG02u7SnAOabslosmYNVfotq0
PYvOjFjz28TmZAAMGZywPsBRRZhyHPSV0pHUgAKCC6CoeY3U7LgpIl8ctdSurFOPRfnggCBEFjuB
Ho3cGirY4pzDhXSXI1M5sJ6S3bVdgOpY9GM/2K4XSAHFNn/6ovDIBAh4z7Yo+k4fqbsFj2+cfp8l
AFeykwuUa9BpUL+UJ442f51rdY7lSek+hhV6DBfi+tlzHye698gdBssa6zDaMQM0yFzlqSNcmL+V
ffUXA7YDwAVYYJCeSbgfSZh74A7iSQAMeoP4gRXyLG5g5SJVCEa9trqCijfNlkdGqjFOY1EGXuFW
/eOkS++EU7LTzuxbdas0kgmcJi4v94cXYj90fVRdAY2uAf9BP2Hd8FOOlbLmFNN4Y/PPGSksc9MA
5XRQtMkgBr6aFvdduwZK3Klm8qizwyS5NW9IlvsaSGXDflUt0yAOpe9+eKSHxW4o3FFrfN+hqvz8
I51UXW88pvlXoAZDHUc6yagNTSCJIOZcnVKmiUtppVpmiBb8oBHpUaxKRPwhY/qNR47NXrRzlr8i
SjTNAZZxtRRro+1n2azaAy5ps48SMq9hRULwNQKh5TM9LD0DN9qXo+qcjkewqlssYBWQ9ZYwAlq5
Dgo/VEjT/XLb+BMjV+yZKhw+DaJ79GkJ7GLoV5aGTKU/Jy3pD4BE88mLgcKsa9N8TBQdLE+WjinR
6R2JqlpCfa0WRiXRIuURklppq18DaRAt9vU0s71I6S93AVi1OkCntshNSn9bmNy9ERtgcVFGdvS9
SlgXfcqLWVWTZcvvqjE++HGMrGgQ4EKuCmNa3Gdk2eL/nq/iCTob9zY8XNWG72810MVMJsFzaNL5
leKfNi7S1q/qWDCT+t7a/f/mugfHjyNfR/GbQpiRPAHFykB1POsq9Ux8FyM/y5UVkSyPUfiJK01d
5EEE9y4TRZhGvq2xYfwTp0avZgFui7c7OJj32g5VQ46CmgFjdLgqlPxjFby7ylU1adoh+GGplUR2
e7q6zxe7CEfFTbykjKVAGNCY+M/P+NZ3KSNwdfUXH18Hn5frkpsvrgQMCd1I+zfRRqFYToSnPlhP
7NRo4baApGC0SvZZ30oxDzIT7fGFlZgJeZq4j728c/q/HCmG3Xmmzt14Q+24FGARdJNgAYrnyH5e
7ZmjFMweDkspCfcRGmY78g/T7jehLS2xQtsRjVUNoeUQBfz6ds85Sv8bLnr2FOl/opP1YOEi5Bxr
rouTstl+kicNYb/UxWlqDowPujLi5i4uH37n2F7FhXmdjrJaUtWajTML6WvpDqI4lR3jQcYXUiAJ
0v9M2aPcDCyWUdjPvi3qtOj0/CwE4Wz2a9vGCOmdfBtWNpQJcqsl47FyrH/SRORg/2WFDix0o5x7
PBbOJQnOCAvl0KbHkf+TmxCqHCLOMie+0TGe0qNH6z4PPzG+NNm7nQdvp5zOeqeOkh/1Ewyx9XFM
lYqajSZjiIaNCTipQ5zH0fmRef8ysv4Z9K8R1EmdJRvpsCD1nAXywKN6mkArdC8M7M/ll+GEWA3N
k4CdQPULpI7+pdM7JSvoE/By/2c74ZFnkGOrx1IT1n9z/PEtH3o3uaQuHUbLlTi7pHsrIGZqQl/a
X4l72ZnDxjxvYHwFHUCyF6CPDwC7/V+IDzd9lBBX7CNDY7TQamkMjhumICnAFNiQMg4q74GR53iE
XKbxfSNSRMvtVsjWj4s7Esomi1wtjzKsPM3qfEhlhzSumsF7T+KH0cN3BmAlbGEUfjFKa+ZjEyzD
GOLufWKAI87ewjpBghgE2bZIca9tUF8UgY25/aAHTDpZWCI8Li7yZGvOHL1SBgvHlC1GsKymXP8l
ZuiXG3mZC++FmYt8hCxqwkZXL8CCtpbaOokHmSE8aJyHO/rwf1H9u0pKYvsffADVXn9yo6EDtVw/
e/Su90tdY4gCY1gnpRbdWq1AqkPHfx9ALkKUTH5WjlQ2vWV/stanmZubaoKXb8h6Kelh/dxjeRnp
9ZcKOymm/aFKhuUioDGKcxTHohiWUyUW2sEmbWPRWEfDyHODoWYWJaeNmOp0SkivAL2+IDBN3dej
3vTODDvzzVRA93cb0rzBL8Eedq38AL8ugPszAvJRHLwLzrJ8ze8vQuGwC2ODfc90V+77W62vwoT6
rEneFqyzTcKk9eNMQsVtEst7RDEo2CGTBaf7jb9wGrNo/EIjaiD70znjqU6ERFU80HOTJbR6eM3r
NOIWt4yLy3LUtkdZoFzhkDu3dcfMi1X5zFdTqrz8e3rt7/Ykj1kethyz7nQbrg2MOdJSumZOJ1Vh
Hf9eO8p5IaS4ZKzxEWFR8ciGW4no+IaRmYnJsqshRrrePsLHuTjK2XcXdyfJ5bOrUUepnTBgycHn
AMZOlR1/PaPQMTLneJlhYkEDt0CnocmodrIs3gJdYpP9UGmjyLpEaoYwaH5LAgJBahQecdlEX/ao
LSsjn4z5gG8whDrrKvGEEbEOjhKfXJrAR9DpYf3w0NlXTt/yMaqu1B9a24muN3r4JotjlOXSLH22
oQlaCNXw/TRnz3WeOQCaa5/jLo9JfUjw3SPii15/PKqiBxhgGpkx4Y7yW9h0/KVIpJmMNnlu89wi
gBWoE76JIckvirWwp52nfVTjazx0zCU7TzbazfI6vSrdNcTRaAhbIuqal98EXRO3yE3MILsCf8ME
mQJ260UWaxuVBzlIsUeswhdPfDWIIEIBwNBQE2M2cMW6wSrGzpFxBdGp8AXREgktkAwu5i0JMSQR
lpiUj9Wdn/wrA2jZ5F+VFn2YyIYAbze8psMpVrxLnfB1XXn5xfjQEt2cu6aZUxipLTmo5WUlQSX1
tczZ1dyqnANYovu6w/zq6Us0M5oNAZSF5Vz1OvWi6Idhn6QQYIYWN56hP+YQj9oO0zW2hOO2z+zN
DhtUGhQk4uh4bsh9tPDvZaviFzDoxcxbDtWzKUddanAJZbFDsGvueG7WknTV3tg3tpHEn5poe+7K
QAEUZnPatHo5Chp6vAQf7Wg8OVe8Tjw/wKVKnCmrUC32zBkS4in130j7UkQ8ZgIn0MU3VmUMll8X
wuL0JqcnDSr4O3kD0M0+DtntSqRpz64/trAPz1hzAGYbfBR0ai3S6EiQGQY8Y2SNPFeamuRr6nas
COAinLE7QbmXpcXss+AAU4cqo9uMQCXYyRDAvtYuBnUPVNoQFWlpBoE7LVjhByzrTB63DTgHHe6w
xfgNzmXllRkCObUvbgxGKSURxoc8T/QuVEZNo7BG/Vu1KZm4D/6yqSE3/e18reF9ujyEP6H/h/zu
Bbo7Z1FgkZ1I9oDnGVvLgrbJqVnbj2/7eXrVVcuIVOZUHyTiem7vuQXa5y4Deqf/KHVR58X/zVq7
KzKBdHo0KXl1nkUTi46EZUIMk0IJ/qdyI+FwMdQ95Fza/hs2Qa1kzBhtcKZqzPyO4MRc+neNUOK8
7QRKrZUuro1nhL4IRmmIXEYCQ+et6A4vR5pFtBKdxdsmT5BNGVyPhzZJZxpuiA1vUODrdwQUdkjH
ooPAmTpnvlSwOuXuZGgsehESGU7ExcZGxVzyu6A9VdUG5O3KOJaEb3zITGH+2nZj/9pqJGEzMBS6
+oYr+NhlcnHH0Os0ThKVvXtoq0te2dZJoydA/YcUZ+mNKF1ZWwAsw0s27HoT7WDXb6qYaIeeTxCU
wSugbse8wGfA96gSRTmFo6A59pLu4kek5uaN8YOvOybgIFIpiHbKAJ+6DVfE4WBcdsZizRWgXiMx
WV7FuUfmpvxedceI0KoSHTZktQK2GPkNfdJht7brSOUuJ0+lgE8+FRm4gaHZF4I4S71uvKfLxveu
+xIXp0vtDFw6C0SGSLCZ2JGxsos652MkpXphrmpZFPXfbrMUl+DudGVdHX48IH+nxiUZ8LJ253tR
2L3CcbmOoNeQutKejCCm0oKUIeFqcS8pSP98AQcP8Ds9+nZFrwr/nJ1a40UXd690jv3JKAtE+WcY
kEYZLmdgyNhuuRM9GO+JweL4hk2CIVDmMFSDRM6qCeQ8tQvbxq0hb/IJvFtc9zFVe8MSgF+1kmSr
spGTt2BB7Ca4WmP3wcXTVyBmnvoWbTDX6p1d4a59+jQe+w+1263pBSlwJwf3ThrW/QMzVEKhH8w+
L4yrVAhIxKywD9Uw5HWTB2r85Bh3kGiQq6/AGJfSVf3CVsi04STd/L8c+4chfhLuD9ch0FQldcZQ
S2JIUmqdhiRhKmUIiZTaTuZlHIWGfD0hVi5xLt8rUor71K/cPnpxgPGpOI0sTJ4JRLb5+qJEekfV
0Ghj7W1aET+DNCMlQymflcCAbVItAB2jS4sQtzMX4t583hgDP8qThAf2EvxEDo2CTFe1gqD4wEbe
O4JbDuWeFVjn36pZR/IVWt8+h9TgHPe88ItU2d9IWXD2L+U/xCm59MeYxBVjDl9jKfL98Ur4QD7J
qJwJ/vssaETVEfXGW9fKe3d0ACgxvYZvrgi/1cVoZ9NjR47HC23GogJifBdSJeHnaKSNE5yLoLjJ
ErwP+BMSNqgbP5IS1avtjbU0Nhwmo7jHkr8QVT59xt2a6dLk/KfbDWcYcT4sNG0+dVqZApF2OduW
AiYf58QK5ztAy3pE11RvDLKD1fZli5UufWgtlbkBqi7v2BfXGtwVu+d+7udog4eFw/UowkQ0Ff3H
ddzsmJ2HKvRVjuhmWhTmn9y/ceOQahtez4gbN44/91tgxNzj9jhmvijyGUhSStlkoCN/8FjDjoGk
k3Px1x8YkLjyRVYyezk7lmZcmHaTlvlwPOWWUOKT1awPLqcLSovIPW4qTcxg2clXuHL2lOr2hfRr
dtm2ep6fBjNQMRQLEYcCuYK2Bi9EXEE7S4h8CBTf72ypnKTf+ScYp5YzxLw3H4iOyB+jVVa5F/Hy
Kh7MqoSnF8ufoC6enl04jw57d7LuiSxOfuf7rYxa3RvqdjHf9B8k/1K0bjvz6xf5f8H/CVq3I2iw
L/0XmOy3dFcWop9s94oPZPT6mvVBQBOJ221SOYe0Jw3MxzwSb3UNc8Sr2vhNd0+KWoDFPjngErjQ
nbJsTXc2Wosw1NoiVyNs8pT29r8IrGIW4feqotjaJQo424GqZky/pz63li76jwk1XG5HuQPcOrIW
PtkpTt8NFoU1sdXCPAYVT8kIe8MeT2j+nfclAl1SV0cVIOzvFpLMkvIDfLBag3U0wNubRNxA0faW
u64yL2hXObehrWYrfDugdWd8AZPbjUby41NQhzXdNopauW81TWNLDvUdCZc4peS2Z6QNPR/axS/r
cf2xFy/MxvZjw70KkPIqIEjM77JacHa9fYouJeqyZv/cPCoc7cXZ7yqwUi6kuG13OLrszv9rbSL7
9XrVtijyEFjI+cpjeZ/IPCeWGQZM/zCa26UjBYcAuKWgQULo1iZBoFTbB+F7nvUtvPFGQtna3Mcf
5JOfR1iQzw22P9wdkwORf4SYdGtBeka0kyRuYlZUGnzCuTLFaIdlEkmnxfJZrbnQjcZPsZhfHNkW
6GtM+wtM3woWJ7fbfw0wdEccT1TiAL3l3BxuWrBEf5nf2Gu9I67h2ZvAkwkkLn4UR4Ehy14r8/ru
0EmB0PB4VZC/TEWeLNUDeT17q31q2t8LyQfQ7BzmdEk42RCkTKVp13f08fvJzEOaCXGvbMqZqYEM
sTmsvXnDJ7vIKJ9k5a7ULhbC0aN8CidA96hh28DtIDF7Wm4CzcxvVXZf7cnnxrJg34wzyae2L0T4
hGWh35Mo6QywXXWMnCeXEg2iAkDj2zcR5Mxd1W8oGX5TJYJWJ2VsUsOviDbjnSyZeBm4JCY5JO1T
buc1/WyNVA33DDCJmafZY1doRLpS04jX0OE0t6LrVr6OwqI1WuVo6pGEscG09YohaWCl8jsuc+aT
eUooBc8arcWenlUg/kxJImRD8aL9cyT38pnRvgVCLoBiP8NM1Fo36ixAIF/mxy8aAg2OF/df9aXc
4oCaq3jE5CwUJLrHsZq9fHfBuZcs+DR22UxBpqAXo4sHzEMuPp0BpdV5UBCKeFWymzguuqesoSfm
lFjQURgkhgwLBWg6H6ifqmmowOm3rRJQ9Xv/7EoK287+x4izNOiaAdZ14QANZmDL+wLXHhMkBTCX
XIe5pazCbi25nan1pX3rOaWDUduG7Mho1aWLYhXN/9Jcmcx0io0Kaqc+OF01xAO2fuhxRHMSazhQ
bLbtSggAjMmIR7NCzSOiHv2OKJhNe5IJd7i27aRX2dVko0jglQ3Jc/O2fGt1ho372EnTpmhzLx55
g2jgqeNU7exXdoPwnW3gVwaBRIOCOwtcn+WehHbwpYZyhHqblM02dxIGVtnVbT5T1BqdLtaUgnVK
CrgLCFx23NwWTjOAb/X8oxp26iuWSR/KEO8v9xG1Y4lhSD9RDfehHC4Zyhu1M4ubQd6IxT5W8ty9
XbkV5b9zXWnnvG9ftSIq89INniYgjSWWsRhtaqkJQMXCeRx60sjvMWT0lZvE0pkxMNTjIZpmk0KA
2IDjYdSfsAlq53+v96NH46DI1mdqYqtSdrtqCGOYSqTK3gSGj4tZPTOK+cPxJsP/4XXTeDy5pDx2
3xK/1PMHKwCPxfqzs3ir0Co3xvXfBRCML80tgUVtDFVhTUJeEDZOBIqQ/bfrzeynNmhhGoNVRPBV
Az7/B8nPHDdntn4PsCXIs0IgILMgdB/cdfcqM+rDGZzB4PT8jANIfRwnbKE0/9QjpBj5amUcN/S1
760klV7yhtjJjLpxAjFWqLr0TZW3o42zM617fN5D9d9HxWxh+i2phliOUJSVhk+VCXrBBH1BLNzA
JHfk2fFePeXU3l0qyxVykSyw0rMUQxxvlKlTIKE8IF6Pu6WKrMq1CpGiq5I+Ejp4tbzFpm8Cv9hb
jXCk/mXMhJpDl/w16px17jPYL105yg+6rv4NR2ly1WuxFmL5f36AFqkVOh4jilnKG4gIX43T9kc5
TKtMBKrQe4BXDRAfY2x/fXVjBYWgWp8CdNaIlsGjSxszkEmtlLFXl1Upl2YKrTQZPZe7ERhWJ9y7
dxHO7OJqmPVi4P1wGAWsNLwbnh/L2StpNxtu86vGTWjjOkBD6f7l5iBF6hQpz7IWdeiaF+UtTciD
lnZvp5Eg5VfK+IDR4gRdKdytkSTDHL/GMAt8hPkGjBOz5EjU4UtW8M+KY9KJxm4VdtnUukrWUc2v
KUtrGCp1jwFn6wOCCyyzUKPijpLBKA5+xDpF8ST12dUYfpwP71gA3mlgELBTPE8Oj0NJSGEvcyH6
zFMjtVXhi0YZYoedtFuj3JwnhBj10uOkCSHvOn/qHuaM0SaoMV/EkWq+9dyrCIlm+hHqzPxlf5mq
qrmI0VE9XQYSBZR8kuagrZZD/UZ2leAoMxxBM+rRKYMeEduaNjOsf2/ERlNChUoxWwdxRE/sTxil
LGvekLJeB16X8he7pZuf8LpsxbXiUxc7To3y4R1vLZbYAkh5lKgdSOskbiHZN89rkSUwpb+HScCV
92lOx1g8ATV7F5VJv2Qvn05s49Gb1V6Kz3Q3qmB9K7EJHoPRNmMDz6co8gce5BiEDm7xkg2IBX4k
y4Op4lIVnzOjqtdX6hdUfUT2H7RfI63sI2BFsj0+ywuRkM5Uc8Gy39n/4tfDHeAcwmi3ytx0lm2W
0yEJ8kBg+TK5oVgDf+9f8NpTdlAoC2XmkhNEUCB2pUMCrFVfqOu0URFmKQNjpwMDvOWmxR8Xm1bP
9B4BrGAXgi0SORXQyvHHlX4WQHkON2do+gsDaoMDY48Dmytz92n1+R/OKMkN+LZhJNsY7c3LYDfW
6Kj1UHMjSpKSE6zdcllGm8fiEcb1dFzcpokpk6iyjV+PuAxiNduN3i3R6XbClN95P+FULoH1H+t9
wbqzmSE2p/NOaDDzqWgRanTbNhck6mCjoaH+LSMiVKIy61gKAfkXBIpidRkNKIout1UtO6kuWBHW
BhZuCvUx2K//usT76Q2PNFe7aPEmSdT+tNiOEiNTt/Dz34LuMHLA5HIK8U/LR/bKPA9i75haKtel
b4c1LHLdv1vZZNG+QdfbrP+OhkLPxSOXDaXKNN6xkw0dL3+p3qKRJhUcPH2JwxoNeheuJkTRqUCX
Fj9beWQnHr/l9pNYZTObd57qizl31JKWMRp0/M7ohumNs63u6I5tahl4gPXRaYbjLyXqEpMN35mE
mWEeEHFydHRAzT3SgX0ycgoDk2mom5CITylluuBv+TOzaDUxIE1KDMpkkpuSm7hF/KRm0ek9NGsV
OY6c/Nu4gX+ptNcP/A2jFthCUl51BqCorm0pBKcwqke5NC3KIdp8rULViLPSFicSTTQWDvmXg5so
23LOop1UgkwUy9z1HtHi4FDHD1uQjNoV8cGe3mYEbn6d3LFp2uYu5nUy0SyoFHhiPHaTTrf0T4Hb
UlVyD64Mf2mxg1rGUgxMI7DK3pnb+Lw1HPbuoNH2zNP6RGHylGT+0yyMZolwaKDhyX0STzsi7n2E
DZwxxCmm11BHwt2f0HD1GIbcbQJOVQn9eV8fNPTm3nznKA8lxnDg1HmuUHtUDXmc45ku5TUTjhr9
VA72S8Gjk1rtLrMJNeo0BMMH8+D0se4pjlOje4daCEWfb1EPVBLFxpnVPXtDaKVDIEI6CK6xMK/D
4X0cfQ2hYPxPxfdgvbfj/SKLYA3GrhJyCS/pA+K+ZoX2vTQPFH4JaI1WzDDALHJ59Yz0MtSdfjWM
h1V9K6YYdvF2Spi2DeEtXY41YPhnq3Fg0EZ/dHejVcFvjdvFevEtoqmpa/QIXdsv6tklLKbsFhS5
9v3NA64hWD0zkar6D0wbdSiTMVnkOsQkrVh8WzHBFKvI2iP5RXV1OIo31NnFYWK1wIvJDR8OjWA/
zfV2k8cyVbGPrO3APHuvCHO6tB1XYjTjTfTSS8OU2P7E+jqvnaAGW/3lHWeer68Fh2H8uMe6Tfr7
lRpxBJVmwsrOcrpWbg4jrpVxJ8bSaN/7FRd32urdSzCjO/xLqRrVfpYbj9U9Lwwbpz2q3ePjoGxW
2dKqDlXQ+lZfVNKqO8y9O+kmfDhg+lK8w2GXO7/yUMMVfZ3g87amwW1lajcdWJOS6KT0mRZgv62O
xAfBRjcYbcxCOUy5q5D+ECFsEg4JUNTWOeHKDPuQBIwUhh2it/hLd1k+MZdk3F6rVqnKXq6OiVaP
VsE2KeuGRL/s9eSWeX0X9y6T6YxRwYrCTaMkaa2DcypXOw+ELZimMyPIdMOKoVshrgcPZ2nNeWuB
dkgiX1C+Z2oe9G5u2AZubvrcgLLH2A+gYZC4rQZFk7e6+awQakXR1DJkc+aZ3UoLnAWQurq6nd1N
b33EZO4CDHi/leA//vY7ku4jD7qdyOQQ8FWebJzQP8uHaAiytiPyFa5l3s8g/iy7W9B3//aKxa71
z0FFQh83JEOFxjimWTMzLqc5f0EvRE2GaYiHgN+g9DdgqbIYqEG48z5LZFTEFeCBRyg2ffy3Ym3z
1rZykvox4O5q3hOPfc7x6PCEahwS4M1lcAG36rUwbBF55mbhUJSVfl0xnXryCLXE05OPtXgY/TIw
CwVq5TQdEY2ZU+NrORVoX8GUx3PAe+7xGT8+1/DU2+yKX/sBM7rVY1CcY1KjMmWFZFrJUvAsHU5q
GwxVDrk4nw+AT9LkqwFezVSpjjYcNWP5pEzQyPe6FYv4ggV+1CWMgk6i2qvzHFGJ+f1Y2JHyrIhH
BlmvZxpOMRHbkYCET1nrGxNXcstL64EOrO45Trm6L2+WIPx2ZCWhcxOj7EYcdVrbiCm5Z5WMVM2D
1W2uWlldjZ+SwWKQtxN1dYjFFBq+YL/TJTkTkjU1VcGqjRQTl6nTCqpzqsMsW9EJBt+S6ZCl8mLM
z3C5xiLuyCswPI9wUzKExXT0n8DjZrMiWRWd9EiiTqE9knzUF5lznDKAc3MbYoa2+k7/xlI1Wta+
suh5U/qPW84BZ/9ZLzYH304noBqIlr7RByGrzxj7DB25qOMk6tH6OmyyK0MM0vEavvzl8M4wO7pv
EE511JcoUAJYY3CDfa9RbOOH96qdXk5mjjB8D1+1FoTBW4omWunwkkSHTLXV/mI4S6n3vUNOgSZB
riSBWp2r2KmhYw84ywzyD24KUL4s7tqb1ph1Hh/2esMNtEneIlXdVSOYIBHuz/Lo1SmFvAh+obPv
QpKnZmXMq47U2g88Pl1GitA1AWRgAxRN89ZZy5HfGWD9EVaDKdz+O48GpeLoicz9/bMGffQfHk1j
fuQ1kd9/SbWTVR+5qBu0kGHIzluEfKwkkUDyRRQdsm9OqTN9LSRZApn6UctTzZKt4pPKWKUxfBtL
P/xD3MQBgB0l/SE85By8G2dqUls11PbEYsaiHVFf4Q4efQ8mg3Qess6x7UMXqyFId4tb2Lw5QZE2
xUIEZg0FBEF5WEDbCf6N1NJR3TrSXAy9g6zehRhe5xK2WfS2zSAeq65GomgoYOAyhf0yUpkm5/CC
OSL/bhSDauN4wZ0hpc8zyCgBjvCyswrPe7/GnLzCT79M7VaHI4lhiEN2l+kaJiUpumi7MORK2ahk
G+GkfMe04KX4/nD90JM5QuJOfMY8olRylDGYHInd07qW3evaF9NMny3sQoMeEzAqNELhrwFq+nwA
398kQ7IIK2uXjTGWzwNOErqohGp/L4x9sRxJ3+XmLrb1HsLrUjnJt87Wcuqg1T9lDLbuKbaYrjKi
E0ssSNG4YWhCa0AFCaQmHTdoDsLrq0ldcNg7LvlOzozfo9QDL9dQjcJQFcFWkTnIkJ73IK2tbZmW
1W0e8GVuHKzYZocYlvt+KOPVpW2P3YH9jOuEoooZQAkUU2JSUniS36utAEG9yNI9AhbrpTgS7Uvm
Dr2EHcYGdLJBNkT3XPX9f+GZqBr1Jdpm76mO7CNkijuy6D0BQpACJTvJLzlGKzxdQ/tzGBXnKFAM
7gqRtwi1uDwH+bTFH58caGgtRwE+ibvjEXbCwB9XltD+ANET6YLbcoEg2i/3y/10jq+k0XGRvekQ
cs8r2VzOM46+nUd/0dfDpIGPffM+MzHoMbKq4nmB1+XF8ROka5AK/hNjLZDHR0s2XtYvm9rp1eTP
6AhFUQSbXFpX8haDtkLFb3CiKQ1AY2hX2pZewAo9q1YnfzwrmHTE9K2VEGhTIeWPTCCSSzn8KfIK
hH9sOWa2cmUs/ps39HTzN8tIiRFtwdzCsZNKQ4hbBTLgU/6HBHau3mxOZLuPiwKp1tvXT6FuTF9p
nUTFBYI9DT+fSE/cYpMobhR9uGz73jJiFhsobLbh5hjqIAMzjFmI8G4aYCv8r7PAoh/tf1PUc9ZQ
jEDv3l33Awpj62qyc2NLThMepd9rLusgF8Ky1Kxd4RUvw3L8KsHDxxXxy0m0dE6DNGfe/n48W8Lg
BhwvpIvSH0RbXbaZI0qdVmTvhmbJR3+OBRRFabFJq0tMRI0stG7PTVGjGyqR1A5DmScCaXW5Tv8Y
IG1CkiTC6yszwnajVoKRGjN79yJWElpIekOyM21Zu24LkGB48xxzS+G9teGeCWwzJ1QLw3Ov+jRo
1VUCEHC33GwCqplISSe+l8P5r+dim9boa/viu95GHoLFcmoKZeq7/8NnAQuLCbZ2hipiGumqjC75
/VaYGYD1cMukEUJg2oROurmmgQ58t9jWrqaCkIDMEz/Rvw30uWEwCCEuQcL8/ig0VygG4ZS08wIi
laQ/P65j9hsU94XVbEepObp5v18Hd3Ve8lpUcVJf+Xmbw5hfUVw445Z/oaq5lnWBrcQHRyfpUGNg
3ySDUlPpVcHxVyvRkWtqvQx0hx7IfteGokKZT4jUTPaRzI9kOoAKcZT35EpZM+bwnMoGupb0yFcM
RVGUT/uSbfdkpMRv2GDUyK6hp7VcHNdlChyTF9G83eHr6iEjTuymRzO/0Soegr+haGAV/T3b4FDN
FtF3hZ5Iaf8df/ubqpcx9cb5C4HyY6Jpto2GbKx+Zp2946dmpGBsgZ0N4GHh8PGztRqtEqitcUZE
Yp/OrDJQbg1lzR3s/zC+IyAc+aGTuoR9cvn+XAU+JQ9Y2Z1ofSpYPZyBhGWeT3LTO1T8FkHZKFj7
OLuCEaEsssltn2dJoO5Kf83cO/wchLmR73YMQSxZkcZnP0AAAZK+NioxD8whSHOQgLZtf9Yuhzv9
sIWzl1RHLv0IWgpakneDehoqnIyztHXuSI6HMuBLkRG0nhfQxG26PiLIcFELGDqb5+IJmOYxy6sU
yzMlRvVxN37MVPRZ8Rq2ottpW+ftKdd3WzVhBcOT5UsS+XvpwSqzZr5xl9sha4hGFEf6MQkWYet+
wricTJpeYhWr6irC1r2HysOvq6mmhmqTMAc6OqLj7fk774kmrziBwLwxjd6RPd4vnPWbHnckx4d/
Gl3pyYd6sNt7wcsL+ylfLAcFJAmh3Qo4kXFQWBoqJu4rO9qRYDKVt7y3I6KdDV9wB3dZ7oidJqRP
Vdex4fwD5ijUSrmdYLpyQHuySGv2PAY6qq4jE+g2uO7cAIOz1vliLYFDSj0zJQS2XU2NP1du4OHN
nLy9LH0IMVbb0Vxnt4Pv7uXYJTLUmnxPh0RYg3sQIbgX9WOCS5jmVHaJqHjE2GXuTeYagGG/kApr
y841FrD85ayw1xCe7fLllAUWpgpf8WpssQlFr1JEXyvo7y1jSAeR7AoYEIZUqG/8CoyVzXwa3vL5
NNLItXJQAkbjzJXBgB6WjSeRjnKneLr0uHAM9Xp7Q9pCQGEDHgz7MIDxkCt/M4xeVp+LTxYc33xB
ZonSvk/7m6cnJ3yTAJFXDBEkHiYYOTVkiExx5BHDE31qylYI8f5qz/UIOkmMraU+x44SKn1VO1W7
VjwOF6dgdbJX66de94bYo+M4r7UE5/5JHMibzP65jU/fs9YcB1b4bhh9pMx7jZQkYxgdKRqwQTaa
MsNLJQb5ebnLqbtnm8QQyllkgT7R/Cx/YL0HKrRErwxoWTnmIi7ZTlZGDK9AgBnte2C4FaQY5BJz
9IvHAM2DafR3RkkVe6dOF5g5fhFCLrFEAuuHy/rWhwfVcYbszBCQWRcq0JqPNQHRvXHyzL5qJQsC
uhu7Ve8RyXfIIMgR/NByo1lvb/ZvB51PodOIRMsA9prc0uhQMKgcm9tzgciONcGcVh4DrBqFV1kW
mNZMSAydGrsxbLCBCZ0q29PENKG8YMAlsOQdCOww0PnrBHxGD0PnOEYqhZvqjYgW7pzRVhVLTuM0
EXutyTVM04/D0kO1uZG6kuO9gfzRQCwnkvuN//USm10sjJN5sJNRWFvDqLUELXJn/GTOLeZt3Z0W
1KIxcWax0jXlmYXHV9RpCG/GNird0YKTjwsz9UIgnFLcYLedQYgp0ZmJdBuJVz6anNaELM9ZcSAm
8zhgoSDDQTby9nwOn8SOiurZs2+3xW5qMrLT5aWIhCyGKngZA2QpXAFERu2HxJfTqFUJ64Ifm8BX
rUWJQCOokD1goBqvYu4N15q7QU1QYYl931P6Bksov9k2sWwjUmJDJ06Q2QWZG9c6agSDmuMhG2/A
J3iYDMa7YnAH0cGcCXOyd2HFfrx+y9rJW0iLTCVIwQKOKjYdN5KWkbrarLzDKrpVBpKUg/oBhB+T
/lThzcly/xZW5J6q7BpdJelzxiHdWrUBs6djKZdru28YMDhzIfMlFU/NMrba3UbeoVvoHLP7VTKK
za7Q6RDsS5uLGUVZgjTLMb8kfNXuMZq9pSCA1NHCx5rx+LYS+96Mdw6tUrqy0S0alLVxEOD7h7Sm
fGj2EEo7E1HpWfEii20L4ezzpmtAzDUHUYOfYKvTr+dY3qoj0fDzma4+xMm9wPYf0936xcpQJ6z6
FNgxf/GScPGkfUu8u5lr77GrNEJT9SOtjwpG8nEW/pho1Mh3mTxz+lY8Z3O2aSMPShgW7/KtKn8q
5HbeT62pG2Bq3Ko8a/SLGtV1kcpbZmt5aOcHmf48OynsDVYvnMLo0KvGzKS51xbUlTk8LOFteU7P
wZEcmj+uH8rBpWZNYyLjzHm7eMqJXio4uH4rn62eGerGUOL+yb/KfY68OE+Bbe0HAmSXNlQkoIb8
DKznlQ5TSQifjBvHhe4BQiNjzR094kxW2zE+aeYaCmxmm21WmsHFd862fc1TyTDpj0IjdReRBIry
S0Rnws9eAxSVIGUP3M+WGsOPAF5pAUtiw/pdfI0FC+bTfoMBaaKhIkn2PqVnT/UE7+wjs+2UG7RI
3giuFizCVboUyupqu7dctKRb0JpsqMettU3eXioqaqjiLagBcxZS8eccwp64OaMKGqUz8iUIueEZ
fWVzlBPpbhwS6W0BLq80eermtd2ehkl4ZUN+NeA77noOOg9Rho2l+NObOuNHNOTmoAxP9L+0p8iK
cpdj7wsT2ba2jqG9LfhVl7zPS5oIA1ls7kX7sSRBV1cc8Ete/V+RjQVbayLNUqLRK0j7lYldA0hS
nNknDnzyTqIiIrrl+BVvk1G7GtNiaq8wJowLwUVwOa16Jrc8e83Dje/UAx1KWMnq5zATyNpJb1Ik
wTkbg3O/HTLmDqzBjZl7UMK0knv/3Vkg6zj2IX1PKrut+SKL9E6XSQDhBdtghI+u24LMQ7iMgTGs
ekzFU4X5D5nX7Lv9ZNZsGECtiio7k6CVlI9rTuBOt4zssawPuBJ+ny9THXFt+pOUmwb50NYjFDFq
9+TKn//QWlLHrWZR0cq5Iy3ArMY796eFlBsTnuwZV2M24W66KCaWGzQimNBmeCOi8mNJGHGzZo5p
Na9yn5ZsxFitnrJWDTnHrT6YXNws9dnIrI789ICl6WvENix4WKAAWQnhNRVsUNwZrWbzDSC1fmVZ
P3n4x5+GSAzvoRg2qVzSiGeAobZF61eQAyrI3Z8ZOV/m6hdHKb6XomPnaHus3hud5bJkS1vROBVH
WbZpXcx2ovSvcFYDaiGs0EpLsAF3X5XttQDy4509VxuNoAZ5HbmJaWv8errczTVfm8fRBbQt5sn3
N6TD0XvnGwkSDw78ahLwhepiM0/VzNolBhgYKPZef5TdSPqpnzY6e+Qlx0c5qWMWak3RZc6t1XXo
/5XVI1fyt1MB6P2lRlaiOhpRlTLOlNKAvknMVQRJVV/Wsz89tWzKh8HT57/R7eh/TWBoKkAkVnmo
t7Li5HN7soeVp1buBy55bn1ImiVAr3JEigjMjcfn9bxzbVpKga7ONMV5ym0v1B1bjSUDRdpzZ5XL
RUUAZaWi5+fgGgsergbL5Zjf8cBcc93xwe9I08FyMSEqj5NL6uOp9O57QPQsjbhXFU0byNjFswV8
X43ryPdXgWCVdZXRoK5rL6s7CSRF7IGWWXc0IR/9P+DGxliZNXOdxtZN/IncQWoBeRkm3U4SqSte
PIJKp6YYYcZiA+qI5aOdjeHaxJ9/BNbtZW+/iM6gQ4q71Cm4/3/wBj0Xm/Sur2OQquvwLrO0aVop
QUUmgiMXZDIKVZvxqsnjpW6k+stJJ+DZgf9Ps0tyah6U/jlMaU08jfrHZ4bY6vOLVwImTY+DF8mI
otXG0W2ByDg6HaH4rjfIjHYuPv0ofc6iXfcblOXWosyyqq8XuX+pksJ9Z5oSLHhF70wNBJF9o3eC
3XH1p74mwaQwj4Xet3nzIH5EJVM/g9jIi0sryXTp4c1VCeUrFqJ0ZED6FfOkwot394OB3MeqZwqm
3mbR0psG31fNvEiE/SKXil1iqpVngMlYawDeVePh9x4YAy23OEs3o7k03Oa/zzLL/6m2scuIS3m7
Lchpdd4aDU+68i9arfy64AtekoWmmlhu7GUIG8JB2yQhLBvoVjPhgxm6Iq4k0o7cSV6dpUFZ6bJZ
ztWZdQFECkipi+sW4zw7Web7hpCLw9QNAV91VHG5WJAWETTyVUrUUrQzFWDBTIg5koO1S00dGO/1
bueT4xVO6r+25S6/aPj+sfyWQghOZt3N20Pb1LGTbM/kJ4rFVkMkYfj1GO8T6UNyjAIUb1eFccHA
ECTUpMXsnFXbc8e79UhJ2jMAzMMLIOSrjG8A5fQQ+AkJvpljM35Ilzp/v9mYFrkV2Mt6MVBoYqd8
2BWAjwTMcgdEeGmimBBR8ccySyZsYPrGlEyLarGDMGiM280f2SndO9j35MmVU8B2b2dIzr9QqEWW
1Gp3GcBu9Frz1XGsr5VzXcNyUnEQJM5iAbUgf6QQjcAXu219seXG1pLvcYlZAzxCBbFQNn2dxEVf
jGCy830v3Yb1CdKxvEzAPRoI4FV+46+KUhA8L0oRhv1tEHI0y/AIIbnEndX58/iBv2iCp0nUruGY
KVt/gs8H4q5oeZzkZbtxy8xtaLdrgb+nnbQNa1pNDcg+8ijkZHHIyWEGYTrULb169JZGnxsA+RQv
oZ4Jy64Un2Eq6QLzAnDeT3Rx5aChSxqTaLAw587Q4vAo9soghrtwcnulXbFj3VSgDDMUI0PSxwEW
AD3wyKtzCV4PWqEVPWosCmSC9ua34UAlZTnoRE0IzVl4XMw7aZcd0ELbnEK0siCnjL968bGbSC7+
55rlkEzCPmkVlaZhhjFelTWN9QBzeMzolXMli2Loj1FgUSfF2dh8YbVpqiRGUxBwakTnEM2j7k3Y
7vX7k7pNJ37uWgfNdevcsBAKeLuL0zwA8t0B2cGDvVL0z2Bieoa6neKBIQOcSMa2wb0Ts1/dpVH0
I08rUdqjd7OCn9dN6XGT4SZz5ii3Y2sdqQAFX5Ack+kW6p8zAoVVMUXLGsQPP19Q1rCjnzO4BnpN
7e50eEr6xlRoAJqp3+SYxdyvcos+Rme63ZRHOfODdKmyEd3yumIAFYORoDoWs74ZBIotx3XktMeX
KBmQAxSikWz/STRF6Yj+F3l1hgvbI6XY6Iw67y86MW2OkzYBmz4hOY2tSa6wi5lSs72VBSsZcG6h
mpqGza0cbznhtlrPGDr1RUvz0IHuaUGmUOft5j9+0SoSVbmQhgSkUA1l0rPVq2SPwlGsK425uwsB
Em3ItgUOHnblwl0/Eq46T/332OFnT4FwdFu3y/3Hu8Ln2M35tqT5AU/Dh1MvA6Y3tK17lbVagVJx
zo1axfMOY+6t+quOqom1xDjBDtNi/byrUqmcOpAZjdwxiCrvImiIXOwxtC4MIzn3vhwFuF2AcUOW
uOFBietsMpWmYhy/WBylQHCEkiiA9rniH+6Nl/mz/rmSCVhx4mojikj8UfGNghrnEZMkuGjebyMG
SgcjMLBnGb9hFNFrwrmmrcC+COgSaKKgtB06mEtvWhwFb+jSvEPCB3L4G14hXALUfNELECfHn38f
YuE8zH1vQdeHScDa3Ovt07H78H/YCmkSkY2tCmeWxw0VDZmWBdSAvBD8G5v/Gu7DXo5re0Il6TGR
KkZvckEBFFouAfG23vLobDYh9k08Qa8+TtjUK3AkBQEazpJprkOCTGzzEwsMM2blT+UAYgkZi/Vg
Ugv0UrzgKXl4esUq7UA/Yot90yFD4I5bjUVchVSrsxnX/NDGcOSx2COgAHNg4S7wl5mZzQ6rDsOv
cx368FS0B3D4bjwA2mgEJJTEC8UKd1/q2OT9ouBe4icuqtkRoRmdgxGpM3LasmiAaV6A/mFLSell
0TYojdyRQs2TZ1fW5OOgKJ20C2bZhtOqZ59tz/3FB7okS5cF0AS1QiXmGnp/Z6hlEgexI3+EkliP
KAD0HmRIF8KHWAviX+lJCoo5co+SOnr6yud/fvi1HHy9JcgczHP3ceLPIA+PlhjsLmpqR3kqxWQF
bU/1cck08JVZWhT5hqYvmMYgE6ls5OaypF+lCfKc8TDwG2Rn0NGhtK5Rk4mzTC1CdtPBulslABAu
vuBUtdm8joGZX1c8HxHn4qeWR3xgSqLIMzI8uzWMadK4G4Jpj7uL5VEwzzn3OY9I8bJ78xZQ9Vv0
b1bcnX2WMIZnQ548kmAX5W3qlKgxsLc7Lq3bNNuZPNvZjUc1x2PHJiaPOnu2vyUwKXp4iTgfb64H
CFKrwMpo6sYf5hnQ1HmMucpJ8fzmciG0UsjH0hx+ej5NBT2seVls6aaVgRbAkzpGGO7Ok6w8MGLK
dqxfWOi2H7iIGELJt6+pUp/QbubR2tH+LiR5I1y6r4rNQzJz7jLIO956ZPC+MVW7eoKsxzXLiIwf
vkM9LyKIvTorpaKHRevgUcFikgUqzKbrxN/ocITvMEKxUJnSnYp3R0+MI6kZ2ODGbM7HlTTdUeTH
L8Wc5PJCNCZ1iGT7/BJjvEwYbOeb6FomoCXsOyQ8abKxjVlqSc5gJMlxtjdypk3LH/YglXsRKU9h
5c54iGWnS6bLl+c0GkgT6THDlEfPMUf8UAF9/tzkr3ZTpa0Zlyq2E/7Eoctw0XaOqHG22JT52DKM
5mTS1v5jd+xIj2vj70P0dDk+izuwYvF7XhuEwm5U62ama/ho6r3Vt2HmRzWMy+Nga5KcIBO1UQiS
fm7WDegiUHS5jGQkRNkKPJh2+WJ++lrEk6IyWj0BFex1hdHsgVtlqCgHh9bT5T42/tdMmZwaCRND
Tem8cXNY79f/iMczc6W+6zv+2QDhRlC/s9mDwXgacFEBhKni/yl1bKtQy1Ot7O7nLA8kjfAXdmY1
CO0VtjUmHhee4aqRmcFaBejMuRxtd8RTwYYjAtojD+/HKX55byIX5XiVJkV/uUOOdXWVLnTY59CF
fYtzIzrqp+ELwepz4BQqSFl0rfanvE1OYrDzKDLk4ckQajzfD2Z2DoQyPs1JPkDQ9DIdwmJxlsfK
5tm6qOVcwwDL/cY7jei3VKH2lpnvsweLKLs4tZgFa1ltUTOlGTXAFP88EnrXUokf3i4SUbJybUUW
/FB2MWtvVnLZx2T7FNTa7+lse1ZvDQepzbIWP8iuVOs6cbXDmd57F3anrefWsHPu20FC14ooGRV+
urSMVk9bKYjggaJ9veQ91jpR8VVKhi+ZHaqVs90HVj9dPEXg6xoGGpcGAGLC+Z0ZqZosc3nhvKzJ
QMs86YR4kAJGqo6aCGWA0erwsxJV5WHgE/iMG/aymTuw9GRybdqPVc+R4Z9FfldH3+xAj1QpDndY
ZvFuKsDLM0tzPMkjN6s220NtZ648xI34fDZ/4/J6gbfRhhKkPRlr0/vG4Ary/WdZA6Y4nCsGj2h9
RaWS+Tz71y8YarNc1U39TiLmy1dd7ICuOoEVXqJ/JVrwSQrwc6gnhsY2qq10ob1eENgzjFFswluy
MOwBic5bU/yaiJ+HfDWDmXLvtmi/00EAytlCap7GYUWawKh3SVu+JUTP8Gej4vQgObQ63tno2Ak7
Ri+fr6cd86vbbwcHjLiMx8CsOCRWJrnMFHKHTeDodr2GSTI3llcfMjS6KU45Hjp3bbZ74V95Quzv
20DCWzEk3HUZZyqcmh4gabDfYTMKzNlRI5+90h86WxV8UaSEKodqSbubICkWqlzZ/dGMThnhn8Kt
lP2n6sxw+4brer6UB+ga+8rxbEW711Nk1uhsO1WpTsf4rIAJmWCNw889s6mJHKBFOK2NpZhe9OFy
yyq01ckqLJfVUCQK7fBhEZV8QokzUQ2DumyFj74MRUk6szDIja9OqOYu10gmUwQHk0OsAJrox3Ev
iVyBi7XgudDBBYJ8VHIR5l06xJERFlBYwdxamxAJQ+VUZVMkvJ9qIg5bA/QuNf/NaxTdNGZaLxF4
vakjC3cqahlfyh2busvreYSrXCVbfs1JuMfYGA9IXEz/hblAt3uJQYIc5QS1NypbXLHCbrqzA53Y
MCWo01VB0J3vLO979QIEaNJQ427mevUFzDyvD0WpoOlvg4xxbLJGu33pw77UQDvb1c/N8jBAZFiY
xHE+RGBbCifGDEA/xOBXTONM2ZHq0DBBzPtWPLFtjfa/MY0whlD53QwSFk/sMa5u7BM/wJ95CXY6
wMrUjJhJulIJpGmgACxcZN6dldXsOgPEx6kdCB3T6OCFd0R9lCwMgHXABVbQyxJd0YKJuz/0vfR/
steSl6hsxNGDrjzlHAgKHXPlOa+M4AGzx0UCwl7TncY/tQEwnj/nG/cxgLwTSmHNZhRakRGRRksD
xDzGDnC45K7nGJwsnY8T95RF4ZtoHdlPMWtRSU9TE6D/hdtg3Ij5ZqsFI88SMlkGQO2wHkUUr/4P
i3yboh/N+AA+/Qw4Gz1M0QNIHv1HAtNwUNMH7fL+FRsDPF+8fuhj0mIzM1TWagax1TnvdHvA3scX
xqICbwBGVDtBAYsWb0y3wfNd65TYvOjvlcwQ1bGQ+f89+IrEfruK56Gme+Z5tOwX97AHNOYLr1z3
xNaqChq4Uap3PTml3NMVULVhm3QTX0qMC1xMNomWjVZKNzNONQYDU7L1fD3NI/HON7jLVDjhVk5U
sOlZB9XpEu37sqh3NV0jJ60iyoBcq9Z5HanzouoXRSCMUorBkSJcCPkftnAtNUA479wyBfCZHEK8
1ly3dXcpZ5Wa8JvFDzsdDRlpMwRCciFHg3JuRNVRCg5WAGj+qNHEqXP4ykKwnjp/MGmmRyaVfsWL
mBeH99JPWDz9Lzwp20W8oeLcYpwF6umDRR1dlumQT2H0CQYWMw4zT3z9i0QY+CkKiffyr8mHbwsP
FvQyjI1W3nJaqhUZjV5q1sR7RribpxPPKLFTygYtkdRS0UFlmh1XlZ9tGoauhMPOkMCMS5kh+jvu
PvUPeNaGdaCUBAuv5yKJtezrI+X9WUcZq7RH0xJoudZcN5fY57KmsKhhH5eJiBCJ3JQbSsNMPL+O
yKimK3ixGRxaL5X9R4LUVvFt4/OZgVKfgNOc9s/yWaZELppcJjWryZRDVeMRzjH+or+YVYa6QZam
nJ0ryxxbu8sIHGrZEUakW/j3ffjU5ghaA+PhA/iUvgCXJKRHzLfMZ91OOMjKRfOjD0i7fK+QTYb9
kevkDuC4zF8833Ta5I44KxjpJG37PESDhqxeCeZ3XvBVJlpk1EFCjExj/dxjlcUy8+8KATnCRPCE
DxyfmWfVVrsiDUUfQ2Yckldxdl4WOVVU80Gib+06w8/x1QUntFXuy1obEiPaE7vJkxtJhRIk5GRd
i7Q7zCssQ2QxTGAgTZ5mNrDb/+EAEm9bvwZTsyWzoID4p15RbrxefTzgHhdPRDIb87xi4WMBWb2M
BI2Cz2bl7SR4Kn5wgdIj0kyEpBFYFrFMCSyy/8y0Ilj85Fz2htN0xSmjslGtzw6v7/0gmCO59Yaq
yie3NmuPKAKj3pWgLKZPB9HGE8MjI814CmTvB/d3XA1TEfXcBcj2e6wyi6yh4gUa/ReHgMn5kFCe
7ALwy1wB4pWOw7+cmOahf0Yx2pOtqWbiqDW+xyDTkoFtPYWt2ThS8YFlniEDUMA174v0jo9PodJa
bOIMht9apZOyJEu81k6GVEDffxDPIa5aQqNDVCOPWclIPienLMuTLssWJAf3yGtVpsP/ggX4Z3Ti
1Cvd8y2aBOFgVgT33rcKbL5lGb2Zrkp1mj9ynx0udOoMENTsQd8kuLVHSWZ+P+jiz8UNNE67ws70
vZBng7t3uDEbXgRNSidqGORqw66cYj0fRsRHIlZOQV6X/Fj1SpMz5KnNwKkYGPpqbhWL3aADQkkD
Mt5giXiwBVu46bzJ9GbHC/JKUVJL5KmVDG0ZsjBDOC99lYn5tfnJUmWHkXvTLMsbvGaqZnN0ojE/
+X/kdyIsIgdTsmUaWDXD6HpyKrQWw+6b0Fvh2UyaR+BFuI3+CuAP8KeFJa9jFeQ5SC0l3mlVAXj0
xZ+q4Fk1mTgAN+sy6KoKZPThXMVzMesHSg3CD17FWxdMYNaLXNOw52Hfp4/aEEoQ1s7Ug0y3+7B6
8yGZwgZpGRBO9laQVvHT7tLschupgx4ljg2v/BSkA/PPkBoOGCrwvmpncEYLf9akAGANTf5qUOBD
AwLDsl5SiHEKffDaBY5HEv3YdyqO1Kwl9l95qKVo8vGmccU2M8zzAAUw2QJs1Fa2LDGtWunQnf56
Qf2iM+T3HL8gQvvgmDsLj3woDwBcQZwrChBE0hpc92FAXbzj4k6OsSdKdDy1kX5JBt2BtBN+etaB
iQHp1TucZaNBLm/NiJ/DbiePgolDWDP0XOMV7xeYLS5/u9qt55u2XfGSZgk9cWLnEMApQFGSa5A/
o1uSqdsgvIAh26lonydjQ/2Y1xC5qM9u6wjND5GbaqgpUpepT9JOlJh3u8ivCl8xiq88OmOU0/lA
UXdrOoXDs5cfZWn060vLUtY0dmBYC28hAJZibniPRdk8DQnP2SAJhs+fg+xhkEbx27FShXEDSMdP
whAKFmKa4FU8n6TuCQxU3gimTBOhdGQ/B4mOtBt6K1yylyPo/h6tmPw3PKG8JmAzSIhmIMcE4/E3
qWAvgJt1Z/w0SNTWnqAKHaXtuGOTAMOOO6rGnYJCHwcRzce/zTdO4wd5uEjq5TAAi2WwmdfMcHnb
daZwFxIv0w0VGdYiwLqN8JyPaaSK89PJBJFvuWaKPwcibbQhYKBPgbf0tuMYcqOT2eeoHwgKxolM
AMUdQGoHA4nWldLZH+FPVa5tToYUUcyCbJbQsyCCAtGwXzx0ihB5Hv1+qeIN2Qq5/Jj+i7LcuZRt
/uJv+P71uC3fhfuvOApYzOfWSxPSoAc+3B8uApcsMlcdNpOoGJ5NBNphJQ44UjmDlQ+xXsE8iIM7
S67K/9wEPd0x39RiXlcB1m0zyIifSirPvveNhN5oYUzPFkAl6Q++39XGfJXG8PlM7LrTUH1zZkVd
FLhsmyswMItxKdGzXw87bRt/yJOQNrWjGCqPV151JBe+phZ3YHcM6Id1frtp3HdzlSQEgN+ksOLz
ZSHvXn6O2MHZ9RJkxoEjFuNF9KKcz17XxUfRfUxOP3saVIRNgIdfSDhKB8Yp5faJbyWv+XfyLYEW
ZlnmhfmPdWnMNkWMMX3JGO+GjYCYydud6rwn/vnpQXI6/Q2c7k9bQrauCLKuPDuSDZwXpFenxpNa
RmEZaKeWMg8NtF/vo9ZpIl9hQd8KMdtkY2KvCm+tJiQSWx2F34Ih+JbU+ZEbsCX1fb9toiHH7A1j
DWLYQTbIwCn4qVMSeuxVa57mU6DRqMsbjUSFqOP+54dlR3W/VDP7R8Q05EdoBmbEEWqxZgYBhp6K
yG7pvK0/FIM8a1b/HmYMCtME18o0gXjTXxsJUR1iKpj2oLuwqtEOl/9TP00wJ0kBIm8phvNtinTm
G6RdN+PUPvOQVcjhlnKRU3eZL+Qd+U1QXmJqNAvTFjw72jEhwS89nvY9aqtFIuHOdPxqll6WEKlN
ekzJj8WnGLQmajvuwmOl6mRRcK5ZDkIBtBFUPmr3uFZmVDy8pr2WJGoQHW5yv+kT9WQVKWbVjXzQ
iMlWVamcNAObLMNBH0hueOl9vitOw8fz9lGQzP6YQTiHeRUSdoa7N4ztwvpmwwHmQu6PpEQRBli0
R3ApODdWXObjI6eiP6LiqIRP7nI6yAhM6XFQE6ARWsxfzti9d3Xq5jyh3Q2IUeWAsAYyngYZtt5s
zFIZo2yvOwQPHpHzLVd9B9vZfsDqa7bdol8VZZCICtn4+l6GE1Im1/e8wXc7LPirBrvmX2pSL71j
9wrV0HoZ5TrOyTu4YtijAFF/N7OekqPdPjdqvbCMTmlpkNOyqJ/lKTipDCkq0Xud5a/3nSn/MnT7
Zb3Neh5keSVsgQe84b+sSMEpuJgIessHoRq8FyoHo7bzHEBchW65G7sqlBvq+0C6gtOqCKb7hKsI
eJ8/2/lYSrjFy1Bg2N9X1lixkVy1385SMD+vf/RpvNBqH7w8ksdI6TgimOwkv0fsxEqt5665p36t
JUKpRrd3S2JA11U9DFz+V6VNGj0TaN2fPbmj/ukHVPoI2GT+mdO0NjfN+4OH2C9p6v5qJccMHiZh
39Ao6+0evxtV5++QEf5TFQh4ZJIRfC5sKwH0c7RELTgsm/KXDns9CF2TfhaoTCFFy0YBe6JZBAfs
HvBylMEujdUgX/yaJfiGxxc562HPeRwx/oajV2Ef/6a4wJJUIlkyPqbXRGF+BUPGL+2V5VSGRJbz
AIAl+Lr9NPDDRAVy1MYrjE76Ox0fApJ5kC7qVVaJPdwqgKeN1w0QxBCj4n/b2VwXEP55eBEb6OgQ
+g45S/3vEFm6vlAROKK6D4V/RVuNXSHvXNH8EQHSeuMWgrDS0zKUSkqNTUnM+urWCDeyJAoBqbp7
n32RehDSE4LS9uWpU1BMNokBv46N5+wi0UyLiUBj0CQ/zQBvczJLueC+3XWq1I2ZH9irdGxNX8r/
yZ3wrwerYdNXMfZPSx3vqmKbBLcZwRQwQZcnGxrWgUAXvfDoKpWJCRUOrOSk2d1FMf0yrEo1goUQ
YmmSg2UzjJWH7nqsmGRZjp0aBkqwaQLCe8WK3XVmbaDwsqZ6aFEQZrIO9KFmO2YYJLVViGoApNtj
4hlPCzUy89k9MAaeiJpWt4pkw39qVmimlLC9QVztm/MIO46EUI5ssH0HIu5quqlz+RggYfCUr8cW
ORbv/zufO5LD7hilHzbufO4tJ18F9bIdOPLBgBIhIUS8ejkgp+Tn6PcsxbwUbPJcA5Nu1XdkpTyv
Hwo0pdLEfIKA3ZOr8gv57q0YGu4UDkfAphBmXi1fOTMn6ghfYbxUaLHcNlWtxDxFPT+EyevG31h+
e4ixdGKIyS5BbECuuRdqs3N82Wgwix+gSBZu0qjb+GOeHMj4nSs3v7981ItkU2VMZNYnyRkbnaPY
+qmurFTifa/1snD/WbnxP32onkIbRfEGHNv3xdhUPhokDWX4P4mgiixTn996OIDfg0UzkrfriFeL
gDfoXrHgAgEHgvcrqWO2UqxZKsgmOROEEMsEf0WMfnkpymOtrxJ+QafjBx6fvHnjpY0m7yGar2XK
H9fp1T8jg/69o+aJEO/La0cc54EiiJJDMw4cQRaz7BfS/dYbN3gNToxG9z26TCuzS8rsTt18tx8F
8zQtJIdUIz68wXlCy0gUhi1tPFwgBkzVaEOrnTH+xP6/TBC4p9sWOWgSGUMH5A/YOnlXYkM1A2/T
FV70RXluz9qATj4bJpJdC1DLjPhc2B5lj5zxaetUj0Y4W4nIJy3VIOjV31fhMGDzH0G1cKeQsiSm
hV7WpEv8VDPY5f3dgcvA8m0TH3y7jJRB/nVYsG2UcSfBznuVqefPC2z/nXFRezlXhnHFaUbV0MPx
5EFx/xz6RxryFZkjGVmjUmH7XIHWbJBw3b+AjRQmBrCYhM6GCM11LMHBqugGUIS59NnyIKn2ek6g
dgeTPDSXt8AlVEpePKV5PVsKNR8whYwuKSxYqJf7e52JbjVE2JQKffbRGMZrrqKgkuhZ390pO62Y
EMFyOb8EfdTeqpwO/2eiyAJX+t42aID4UtTIQIh36nUP2oJhDRv6soivQDvIQOa02MlqjsH46/kt
Q2Aq0KbGL7uZpZ3JNKQvtnGUoDbhSgWmBRrBnBoNP6yGZU+MmqM5nJAYCJzAmwSEP/uBZm5OHroI
vyWxxaBLsCDoFgjcoV2o4kSq/zlhtafKkFP5khkAi9gsIdF65NRPfc8ZPbxmX2iEeGSChLUKS8+E
DhBrz31nfBptjVAfU4HJcikLPG6f2j4tDUBqBQkpFNJz0ZuOns9mFSTCy0IWBwOSsq4Wd3XCEY8W
Q9ftFnvhLEwLe3lmF7luqYQMcLUSX2XeFZLluiXmIK49VkLSADNUgR5eiP8vlh9/Rg/2Fn0+ESjI
HyLGA2MNqfrSeAekbsdc523/5UlJM/eMthFxj6VanWX4QvFwAE1ovoZbiTpKzOIMsvGokANg+mxv
6jqKU5MzkXmU/RP6zAEGX0HNSbNdsxmL2vEQNvqOqdLr9/FeqpSJugEGN+Q4JFKqf03x2esbUV1p
/QzPv/4hNU9hwEs00id/MWDEnJ/u+gJr+0/1oH70h+IuVCayYQoC80xlaMnc/9pmZJnpUoUIfRg5
rIJW5BXuzBbM7sJHS9DdQJZdJNaPkXn2iK1dKC7lSnW3CDR9B/W9vXLwBoQL7o7q8yqx7hGc2eSm
0GHRHxtK/ADBGZ8B6aEEDuBAkqY3ZuWg1f2tt//pbvNG2aX4BR3N7zhx8U4KCwVjyUGH/nPfp8Hh
pXTjebG36tTk8LE0yb0OBXfCv7hF2xnYfz7ooh+Xeq51J1/FjpARm+oGC5gXydX+LG+lRhNvU7Qx
qKexbIJFMUKJeJesHVxBVCuUyvPUfynGfVXY57m0UEllGV+N3YhY3JdhZ1/pWMOwcadpcsvUDciX
4IXG85FXBbTxT9HJIRAk1wgpYQ+jxCEQIBXVv8v6vdWvg+cLPDHyCaNzYeLo3Sw1M3kB41XFKdQ1
Lcjjd7HETy0Qnd6y5A6rKt8hwlJXu5REFNW96wsgdeuoELdu86rq7a1czDmnQ9rDj9OFl2lgLZ+8
D+arKj/MPyFwdZPVANcTJ//QARymX+pqISt0c5dFcOiESh0t3PEmVgfACN8YHC/+ZswGNHqGKO7c
GwGLqvbpAI7RXpQOZ1Lsu4NblNBbmiKePH/Jqx7kcHnkrIZ2DgkKXR1YFaAm4wwanmOUqH7yA3VM
cp4Fvnb+rG2pmUSsvl+0VELMDMetJriWYHTUbrBVcgGgBnFvP4Eo4FRVy5XQwgnQFUKCH/j3E7eX
e31CV0LVivcL1OsI+k3uNAw9aJibVIhDcRvrKXobVNJUtDERCdMtKPty7inbLZ45yR7Nw/hTbESE
j/1i+d0DAbZgmNwFBtCMC7klwG4i7eiCU7d2XVzpByc2pMwkZvw6I1z2H3nzkJLCZQ7jLfD8kxks
b9HeJQ2qWg1MWHU+u2dm5uzB6VOCiHdR3aTHDOodjyiKQmMtwdobQ6YbJ8VMz/8GZxYIMOUtBsyt
+Rp9dMjQ9Uzbk+IrAJ0E3HQNNQMCSWEYuG4Fr5avd9L1WGO8pEcgQoWl0gUg4LpOV1m1snNHVkOY
y/Un2y2AVEsJ9y4uTNqlQbzoAOElBxNHDV7fjU517gfEO6RrA6qHLoSSW++k4X/Eb1OQ7VGHCHZz
chP6YtVGMtcWeuQZ42UYAOs3Vy/h9LXT2NPU/dVRJz8ZciK13SDbVZ/fSM08Snhela7Hj/5K3Jjm
YmtS5YHfUUq9XdXFw24cCeRGDl/338c7bkO6/wLew1qTpO3Jpq7sEgt8vNyZfXGET5QghnG4+8WE
QYvsfajb2lfCn9ghWFndAF1bfCs6e5zYb+ekBdpaWhkYlGDCAcXOdKGNuJJDiTY+WGrz9SC/y+Hu
UbRyCQhPLwkSfE+A1jPwvOFQktD02MJpDR7USN6pEwYlOMcRv8+TsfCtCGjlQcR/GtGPZQxNcPEg
DCf2ARvnBETAX1UDTl66OtxHZ15Irr7e5mAjynh8zqtOckuJxEfgezR2/pqo/cSyoQlfy/ZFs2AK
S8AEE+LLDe9Vc+meismtWbkVyYDFK7H/0m64sWD/39vGqvRtz+Y4PHWOK6OhatMGBDwUTW7f0SXC
8yrTYnW6y2+xtDhMFeaNoKEKIXBH5vNb53mIJZCUDa6MV6OUJ2hmCByx4S/nNl7+qKxMnti25fzH
nvKwKQf8PJcpqEopLNkt7bfhVKAp3YQmP5cyft84dQJYC+jsXLaW7EtVyYES9D6N4VJPt9Z4LoBt
WMWaNUmY+/K369JcjS/N3rA1x3DrlQIwMPrL3jGhiv9YLuidG97//nzlfthdP/J3mZbH9pCi8kvA
WwpufBwAQPLwQsBIsykQ9KgBbR6VAsA0FI6v1BysIJKRahC/0H5MjBzhrbZ1Ty8VH9GWRj+M6BAF
YRHimjQiI374tB6NF4UfIEF/zZ5gyTCGH2hYtNHhkOGk/rRVsI9J7rEfPGIZsxLk18iVcL375HA7
P8MqItPwFrgaO0j0cepnzUL3Ie+YknKChvrKuoKZwTF2GE9mvxXHeShtF/QXPRpC1a6bXJ9EXucd
uEy5SVnR7m7A826lZSpmDnWQAKHUBby9oTRfPJw7HyOQVlkZmT8oi3BKrP273lz91wumYdZ7H23Q
rMU/+nQYyQt1sZOFSw46ZGxvZkez20b7AVCJgJ3i6dboDJ2SHsN4kN3dQsqi7d1+y9XpSvkkw+El
amPsZVgy2Og/kNnW3qIAwXuEttYWYnm1qnc6tbun/bbzGs763yQkF6M5e656uiYH1fLKupNAAATF
LvRt3ogzY8EwxI1wQWXgM6cQkWhXvME8vW8plUljiOgsc+3V/vucZvLFbGP/KYPPO0PWidf8rmFd
vc2yfC4S+I179GKsoYQewwQCVQSnpC+a5NuL/X/fnt0G0IL4/09SE0SrIAbZrtparj1gQZljSv5K
19mPiUG+dksTtGbJcPJzUDY/oCwX4QacTIFRqLjEKxKqMkrO0NrIZxBNVmj51j16RbbLRgB4qBFo
6UdOEDi1LKvKhXB5Lv1igEaxk44oll3JnAWZQvzH+rAJufw6p1l1haZsJiw4IsMGbFo1ofOvYvsC
zqpKv0abLSrmu5dN7hRow8F5YSTU5u2kd07MqsaGEWMj9P8W88lmwmtd2OH+8vPUEUydr4tRe9Fp
sdXxqaxr3wrezT+c53i9WS21VJ13YKwtB5H/6mwTphdxyAZZSDUA9iiRE0CPSnIdBs7aFmxPt4sX
mDchfe/qvRMmJf8Psvl7s7lROgvm21bA896iKBmvHdNIIILPcVGJoecibZO/nIUP07sSqhQZlfxV
/nc7Z8kGJWM3FVFqcuSKyTjPX9PHtUBSnOO90ryN4GcOfwB1xvt1Jinof1/7k+BI5aF3dGMM+I9v
FgZErH4q05AxbJ4PGa4GNI3dKfeq2kTx+mDMxyIQimQEpLcaL7bae96rTQEzN+/oYGXSRX03VP+z
epPAqb3aAnJicepCRBW/ngADA4u+egoFgYnM8qfgGF/ZTJmHFnQDzVhrLqbXpd6ziPYJcgpfxEKK
8yIh/7cItCoIiYy6yJHHXbFMTMU/7G3t6qT9lZh9g/fyat9tH86PqvPr/uvbVHYOv2deq3ytKpGi
Spg9V8zjv1q0F6hj3kmNYWyR65hFZtaG5h/Oy/om+8O6jHPt3v44UTzWHWPAcrh7m0LajmmHblJ8
mK82g59BJALimhSYQQhFdx/BK7yz8UlflbEGv4LuroBF+WFBwy7DIKRsjz6zHX+KigJezFw4n8HP
NXwk2EcDG/zAhOLqtpS9GA8dup7izWLsAnNln45jU0ABVszOW3bOZcre8QY4r8OnNrOOd6Dc8PLK
MgGWOxAPPi0Y8+zEG0O8rom1uci8amx5GW7yhinfzfbiyGB2vURPEqf7RWU/VcoFbUeQBM3AtUoh
OHv62chD3CO6g1VUfHTOhSoOdxlDiK8amwImOp0+4aJ6WCE9UaLw5b9QKD7wbJmNp/Qbpay7YPZw
BrjGNFOciTnbmzHQRPiFCw4Vsg1QGSfHi7a4bhucHIW4bFS0SvCru24bMpruw/yOfEsU4+gPh5ev
NZPCWkZqQDetMkkMrdFyHABjBFwHkiyrtiYieZ428ABufT6rs6yFgPzTF+fU1gZGzXLwU6vXD0cr
FN0x6JAXrIloj5k1PxnYadbOmNZlQroGQ0+nK5ssCOAQ2SCT7EkLg76EtFblPEfPWJSpaY6app2C
UG7Xm84y8b3rEyLn7yBMkZ126+/fwQGAeUH3yPKIFb6aZRrjM9OSVrRYy3kaXUkJ7oJmZAg0RYft
gfp46hzMVm/Tia2RbFlvEUj8zGuu2dn+UrL7xERUMbJuacxCDDaymJSadPcrDl08kXz6xE8leijy
LrXWLtRpMSqbm/csHpBiQEuMjrCdVWJVEH6atK/Sp7rsrjKVaoUR1maX+mMv26iTz+Ll0/yBGhj6
TlKioIlmRTWS0bV1VlLeE9L+asecikqtIkyrMiKuKJzqbfZTJIRczftmF7cci0fj7AJHBFQIY371
NwrMcjkPyH57teVnEDPubcPU0+5/Z28QrNk4Y9SUtnbc7sodjn2CrGgLyZPHxBR9kya+SyX6m/xa
RHn0WB/AEhPU7LbHiLqbugzvl1zepumx0lKGN6Y4zcJKrn7iizHog5yKt1JmRIcvs4EjZIkklS13
jkBApVbZUjjx74MhJfqoCfVla1Jul3u6v8f0rPBierGf6WCyKyy4QIh3fgl86HPd9xzZk2gATAz8
CRZQmiFYm0TZZHZTV/hRiZ4pRHyN74L8tD6e96ErKkjI47LFZui2SzqNtZqnIxz0Gy0NtaHG7vq3
OeekM5rd6HmFA1uSCWz9Y8auBSdQB13OJIhlp0qhmbwQMrQqfuTgqz58bc4TeErQH7OFxNQtoZ6D
kz0D+dxYBFlLXgxTArnEy8rxE7Buii/2lkWbXBQV8dLSs1xAX8QjBrv9O0hRviFS90KApSni2SHu
y58XCvkC123kjgN6hMPFamQ6SXjVD4l0z0BWKl3MzFhyQCB0SRJVQBEFrVvzZS0PdyFZjVsRablr
K0MPTQzxdUy7MXV6sjPu6JGDLvVzDGCEGZL0KrtpRqA2KHAIpJ8z1emopVZ39T4PuazfX9LdYC/E
d/vsilutMnGgRpM7iSntFEkrmMXa3Tnbgdw5wPCe0QFfGzgqn38WG47CT5XX11ZoN9zRSevmRLTl
ZJgmePuUb99xj4FTuTyk5XhiW12+NQ+zFN+/CVNVH0F37lPzjfphrcOA9U6QHZJQ4QabVEmBA8cd
NDM7bJb5S3CQzWAlHbJ1HkIPt6ZUdV8NG9nMnsGqMwkPp3wiwFyM7aka7AiZ4N1/6QsolhEJi7xA
PP05Yx+SM1EPd9QjJ5z56mitDHlCWWDyLpF85lu0zmWk73iQeR5lOX0YVqifEt0WCwkXje5ENuH3
S22uUu0gfaATP+z8aao8VvopDI03tIQiAaRnQHncJEacgMyhC/cVSmBKp5mjN2znYdXQeayxmZNc
FukFha9NWRck7J+RM8w6x1F5TzZzcxP+mR97aapHHDveDo2Yl8mv/lUDnLYH421/OYdrmgkFwc0J
s29krii9mZEKksiyTpU346SQSB+g6EWx6Kezv8IdygNJO07E7qYwMzX2M0FTJjEYB2mt8JPSyne8
Qipn9oXMd+IeooyHPgN/twIZPo6gWS8HsRtQwcMtDH+V8Z+BN875jcaFCHJRPBnhXotbi6RyQA63
uafIOQl1j01xnGG7B8txlz0LnuPIU9S9iEeLdxQUL7+YcRY4lkWS+pKLnAPX5emGVj0CiU+h2B85
rsJFBWcynPY5bCrobqcvjUi8Rng5DoNuYzjG+g2vX7SPqEdkqVAFN9fRQlIQBOi/hnhIZra7LWBB
td+qQVHmOD0UU1I4trFfigNEi5rgZTw3YkJxcpGOlVlGYx/nnFnxpVarVEebF7qzTMYkUROTp9zo
OP2KkJWu5V8ypMZGxr3wjM4dKidejxcb+OHOEtkBe9/y63CTLGTSFlj7o+HoCJ0XhTbz0LrQ7XL1
tKRFD1mIqH3g2dGc5Fm0AAPClMeMWrMzNyJK3wUnWB5oxnjXngfyzfXjUv39JDWIRF9W73m1BNW2
se4AwQOaDQTfOO4l8yGWdESTgsjgP9AB07X89j/bp4CJoHi0Nq9wHN4WhX2Hek1Dx0kEsdSzO+g9
wHRhcPwo8Qx3GJBTvtiUU/8t8Ln0h9b/qkDrIP7k3jqZyJ3ads9LHi96mlU9EBMZ+laxQy7pnrun
OWz7ky350oetNfX9d3Al3v+/H+rGn8rM+yZLCyEIdaqS+R8c/Y0xsapYbemnw7KR/TE9jbqwqYt/
askEIxCIC7rVANTPGffXH/lezNqmlO6VOLhD1owgROHGUnyDFsOzaWKkaK1xRG0K6VrWYo3gqNeP
vSjeggLZbvTxRkJdy4ahRA3le9WDilFcsxtBhGLQSLcSZRWyFgbv0a5KG69OO9kptFURDSkNhK6y
i3dBrxMg779reSQKaHW0+Zi9bsXsxuKA9PMXRz43DwrL6Mq+8VZATUdERFgLRu8AwSviIL1+TDyZ
9v45oaZKsGkFFalzVUNkk57co931l4bZ/WokV/+YB6PhuDjNE87yY1AR/yUN5LqmA9da+A6TH/bu
RqaYiV6Ja/ahInLCWfOTDYoCiwtMQ82o9y4xHHkuCpwQ5st4RJyW+OzyCuZXLF1OCwcluVDU7LKP
E7gcKfSlI71EOwS5pt1TVY+EIlymf62mbn2gLtTBVVyE3rxYKEdUPQ1XW5D/40lvjZw7bjMgrNLc
08lvTGtKUek1xlEAzwziTA9QN3Lhc5SlJTMq6m2o3UdeucFddguypKc7I9MobwqZIxKPxwC9Xuvs
X7wJulYYxp+jqQa/2WdEu1jmuL0q3cCwIq4PEuQUky3LjZYuFznCNnQnjy4NMQcTysOZAvt7oiWs
5qgw5apavPLq3XGerfx2XDKZvoZ0B1/K5s0I90WHbeOfEA1OmWAYGf127aSYkqG8rXKdks/z3SVM
xxACUjv/ww4VeBZxIe9iTz+S/tgHTWczfk+QHkBznlfA5eraAUZIURhPSnR3V5IKOMm4tvlEaPYK
ImjCGLj+naxE28iicmUPDaIYckCUP5inbhGuj3P5mij46R4vOEgzUws2Dl7X1EnnghQ4Gx2Mg6FF
LBdvxRNyfxSEW3df79P9dxwC77/AJ3E6gps8AyNG1xTq+OJfxidOESPLOjQxPL+UBpzFnQsgMF3G
2lCd9bCuiwvUV/Ovpn23xYzU/a1F4Zaf5N+Yy6aVs0YAXYNiX3xuS1/rROfOP3oX101iwb5FxOhX
Zic+eL1jjvnMjiLC79fmOcOPLufNfBV+WY8caqtcafA8fHh7xicQQ8QcyOfMLVoK256UhwnbVFwo
MJeNOLfRVheh9hstPxW5vNYKkqeg8714HfttGiOw2AicBdGUeoYDr7C48KxISGcL39iU0FyeAa1k
Zhw5mUkoVYGhBD6yxYED769VabAVo+oqn+ni57KVnkSejJXIvc9uwNHwvSdNep192nmu2sQOUMsp
dAL1xTI7HricH/3gIJeqdBUYIVWYOMMffP9E94s1n4wOdlWGO0yCsY2BfHKBhaouctZMvSCbPEuW
ePAvJzOkGa15xruyswR+PzaaFwbS+xM6nTznDrRaLXrI3PgegdsKLsvtjmZqfFVkObx9Htzbm90g
ib3GtU6CfjFgpk2o9/zJ4pnr9OLDw4UjhrUvaX03yKZfuMf/HCTzDyISGZJmj1GJqmgqNDeLh1gG
7w5yfowERmnRw+SzwRO/a2ERBx+g6PZQJ3DHbynU/KoKlQEzNNZF/Q5QGIn0i+7GTFY4bsfAjX3o
yNvVjvDSxiqKueLCGtZSH7fpWes8kF7nsb7cRSmlDyUPlkcNLwxr8vwdYaCzbxEWqSXj2LUKN46+
987QFnjdMlmsyshK2JXjzkAHekdDt9uOI4R5CdBJrUkrJ2sCf/4oOU4IgrN6ml/SJ54/HFL08LeB
mSSLRlr9zD/y0g3SAbhrEQqEfnjisrRkloulPjDSvNC8lPCqVGOcm77Gxs6j4X3KHJer2JMGN50T
G4lPdqw12i1+ZwJCkyjsynNULZPC2GUZPDgVXZZinISzakK72LedE4RDRw2AC2QdS697KeHkGdC1
6M78yUL75t7bchXdxj25QxWCWfz2IDR2kYy5UJTmEgAYreot2bK0258YCB74DwSJ1dA4gclFqo86
Oy0KYkpCC4q0tNa/yMVXoSLYA2hMeGzS/7yMOd0edhBOKWMXZ6HOhzlkZvMDeUWO7DdZedJqawVc
JSz1TQrTXOPK5Ih8TfKwnfLEzyO9d3x+E01cs9xQnrO984aO0CTXep7UTuHCnhOA2/qBk31jv9ef
GS2G4PdGlrngOvd+juZ9TZBApb37xBqlaoFrIXocqg6HTZwdzLfRNsjGPFZOAKoqFZYXvvv9KJbE
aVMi5XzrmW+irZ5ZedTtIOMu92WF+p+XoR4be/mUv5/mtYeuMCM/vp3XjADyCyBHV3dpzVUHC0ae
TprARtOg5q9jxw7OTsEKXrdt6dg4kKhrgcc8MHPoTFVJfHb5D5mtSboed62Hrzug5Wg8q9fRlpF3
uUy+gu2Rvfj8H65bQKV8XkhML2tfsvpacAMCt9j5RJ2Pfo4Z85OerQnRtQZzPu3ud4eVkDgd3kY/
XLXCbkXTiNcnGHuxfBu4mocqEduA3fARpe94ZiIxMM+EPnswmnlBZK93BCrk8qpTnPKxcDefdtxc
j55d51VbjLG9f3DOf6Kz/ftyIyDUb1BtV4GZd6Y12FR1XIbJpa68Alx6ECHq7IC3WMXUt8gc8Tr0
hfLm9JFaRED0Y0PGgh4JeiwmTdWiPKth3/9rVH+SJwRhZ65hDhim0vM2LRQ0rBalDEV8hF+nNaBT
9s7/2YrUYJzE+oh01vRV/RKC02B1Rma4qiDsCyRIKDmBPXf0hkaoDMGL7ZZuV+hTnRiho3XvWr2i
8PruuLwFnPG8gog+dC1KxedCIFp3Wh44cHoGtP7j9MpE1LBnntxlYnAXC1BLyrWeq8GWT4EMjY7U
1X4FrZEEgWgKXLDvktQhFoFpqDlfHw7du1MwuMs1xgP5bQ2X6Jvhr0Le5oEkaPi46kDTXfheSxzW
NfPtlTAkGYtEUe0zqtQAm8YR6Tp12P4FlkecajWglJwq4aSAso5lSOTKdCbl0aQ1sIgbQSKdqWKM
KZKwjGgwgwYhH6U/inpx5jSrifE+hjSMjAWJenO7PhG1br1NpWRh1gKSxr/3LRVbxgsV6+8mqKu2
XgWwgP8cJMAzcM9TdhEPg0oMDJmxKQVR4DtcgDTsR9kmpp515dFqRyaVJKhMkNpQ69QRntwW1+jP
5hUXnzkF2Ftf3DnKh9ufUarTS0bVkQ7hmztex4T0W1f/vW8hb9gI98/z2M3ghASAvaX4lL5sYOzS
XcPy2FSngUYDCOL3gqY58PxGzSGwuSpLVz16z4ngAXqER1kwy9lAZAf1MBBDpZaAtlXGA+1fX80g
olIOzGLdtNoY4DmBdKrr6s/yER05MfHHXPpq0P0ztBIUYvUbI+tLlw1SKkskL8ShYoFeQeQoE7ff
/vPAH2gBbgwAkVyjYrDZokYbnxci1t9PKMriXxwik3WM0JYgIuWAEQ2ojir1XQa0LWaJc5209CZy
xRs9PZm2kVVcVg5tH/4/yJc/hBjHzd9shfVBJkobFJwT03sIZArYV8anPs9qkp2fFStRHSYnlNQB
45ipAhtx2CU0yZXYRexrd36ihcpMbUQYXnEvRyk8HpUyOid4UshWTBmAYseIO0YZCRPj1O39qZQT
FfxGRc0KATjmMDq9fgfFJ9410LoEYLmJHUrJwaA1jUXotKFgBszKFTQlC8BKV/kWN1Yn1URbmbax
NWurRgey3UloFDl3LE7LXYc0F5KNdeUYjib1jwwjYhNcEGNQSO5zLBsR5I/Vq5yGdnEoioAFvvxw
f9qgrcp+fBaFQd8VTDA/mQG3FfB9QuV/z3TA99EpcFV6lyMIJ0eGfXsbjN9+9rMhPUhubBQJsSCv
0wL2fM+a3c2djzfq1iA4TmRTlukIZldwMrcv7/3GwnNWnynCw0+NOUU8ManEc/ZHeqtQCymTWnNV
rpjOjal5QQEAr6wRoH9Dn66AGoXe+uV2A7RLG6mHQ9/+c3fFSiAoDo6DwFnkXOna8unyRYvwhk3R
idiNWD6FTq40QxenksQhajZZ7onZrULinE0+B2/nfsAVgdd0+tcgNEW7W2Y6lpfc5s7lnoHXaYhr
1VfOK6gylaQwoKGzG41u5I/TRArDjoc6VpA+Xg+r3j86w9Z5MdRozZ7CtKzACyXh5AxmKkhu5rLw
CMXMjusr/LJnVnXgadz5N2ropiy5cYxY18yiN20v14wptD0AOWnZxbFA5DNo5KO9PCNhA+ppioXL
W7mPXh6TT8O368iRlZdbB7kqf2boUSkZiB0bBqQMRqVpHcjHs/MaBZX9JSZMCNDdO1/l4pvhYusg
Dco9AKikN3UJa6IuORkxpUXWfN8Ik7x2wl8UexI772XKzk0p73JKsArkQeTQCEkNjvU4y1/pijOz
4qKq1EGbwGefcuXXsNxDNGPSgtcRD2ZgSPPvKzoi+rhvG6W+YQxB64F/yi9y5wX5LsOLhS0vGkmS
DXRmpArO2eqM//8Z7m05Hiwg0hBbNjZDffrpfSuueWvZDwQwQ6iAaFaRMCirec7uCRjBasQbk/aD
hxoQWUgzG3aBmshLcOk15mswDDLvrE+eWUrOxDMQ55PPwo6lldIGlm0+vbMYgvr7oXtIs7AnNgpH
9ipuuZPhya0h5ivCITH99ZALdR8vN3CAs5J7pX3nf4PnFmLc+yvTcmCC7LmqzwokqnKXS5y1lwXR
kx3a/3XbINjds663sayM2KrUTeYyFjAgf/E4gaSuMx0HbaD0Ow0kr3bxkUOLZDNSUeb3zejPv8wI
xdZ7cVMET4Jvb4mTeOKxc9yNZbE7/8pJ3MVXxc7vabeF3w+UrrOHoVIVEvBVJ7RAJen8uxMdPH9N
pRQ8hqSUXBwjXtiUpGFCVWwXo3rUcsMmliNiKHihJWCLs9fA9Lif/1K2wy9cFROhs7ztWK14o49o
r2ccph+2zoY3JV6OxG/2jYQYd89xx8uqKFlxuZw/7qbXivIt986RddWpO3Mch+E7olBAYCmJfyb2
Ibt9IFXq/lsHWzCqoM8cXzF2S7kCLc+au9QvcXOqcVIb8WXZXrRx+KCF+YQ9JA70wylH/zuk5FLJ
5G4oi1LmjsVXz7XFZmp+7oSViRN3Ot+psMJEvKlZOZGBI+t7NGOjes2gV5DPbAsSyu3f5V7A4Mak
+2Iox+rnaKJcBK03ENJUio1FwBpO0Ym5QnmDiIKPKwM9BOSWcSqZAixNMysr/gLADuXX0tLboFv9
GHY/dXGp3HSfoWkoPgYtajsbAFCwrVpGDgmcZvoHf50Rb8g3t7YcgKZl5JfthT2wFKAHERcxYhjK
gcvDh9e/DHhKa6iUFnDtlte3nIUw4HlYUKmwv93W1r8v7bn13a49LOQzzDb531hEuOcyNrcP2IPP
VDRzv2bWaz0I5K2P+le/2k47tqMjYuMwIoGqwcZAFbyvBEC3fjsHcU2GnuhxwtslwZYIMxS3UDah
4EWKJ/V6ma4yo53Fm8AFFXgn2DztP9k206yCuJ7WYletZyosJUtT9JNKJQVxk2Ch8JZLuwNnrfJj
iQW3Awuukzvq9wErxfY3Xvos7vsqdycG1ECby6GjNNXvnyE+B1SH9gpnr91Jlrg3TI2M72RUNDxd
fp77B3TKf+6yl7xDESmLwhMnMh0EB5IExyPnjawret5NrXxiPVp1OOri+ynvOZ+VqnODp18fRmxM
z5paWJC4+KoF+g4VBeDlzXHGmsXbuy36Zfq5vTaE60V2rasLQ4B59FU4zzpvO+BxeBGKA+hVxWSR
VJksQL8UuIHs557elchgX9BNdDp5mmoR6xE0J0mHqmbqRgvwRO9mQt47PL6pKINWS1mLAiheQ1Y9
XubFbO/rRpkd9xggOEhSxk/jjEzGS1gvO8+Ep/rgdJWWJA+Q/yrlFOx1J/BjG1Vmdw51+Rk25D7M
UM2kxx5VaPyS0g7EF9WAmdvjKTfeWxsl/GOG2jussddEJ3l0LMjQMq2bo2kV/jopBW7bvc4/XwLI
EdBL9Lam6LdQAddcEHxxrnL5oOePTBk2XHC7jppxsBv2MRVsBJg1N1c8OEQjjMOegAB3xpo+dTVx
0QgRwC8dq5OYRAxPJKl89RaToy8KazhFObM8Fz4EtJlWznhXYeXktFDZr2RisCdMsFFZsWYn9CsF
gaofKO1AivuMMRda+JfoLMGEJvucMfnHkTdTO0u4U8ExBN4GbM7R3BQtghL3wjtxbnXO4A2pQulZ
ANTa/zDL8RNjGFPoyTY7CDAO3t2qGVXncWvTJke1EaIQLQKIT39Y464JWrEHft2obAqxdE+YeTaJ
FIgt+AfRCBBY846Q/9T/ZkiGidqvfXJLMBr3qtpxMc7hxza/yWIbwi9Em0mbnkiTxgNXA7Hf7Itx
zPgZklkSRZQHgiNXeZJMofvfN1UfRGBL5qjutEYcAkMUUoN2xfku0NizDOHTmfZ1fegaTVe014g1
N9GGspYs5gJuc4B1/JFNvD6dZUpDWxlRABaa3MaqhVaJnuAturLjFwrICaQmuR7PrElV0pxYKvfr
vteXvtoQ4mMYmRe28V5I4lKZJHjG1uIQ2/ejaLXwpsqDZeZanPW1lSOFRmgu0PdqmUg0VQCmxhID
JclYG0qFQPoRTOhoPyjAsgr325LmxLO289q8uCSwC1HwtLU5mPA83OxIOElJuTz21HpNP1nMqRLg
OUsjBRDaf7Lnt27241I/fWsOIfyzP2fjeT9AAX+wp3/eXSWh2iaNBv21P7Jr1x2T7wb7V1JBuYfO
TfBfG5pWNTqD8YnerfY0/tJmxtqHxIW27z3lKJKhfir2LiUPakQxDsf+7xNrPR3SddJCkydgA6k2
uH+tUKFzfsF5fFodLRzwbnSU1JqzCfpzrs1PFq7EAwitmfjK891suyFugMeeYyA13oWhRaMOxY3Q
mN9aGTHAM0e+aPoHh5mOfT6aU1hTCiBDtYlH2XYcBvjAKE9kF7vNsNdGkeCwiviE+gSHbw8HmDkp
3BI/YLqPjNeshpoPW+13w37or+C7jRrxv78uweLW5q3xeLfPYx7rWDSAD+YHy3ubFIYyE+bLKkSG
/HKrd6RQnFDrQtWDkqe7qaUp79XnR4pWj9DZRMXY7up3z2D8Mhvv1Zlgaa7S/Az9ToovoKJCaZGY
8Y1gDQ3nYZVs8lSVy8XUjnIHb0FBd1p9rDwP13SUi2sSHeRSTt7XQlya0zvLOo30uVnLhi7RZBts
S+pKeawh3/dTBzEaJRcSVqyg9hjCstqgwo2/iB/lI1kS0C2WkFp5r+obexMPQojvyGh/8GZF4sWs
YFeDF7oViyV01V+Y35qem9gkU5WXWNNChi+l/0Jiwhw9dN1WOrDhskTiCDThRtfk2fR/qGVjnY2c
RO6ONY18VF939ZcsjGzkR3KMM20XGai/5A5SfcqmRtfvJiBANFwcTMFuZsclw8GikLINfUnXgZvj
JtJs3UfRMsUvIHU2P1WGDCz7XStRskm7+4Av26hgMusXeh/LKDaal6jclcV0mLju+mpXaV/+HcEt
UEgV4lFFC4eprkAW7inJ689mI4z3owPfNHgEnbD0epEbFORttVikDa5y3BEhxSk+Pevdv88jxv8M
Ii60PKa8KSZZ5ckvtHsA8pA8L6lm6GfPYJ0fZYkeILJKGtEHnMDrxCc1vQj3f71gt8m/ty8D+366
Hf/cjj6PDS2soTKILYV4c+/f111bfxRmYrD9XoTQTywJKpC7Iic+TQutCoDPpPj6spvE/QHIJa2D
fG0+kX/CX3aMRdkmtHMsz4GaLi/8CzoEwZ5djxfbInFEuhuPXlUKGWFqML8qmheDdqrkDN9jUQX+
3goDLeu0oWA7Bmx4Gcd/zdvL1YBw4JJThI8OEpMy/Pa3YMJqSi8SehCU7K6nsAw9h8zu4VShB4zp
+V+m1fUKWX+2wn4qeV/lTWFiwZqvzDZZQ2ZHZCgTvaZtnaYRhWx+KXzQe2s8VWRCBzCW8r/Vvetk
sQZM2razbQ98kEfltrPn/qzgMKG5DJ4F7ilR5C2kITsCO10ofShdtfmL1V7vaWiegDjIkDSnnYZV
0bHLUfoZADtW2c4fMWpaiH+gt0KnHYoNn+HQjsnypZeW3YkJcbABsHhBMjOrIJcign6iUqBv35IM
b/T/fs7KtdVBis76KkfPwRhnbWhJdtLYduLQ0pPgT94R/zBfYzo9Pz8N/0I6j9U3rmDfDwPUe8Y9
Yc9dE+BIuy9F//zq7x73tnysge96YGK8S++moNlrns8ilntW9wvxfTYhDLM3Q+sGBq9Efu1UzuHj
svyG4smYm5oL0dTZvT2i13PxGxdJHhKvsUrjH1r5ALPsXQeiIei1rEUQVP+opqFGIdZ8KDrh4kPI
ZpRlxKMlUr36Owr3Bat7J1TCDXnn7xd4uYSQTLLf6Igx7kN+JTRZ9WJ7EgwJEioq8AisJgoymRqo
TOieP7ODJa4q63XQAS5Pgmn1xUQyTsNDIMA/m8r2UGuQLe0jvmIjNyllyjyweAhExeVaLigflnGk
E9SQoL5gzSnXfpDdLQriNeR19sAsxamEJhtqBi14dF7SuFtu54Jl+HEfw8J/e8iJZiHq9PkVkGZ7
L3kdpTIPZ5DSc9LKKTglJLJ3GhS+MbL2PXHLyFQXZRX+z/6ws25kf8sdfsJGvozek0rBJkFxsM2x
liqXM5eQm1PA/lsfEM5XO43qSoykDOZlKJvK86MTltAYMmlizzemTT6JURptz5trQHJDoj4UPTJ4
2cBnrkKWEMEDfjLBtjHg9ErO/9nE/AjFUFCcAwsmndJ2SwS0r8M7fhq87P0yajLV/mMWjdhcEUQg
yq7DNlk6HSSoepGSV3+7162LODdw5IsgaybnJ4xTOe/lDGplN+hXUoEaE5Fga7CzYRZScLJNv+y/
aLCQ42mjjVHYLTGDf0+0LUQZbxdWA9x8xr1egDKjBCH+uRDjIbn9caMhUHWDgUC/38FxZwHvpbHL
4PehyUKFm1jyaInTMnQw4U2ElkIwdqy/RuSAW4rdQvNk6FZaxK7HgJ89V8XM9SRisgjsPfTtlwFA
XK0Ch4wfWAN2sPLuWjMEmdGvOiJvtUjPvwrWaZn0VEXF3eL+uFrvfXEKtpeImddAd8Iw+tJXJ/bU
MZNVMvXGrZUT6El+yOgU9MVsT1BKrYGGf7m9onaM/VmvyEMVr+a+tvGx5sblkhaH/ReCUJeQq6NZ
NdxvYEMqZ8MPGiire1Ie0EG+hN+ywxRPQh3DsV4H7JSvVsPOY363yiC+UUy2Ss6xShRoES5ZwZhF
ElPlZQl6OoDvypmh61+XlPEnB9b8CVtoBwJSEChw62VfVdzPF/G+oMNSJlh8Og3HdNZQ5areOsUW
GbMBGePDwSysWtAA8VB/RkCuoV5P2OyeR04doyzX4IfytUo2cGxDVDIpPiS9exRlMRRGbRny9MtA
ga1j1gxmOQi9g0oU9PqLfRWetXPUqyV3lBHXpvm4gaXQpsYzgG1VSeQkxY65KBEQnMBBjPG5gvvw
ZTp16BSlBtT2XKY1050TmmaiJ4InN+rN0j/vqdEqDH5APHUDbDvtVxv0ep35Ipo7DD0NbHSDlpq2
9sC9NywEbCKoJLHGs3sa6BWzZ6m5gie5X+RvyzUYbBvr/3jSe3dH9PidfLDaAPgAdkLhwK5eY1qn
wr3BVkVE/1028X2cIyCfDsmFGxd5nmj4V50q/DO2/rgGRf5NJAaimqiYLzbt7AYkp3rd6uwimyS1
92PXekDbGxApF5do99r7nEY7SCgNiRAaF68xtL0clQHApDePFse9l0oGuAIrxO/uLwoqOGnmVwd5
IWNtM1nMW9+hG3w31UYniThCy0n04Upqc5fdXNqGB5cOMQtQGZ6xWYTPBCwE0KWlsB9Zn3FmBGRj
FgS7/YOqnMuaeXg+gFFUSFCz3SrzhkSBY6ekAZ3tTy0ZVN9/8yMeNFakbwuh9ypA/Q6gc49oE/7N
QZQm32SnCdhxV1goLMUKcNQMmbHctdb3rzZGI3xk9OPorEmLzeIoPjAsVaTvnRXECNz6t+GLbptj
a8/VoVkphGoqB2/DJVoqYMPOoh2fO/hQ8JLRQxYbi3ajouaU4qyNDrtK1KpjCQBYxldkV79ombOE
/kyA1bz5rSPL+60cEnHK/8FMS2ZGg/E/r4puipqBTcpkhBDvlzyxHd+iK6QhbDvScuBZvGPm8wF/
fgQGbLuWghUF7E200/Evll9zqKsp63f8+4HCJ9z3qdiZ9wRvoJYbMPLeOx0TU0Lr/TEW+gPZ1tIj
/evbtnXZ1Nh9p4+GlaTHxEKwPmILhNUL6k36Ygi/OsxWXQglmJaE13+4DE6TV8W1WSrlLZJK3lqB
s2g2Rz4sbgtgIGZJ+z60uTVtCJ0RkiOmznG64JMKE5HOM7aAMkTReBS3oq5GaMLUQjblVLKdrUuH
0iNWbPy9+0CPsuiLzaQy0yfF8vyVVtUQBpEA4J1P6HmDzeq/F1iFJBiZgQHbpfwf1JLTsM+RBSlD
sQfKzoxV/flOQf4Bo8PqTH+Gh1/zO/0gbgmpNhfF0EFnJkYeBM8HWH4jdl5eb+qRSZ1UoLteBSH/
XPR5AfLyzNevaKspLBxtyTn9CGO+R8I6WptRNmb2GvotuK2EAp+jw9ijJQiMyRMBGBJ5jcA/JjQm
W5zUjYDX0JkCXmse0fRRgOOMJgOdQ1Q54vo39Oox7FTqkWtEgziWV55CNXTU02lLqPuf6NxMts59
GxBTZ8AYAirMmEXp33lQpdwoMpBty4uFxPM3Ap6ng5qiZmU01DI1ZnOSY2R762F8MFnvooFdnbxf
1QCKs6uop91YtbcRVrvnP8F4DCwdUjhHTEBX2FhGE2uhsLBsgh3gXzxF7LRICfof0oydSf6vBKhy
v0cE9EV/4q1C0FNdfjq8ML7fjaPsKfj62aXstFV/B6jfoCY6iyAEi7ZCYr9YkIpKcNxVzuzXQ4Db
vPC0e6QJ51KWS/dPOv5+L97P36obuBHnXyKaepsCJdGCu0DmD2Vc07nRXM8s2ISr/V7Q9jsSLfWO
aj86wbpREXm7jIZq8IK1xRj8wUQvX3sCfdYYtqdHVRAAWucrMKVetE+mTkybR6bZj+5lh7eC80YD
LRg2Q41slWrReHUCMFzHmm7XmxA49cMe/w3wFAW9Q+cPvhgJ9zJIBos+c49faFebz4OfPmWLFSIJ
8hLfyr7vG4KvWVQMb5YhiKEdCEkMJSPfCrGVX9xN4LX5tLpPC3BDnKKWQdSxzyjQECza2wcipe+9
BYKfFfADYZK0tnSBHV9ZAWj+m8s9y1Xnl1FZyDNXH3GlidSdxuDXrh6tMV2V4r7+5rpScAlelrFE
SNHYNr6ZNClekWLF6hascv/3Rbjwkpus17MzMhySiBvMcX3V9S3/g0SxMB15T9et7h0ohutcV3le
P0ST+d4GLHevEqhJ4SixMg+VJbqB+9794bSRIqZL2L8exl8kGUvdoH0ydYHRxlTjx8TkRWYyp8Qi
0MzlUdBZeEOUzlH5+RK7BDpgt/23lR3CzoLFF+gOlmj6y/Zsy2YfHOunm13SnRN2BeX/LX332R2x
0uL2XrRGZOjB3dPBtct3WeQV7UsmleATvAMy7PyohkwNPwcaaE6MI9TbrEQOVcQcxn4yVgNtCIYz
HzjQNkrdgd6y0AYNij4WtePnKq+6KONpwX0N2lMA5TfRiPS82GqcLOlCgZFo7tyEq7dtbfsKUzin
E0DH6SqthLoTAvhdlzzlxyYBiLnA0HWLXOKjoYhYOQZODylnnBoKVkrMfCWZoXTmrGU+7kgTO0ES
2cDttdOXJYIYTih7uny7h7UsNJz1dLW+pSTKCG7M6vt+j486RY2cgjtV5DzIaqbTJFZt2u9p5Ecc
C9FmYzaOok/3g2i4myBW96c3fQ70sdwNg9IYTvDift5dUXtZHAvdAICyc54SBYGyRxOKteHVV99y
hvKs5iGNeykLawge7c5HAmufJDdFWXQ37HPpJgvqcT8MHgvOO//hlQo85FEV9DFtm5p5rAJ6HvUb
02pefV7kWh77LHvfgDArocegdoWyU/+JcQ+ELM5E0C1vgTBzRuKef1GKyVzZTBJsOg8V55EFxWgt
tCC2RMApz1ytVRCaS2LTNKADeOr37XO/ts4tnSQOLuY3SPXBC75io4agW05vn/poGd4MlMYUQFID
01CtzSOG2TVLsitysVJ6gQQuGbI62oknw2ZbLRTGK4NDg6u23B7rbaIhESQoOIg53b8v+dmbmkGW
eNuhUp60ukL11dE0as0r+cNbehhSXMrnevLzCyVAnJSkk3+ffcBwz9HjZ5LOEKhSyG5bvYzcN+6o
Zk/i1Gh61cW956/ZFwrDYtWmYvq6MJyfo0DIRK4KCENIWXOY6ALFAB40g1tifgUhafZz8Jqwr22b
rhQT3XRMw4v5VaK4BhXgUP5ZVnQVQsTXmr7oheEwDuqCvodnCWbOttOdb61X/fJSW16J84dxsDZo
v8YBIsKxGrALLPVDNrKbXiqodrZfwq5//wLpBGNQ682OQifM4lMLEkgOcixvk7nouNihaOdZYf/O
W9txUtsfoJHfGniYV/Vz+sQkNKFflACMjr+T54N8tyZsNDUK3Igis/7N/kK8WsPCukLlHuuHiO0K
NjcEHjY+pmN9gCQD5yeN/SqJuDSauXHFrXfLn6q9rVXIpQ7rycXmSwvX+pP/2o7blcxJ4NWDd0py
uJgiIeLRDHlQV4tw0Z8O5ro2jR6TZ08QCa/TbiHZ1IDGkg2qYIRlnqdAuNA2Dweljbj8/bFf7zXP
7K1h7vCFcvkOCpu9nSoZeXfCFAGHS/W92bXSXkHB/Eotn9F3kq7pBb66fXbgom3j9P5UQU0Y4OMJ
s2jJGDAW9giqTGzAbFg7xpwtlF8CuGpQxcgoIp5GxLp0Ig/qmHYzrOC58X5Ja9cqzT2elxMt/fIM
TD1Q6RHiXLa1Uxq0RNdwiKeSbfjGHY3XovmWAY4+B+f2F37WjsZaAjp4QDu6kyJb6GwuQb+NhmWo
6kf2WI35lcrPu9ilztVP5uLldL2G8VD6vya4C73yv7IyGao0Czjzf+6OHjazE5NWxv06b3qHsqyz
Zz9QeM+nr+P8h7FshFZsIMvfd8ed2azdIbzPBuA4nkieLq/hyaL50PnUEoNGHMLO/WD1KCnmxRuE
f+P1wDNO8/ciMkcgtcKzOY2vYyRDfzXiaR0g3DxUv+y0tiSCl3tOSq7SBAOw1arLlyBXCbhYtjyk
0ak7FisRT1PONIrfyUjA+AW/00JQOCuoqnTzQPPvtqPif73XYlsTKRbDCoqHMdZAIQ1wfvj6NjON
ZR03orryQpOs04mAiiQpmr2THiiX12bYZMaoVzvGOVAJRqp1x1NinMY0HjkKEZmGqt6MdHUjSZ3S
LIpgzD0AfAjkreUhAyXoPxD/MkcPwwgB7geunmBJEU+hlFoueiaRlHeO/a6Q6LEr5kEEdWHHNvSt
0kBxDCbLX0Uj5IkF8tMbJNDOpYNcn1KVsDpbRKEgF9WJ0CbmfCBKlfp2qk97Yikdn00BytTSNcLO
WGSUyRx6lX/klK2s1zkkPkDQJn2r8LieXy4D9t93+9Wth9Ir8iD3piz5GCFORDsmTZmaBJIQMypX
gjuYb5YNCMwg/hjd1+FGKMc4NsONE6VXwVN/OuQG2FBT2kIXeZnar41sxjU1GdVXN2xRXWjqlW2v
9lRrc1pAleXBF43Q6nxHUm6ibly8CKqxVOGvEG/8sFIdV559vA9VKM1eEYR2eU/LFmWWTCYuSVJk
0g+U1W+YhcskHAv8wx6t7o+U1kIM22PBzd6Ag5iOaosJPkZ6JiJhXIMEnyERjQAfPHhh5tNwJgfP
zm9mwhSRiqSH9yuT7Dwnl//EqT6Xx03lWTqUUrgufQR2wZOe+epcgVDWsuQdnShUj9CC3jTY9J4M
FYuMbpLRDIa/qguEh+hQVevUl2ekztjWd4KHx9BJuDcRx9CtXpEHacXUdu2G2GuU4WXEUKo0jWfo
8FPELGl533NTSOL9Di5uaUiG3iEQfzZubqk5ZutxMJCXV5tGLGGYX9ifSnlZhKaDNnkEDgiF3mWN
8xbgnGppNzdfUbFqjxCku06vB0z0lHOR4jXKjLA39TnvvFWgCLfCJ4vjKgH3kMJTUaamATWpHjM4
Xn8vUdOxs7577IjPAD3v3k/NJH3J9wM6AgffotvtgTEbtZh22InNdeLcaVbjC50HHKqYq3am8lnr
5vk4l/lzXwEO/xvFjXnDstkKMMk8g7PXeMHGD3QyENVhZQ12Mz+JcKhafROgD9kBvjAjaLL/bbIN
kuGAl84I1TKlTBesNXHj6g8Y4QCehWPp3T9IGksdeKIX33aC8J6iUi3JbXgZtlt+ZC9YnxqmKHMO
D3PtdIiSSVITxIv5TujBduo8+ZJ3cERwxUr8UZgv7twwoEwaHk2KKN5wOA7QSKPO687sl1BubCgw
YTiKwIAdNa3cLG1DFlk+JbfwWDpHieWywUggKf7163MHr8EPOogNSvIalE2l8EEyk8Kz6UIx+Te/
iiD3S67dauIAX9Iz0iI2h3+8AMArFybnUFvEpruxAwQBQozMdGk2iVX+jLJbN1vJQxDKCpGo/m9T
mODgih999doKcWjlDIvZvCtaod5OZ+cyVX5TzsrnrFf4FRa+KFoG9s5SNVP0U0+AZ7UeXyrC7EP6
qY1xuo6xY2psmhD1SEtpa6nCO3iOYy4s/TiPXSXC8Xw5v9AqB79849kDN4i1EjZJKKYZzL2fHZfu
O+5sGBggElo0Du/iv3Bws9LSEmVqNPUqETLz6b1rSo3jeQYckRhg4HsxxXgBFL/XZ7q12P4CsQoi
kX7UAOZOjb2ZnG2dy3JcDLm4RU2wRRyzcUm2nmNyTvnu/fuNFA+YfIIlvx1/QNvk5Hw0+Pl53jfk
HesW0h+ELre1Wm0qJ4uICLzdyYgwSOq/3wlfXXoLQmGCKaniTGHs5Ph6e71njFgPYXaI5I1gY0FM
0A8jkt1ucWukPRVpxIOlKEOcpwgQypfG/ge0aoe5gXamE7THD1eNLAWi8AwYwiHZZf6H6MzrOY0M
M/8LkaO6I9W1EFXkvGcDQCUcvx8UvTyfaJAo2c7hPlWqpt9mk2COwonorizRAIiNmaxs5JDAgpPA
gGzhXh3zrIKs05jVA7tyfE5PeMeVmedbo+yoKZ5xUW7i5JPoraqEJWVOloJ54vYONTlLkJk4Qy+L
dVv4B670OmPyGMYYZfRUSJXkJTpqA+zI4YPCvI0Y0YiteciSnKPPF4sIk0KuZi09hTrALY0Srb+D
Yk0lS5vPbUgfTXpO7jnM8hvehuRn8snWDUpLJ+Xuw940+kITZ33uKXMqB22hcCoN8V/1Os+LfyuG
wqbnk0zxRzwx3FdKsqpCdXsqb3wf1ugteq56nfDve6pnF34NQ5Be5qqtXxladQTQV9u/SBotIBtU
EkIBgIXyBVzxrhlc+ruRWDD1zqUqSVzZV4Lftufp+NEeVz2/s8N9ZDjyFHllMUsfd86k5rmNVfQ+
tfNa+n9aqtR2dJ8r/Q+co/A7ShWbzrl/PFb1vuftXK/qHMn8phsVJdMQmbDYttFAU++S0Oof+SIO
ZtUOeb/9fBylrTH+IB496de03SetpaNzYd+4giLlZRlGhJxlFEI6fbMdx9vy+P7sVRIwgqQVDFda
kVnO31k9D2yABdU1EWjvuRVOy0FCyWLxUD53vmjk69v5Di8e3ndvkuLI0m2DfJZhK9E2ttQ0hRGj
7FTj33AyjaAVqQpDFBi4UWNhK/lMMrr0y9CnmPqt6i/DOZwJtXcLdCjozLCKF9pWP0Pj1Vwz/fB2
+tXAwXvcnRLjzUdxRn73nNT4NbFEkGH5JDttRkjzK5hGb36JYpp+li9o8vIzEyVSFjml865BSERP
9m61SodTu3vQx5/1xFz5F9ZlOrnpWx0SGw4XezFlmvy6/pX+aVgoNfcL42ykQ6a8tBoLurxSyEK9
jQDxHUjI5p0RocWcVkH3VgiN05lhEWaeHq2480gvoaacDQpA9lvaONZ9YNRw8RWs/t5LRWHn3Glh
9/oQUAbF1CZ8BWXrUd0QNsZ9jWdeFjD7dqx4TSO49QwKCcX+eDQDX0k/sqF+mChyvK/6L9JKLKA1
9LJvFJ9qpQ83uAS0p0Bcszw4VxzV9hQNz+n51ZgvwOXjhN795UyU6bavRzNUIJOmuaFxf9yMjAQy
Eg5ne8NnB0zlojL2YJqcx0cyobjL/carW1q+8PfoO2NR+4VPTH9lzVjFmknRZi/I+X8HXuDD9Y6k
bD6s5DuBpSHB31GF8f2BX+3WPFkU5bXgXm0M8CV+0eKSTQu15zHgKbfO7fLvC3bEjNEsp/TsZuCg
RvseOxwZ53p1ux2/QasB6QnJ39qlPHBMRNMI43mQtBkIvFKmHEekCRaUxfAXkLNj+mpj42QNhxH1
rN0MpAHsddq6vxbn2Ns8BlHsSmfzcjFCG5Syl+6z9VBc4m7k2k0iL2RpctGE+5C6F1TUh7MhPWW7
VCPM/PBwn4GqZILpvD/wBVxyR+/Vz6MKRbkHwYMuwfigl6+H0GqCobjTUCBdC1d0cBAtDub28K7i
Z2a6+kgAlUR467znrRYNmsCfTztR1ONsdy4yKPe8sduzMH/gtrevK+rcrwFSNJk2gLxTbsGty87b
P/o4fseSQDAEC9Of64VEXGmD/DdFee0TmDTOvt3aswIww8+LUCwC79bzo5dm986hoVHeB/+P0+X/
UoWLy/iGdV35NBLFCgpU1QqInrcQv04eZOoprQB8mpKImZCQX89x2VX2De1RanqUwqRkOpe0cX0z
XZmgIzqFX7/hx84L15tnAXNvkgCYaFJvH5ZKITA63SoQjKQydwMYjtR0JKhDclxBF8GHR6kdCTYG
Q1b6JKDRYMDXO84wEVlE6+KibWUZE9oyF8K3HVaPKwN9GJXFh90PeyRvlHOrj/lNTt2UdmP5qsIY
om0y4Wpeui/T42SPKb+8c5vMXqZ6kelcwRLdb8j5g13LZznvIrJIAYURsNtwK8vZry0EgJKSG0Nl
OkiSOGRqmwZpHZkNFU4rsHh5IsGFe89KGumXN1ohpKuccUERJ1v0H/3E0uK9WtoB5PrR/qdtD6U7
vuipjmTiuAMFZP4qQ5QJjlCnWAe/EAtCh/yD+7mWXmPrfSTNRZV3+rrOjGti+hLEB+ArddC6CfzO
iK5NgPfWubapgWWeZDsnvOS1gGTgENNpUAz05ZdFGtlIpMZXtyHIxGwg4V9PotxFHE9Lr9oCspIm
SknA2rp9AWhKcjq/7MVwTGAeCgeB22vSO4b+wRZXNzRVz53D7uaJrzOZ4tSYmfmZDQCtcL7U+t3W
6Ee8enfpQWdpPdlYGCwSc8iHGKcB5fkqxmhe+iLI1SynBHQO/pFPEv830+3iLvKuZmKq/h1sB/tY
I3i+H+1W+EX+mAOwVEVR7whwmgr9XnmI2vR34Q4kITRKUSMrOzSYTj8RIbTRtJ3YAuLshejMrvlo
2HUHzpUdD0iIBNSPVKYTWdhZDHfe5rnyElvVt/NJn2h6LDR/Nfzij8rcU6kvIc/DzgZNintKZg53
MCwvldx7j+XPdXo3l9uanunppJCxv5perFqTD/3HIHPvy1k+aPU63y8dhX6kzWRzuwh56BlgyDjV
UggG4k2/7lp20T8YF6/agqtVrihYA+LYyJjLv5kSA8wgrZ8Wu5OGYK731zVwmk4Q8KVru77Bljpt
9P9i/nnYCrTZGRty2qpnA/OZPAMJ4F5CzZL4Qj7+2p1ne5UtA1FLwJm2EnGDkY/wOHv6RCRPOOqD
XCGQ5y7+vvroXzUpHdgBndzQ1apxnFOJfles49Wcu1b+BuOmo+banbYJ26YS4eLpSNYYBr8hs++d
Y8Kgbxu6zgb9wrYJQFjy8QnR1KE4X82auFCkmtcpLN/lMkSPjIMSc58xDRl6/b6h3vvLauVK2ums
hL5ZthepjQO1B5o/71HtzCweJtRWS6xr620Q2xKvdvvXewybwOfOATPNWwVCSfz+PhxJf5wKJELS
LFtoSTJqLV6IOfQPdx+W3jdFmAMEcmgeL+LlBsR89nJUJnB/OP+V2csAAPA/9We8rswAzjTaP1Cc
MkluS0K9pP41F+UP7PLfYcGvwYGv748lYHBkxPiA3GjCiLCv6nGwbqXXJ2f1KqaqLSe1WsucEcjE
gHoLbobAIZJrCx7t/A0ySZp6IEJPCHLR9LqI61vtIX4gEmWgKc4lrlNkTeZYhxGbW3cmdYt+ID3w
a1jcv7ZgxD83iKvE+hMh0idlD8gwsQT7E2+nnGROcSMSAlipAgY1o5Sheyz1tgpz5oc7skOmaRTZ
/IWXIc8eowROfcwSPoYyGzZ5pPFfTK6c10ccvlEufYbhqhl6kEjh51tjZQ8IIMWJEJb+hbPSdNP4
EvIB2154flv4m7It8M+drDGQ+Vcg9VZN9TJ6bshisb99H30Eg2NC4klWU6M963wC0AR11E462RR4
NrkVb3PN94U1qO1MoasOJEZ0Lpc6Yi1ojT6OTGEOsKNMomUSemc4ZJEcr/AwfwXGzC2qsC1ohf1e
50sGudAKQYHK7nD2nX8tDI8qHThV+jMzPx2xY/rIn1GVBy3LWshfGzZeXcemGPrY0oKuJ8HT1x1S
EkcAMNRDnvQQTC/DBlQx408gpqFvX0EJO2k1MMih7KhS9ROPca+pkdTPH/Lo/lAAN8RrdiTfIHTI
o4sPLuvz1kd1jU3GqWkuNZf+GRxuy7lpz7MlFanQKF4q4B2KZNm+x6R42c8o5MHCmaEW03wduUXk
iRMVwOim6ovwhHqc+63WMxBvJ17YSj3Q9pd4XjtK/O3ZegVqhH4UcCsqyTnMFVFUpFIcwhvIsK5x
oQG7+QlH+PVJOMOdtGP6iorhSSXXczCGz5cHKZcwJ6P9jZaOaBcnhJNKNO4qDi3KGU5gnT6iNM4H
viDuAzYlm6DjsmMHN+o5LzGbFqhz2TD1U1BI9F3xLgd3cYehL0sm42W+D0uuzwLifQSzAGSoCoJ5
lrvxBCbCqo7LPquyrTIQH+LdjybaqQyi2mF4lHCpzxJXrgIaLOKAjeYKG66/Mfo82bBcdtBcFKU6
0BRDXLWYthUvONackMX4/Dge1wzNC1hizNZrPuNP5zQ7ukygeK5d8qn7vqc0yw9aRA5/d9p07kJb
5yyKynv128BecajN7FwXxccm63X0//R+k3btXUbCEJTY9K2y5Lc+iRDXFIihuX3EvMbRBG9QDV9l
oUprfQHnvXKEbmczOVf6nU+xwSpPh7WqOysZzZ+eVutxli0UkrhoMKyYuF66CXJW/5/nwhhxBOgG
pMrwQRPeuq0WN38dhWSt07jccsC1gilpWvqFo2UxaKtsJyfljFq1gG4SMkKneU/aoLXOzHTyEF9+
F8P8mg39I41tLH37IzbTz/5VCvZ6GbAMk+cKfbq7S8WB8jpoJQpoP3g8JL25D9x+QKDnrazXamZO
bRHfdJoHjzHAYG8xHuj+LeFsK5oqszi+0Gp3U+Q+1YxZpToaRmk1iqcHyYRAeyb+UXSFHooqZz7E
lILHPfVf4cFfWmBPl+i+3XvdRsz0apmtpm7qJNhhkmMfpc6mYxG7iYxX1z/C3T9dmQycYBlzcRj/
UmGQO/9x63oKOc6d8S/m3/J8Z3Cn5Oe7sw0XZ4C01tH8gzaDR2fVwCGoUFH2On44VTqqjdlL/OSL
KcyLxRzq9F2nJElMDzFTefudQPlb3N3bp0lc75i7H9lo6UJvhVu7IY5c/QYkWegUt4EvVdtAXIJx
m1vyhj07kAHkSTgde9Eb10RJoTL0ALiufRaMYSrSWgk7U2BFqb8Fpe0n2iHQXsWgvujhcHG2MA0T
gouq99HrvFvsVw4R9RVKzDz5TkXoezJM+gYBPC+vTwSFY+cRVyuzIpLTtinogyO7NZ7zm3maMMuP
zX/DwqGqvjWoeKipLgj30rM6eu9NY5l36KS6NmxFW2ZPgh8D4VhzvpwayuNcuO1BMa77ZdPAHEg0
Dp3LY6oMgSfDO9n7Zcam3KPIhVlgQZhgwKaa0WzEoafsSIHcbF97Hs+Svv46DtDGyQsUEjvHJ7h7
RJs06lmp+WwZmoLcMxrrmwti9D62qoRS0FuyM1LE4xxunrsPEe2dr6p2yiMbM/66+xUWkwzgLC6i
7AyCWzsto7/EuEwIE+BuSf3uTehWBfX2TffxYk9TrLwRHlPiIKmuteZzunm1I0GkLwPwv4i6ApR5
WyEom+hRazprbDFWMMIfq0vnidQkvAxRF4Kt0+C3uI4ygiMfVQB1wVVa3Fy5CN62AAnp3Ma1ZUa8
CmlFEhilFUDf7IrtI8Weo7slyfw9smxwFzh2HUCP2BY1rF4TgN8O+c9CB5TrHwx/ZTx35JgGCXbQ
Krr0vaueEHmU7rtAiigdP29oS45I67jUaxxzSBE4gD6mMkyEvJLZqi4K1ePlNzfhVzkdocn+mkHV
QPYjof6wA59/eTn5D746+NVtBVp29aZ6dIYNlywJ9gUU48sbwgiw3kaS4IPBefzbeBGbfqMJi5dq
CEwwmN4PrIY+G3p1QdIagC1EjmFpStlDN3+K5hjxkDqMQNziqdtrZICyUUwHvZErHgiqeaw0XSnB
+XC3HovAqeqaTn/dl/Tr6bH4EFuZNwZdsaFuUtuCnccTogFWn4zY/bn6gp9CfnscH8JGPrFfYKNw
fGilsBbS89Pz43OhpKQ2zSEsKmo0jyJIJ6foSWTvFPORyE49HsHWX2OaDll9AkQz5sHzISZA8c3c
ESr4xsYLW9fKkAeoRoX8gSqc4g26Zp3n8GRREEdirrYIMKpULw8wZBVKS6fPTlPG+LIueWxOULFY
ThOdUVpt1oQoUDT4iA6qKD2/Xu5xvMXWV29nGwjjDCWbR8n28keS+WXucLPCGXhhfyilQT4sdMtp
7oJazFGSwHMTZ2wkbtKGEEZCaRa+nsDnjDVaNlZLzh2kpWrwJtjKftB9rru1Hrz1+A662CB7J2xH
oaVOPFmvohRcIzNZHYTAYU7SCY1CEbrNZpiCaVRsF69SjbzVP7Vs/N+5Jk32bbKZPMJ4C+F39u6x
vn+DzhTPItVQg/iIBJskC453clZWtFDNDFXBIhVNLjciMGu/POmI37oiupgmDiPeYAjZ9EGfZD7W
McjnbfHuvhVTYtDqJzp4IZjbQMxF45Ykc2+cNZ5kmOKt9Ys3rYz2dFKiQXPycEqjpv3yIazXtjJu
KEE4G/o0byp5wOff4AWqcpafz2DUNcXn5QOPA2llpXDyunSG49XPq1EfHo4YyPr40UqwMbN+ssTR
gqRHKVXf3kc9TwFXje4RtxE+m1f1JufaSCwhbeMxgLqHHz7GbnKDB1LMb/Osa2CTrXOqZmgUE9II
S+f61RoYRGNIoNHQc74YYNVXFj8WOgEVCyW9Qrinz27SnJ8B/av4ITkKgqjZdqE9UDqsVJ9BuS3S
Or/6mwg14tdIgZ/NRXoUh1GI/byRiGi7oZUKYo96arDnDeLZjuQzljuANdXquhEE58Tur6c9JHzV
ZtPFlEDztMicUk8r8dEsggfkBmxDLjNRrYZ6XLERt03/Gy6flDOK1D3imnKJzQFYItkFfeCFwR7H
TY2cge06nRZvvPFos174AMpRJIQl/+bkw1QpZdl8DU2U8GP1MbtI7C9QQxEualp8VcwExLZxOvvV
n/SRw203QOgJO7MX/phKXIq/y6ROxdXEpmMYoU8QxXvoHoXRzSbQeo4oQzBaSDaxHKFOP0n9OB1G
PnkEBFxNPgD4ixFxFHR9+mwrQ0Ho69uZS1YYAr2w9twKNBXx50CPKwholIR/X9eiGrNxvGwr0sWd
t9rewSVQyjiYV4H8E0pmUx7rFVUOvLsT+4ek5fxDfZKWRXo1QxaRl7OrtULv3Igj+GA7Dz49dKrg
uHTpfLya0F85hjv4cltg29j7TMm9zOanisGDxUAzkCXN1Pb+14IVsQfM1nTkKhEp9sKulQAMF6Gu
A+dfNziZuNz60vZtXAW3wgrfW2ervOChaEFe7LPNySppkkCiVOBIfon33HvKuz/q8uONyCMq3s0z
UOvjbgmvXVuOUihCh4ImXCVZtLin/5EHuWOHjjn3aZHgZ1pXIVcJvXkh2uAvTudHgVxn0P59eXoZ
L6i2QhLIAu7e6JbLHAwAlutvKMm/k8GcNGOeZ7tMOWECCkRpheyLavCShcuLONb/RBEH6DYtAHD8
FFz0b9IfdPddWGO+dFqigYFj4NBZk/+fuL/vC+xngLLZ8G81Yc+wHnXhrsdWkVEAwT5LfeVRO594
v01nDX7XgAhqharunfr+poZZ6dytPrYQKvvITVynVL4q9RtyTHmx6oXdBVJR+str9H+TcSjHAHRn
Wl/K5/kFUXIxcgXJk5wX/9MxGZw4tZQVZO5koQze8xDrm8iGVCTsJBfaPP49F/sW4bynFEFWq50N
nnE6ENNAF3iOx4nm4PzglAnTBFQpquqwOUuhYK/tbYmxTfC7AkBY2jCjyq+ELFEsjuofmHip9AYg
+VeCGTj+5ztd2++aI80DDVgZkLEcqeiOpavo+HYYS0BljYLYaEhminsyOIRd1GYS28pHCNYENZ2/
WsVa3dUoqUHai5iS9MU46EE3FKpG+UGLC+wYo2No/XdTjQPz1sGMMYecGXjdfhrTtJpWT/5RDaZO
Bw3rUvEAJMj/l/XX5dqRrfXomZeb3+xN50TLKceZsIP+cJYheB6jUSKoLIISZmD3BPNUUVWfh9hS
j+sSi9Y582glKBzgU3i43ENBMopH7iz46v89rGAv0HP23Uag3em7uc871ddRaC0wQXNqX4slwJaK
wRteV0FiNjVcGMyrHUjPTaOEmlbK9IiipLumROCuWWugdkGS880VI7R54K9hcFVeMPxTMDf46e16
S+w5JlHNgh5bTzNuFK1px6TsIm86TsBn4vHq7wD0mdCXi3TKmdsR4dP2M00xo0SWLmqId7rz0dby
J+3+3RkcPyI8daRVL5KbEuFmzZLw8UDrAWjvT781MFwsBU+LLfiTomP4U1tVMg7bswijASR01ynO
dCyIrIUxcADee4DoucXA9Qu97JhYdX1LbO5Q7/J/Rey0jXbEXHPsQPySfHKf6NpDaQTUK2IS/sKt
NCXn/ZfdZTi6ygiaaT1lUpgB9k6RgFdQcelpPdjFPTWkk3fAV+p1Fvg8DyM7p9uy9g42O3qqORLU
NyiZVTM0ISfNrpgUOOEXd902wfW/ULhYELWc3LMwE4YpZYW8dRo5fg38W5fHeZsCDQBcXBSUaBpn
FULgdL33lyTE33neXpP1prTEAgD7Ym1wsJR1HCTwdOVPEEpJvFaF672bzurydLDLk84zWds6nS23
K8eX4qRtfr9y5n6d28OtwO4f1wGvd6+XWLjW9uYHMLpCFPXqK8RPrprdt5Vxijdgm/T1dTEgZFiW
e3AEHjvdHKVOOPlONX79qj1W37W6QWsAsVn9ayHRLXWfTwSScHqXkjRSZc6VqLSX4tEFPBDlznzt
/2P5nNKzDHO68mXbICfvbx2CYE2l7nIc8Pc50WPkv6BnSEYIQEOfqTwqKtK+C3n7kBTcq5MhCcMS
DroWOpUgGLG3HJ1zFJP9bJZHdF5T98i2R/ORyqb8vKBS6EVjR/OkY/VP9/mTZKFCHkICxpkC7mSt
oOkAQeqR8Enw0Xin9uclGbx3rsVc7HbDXk5vnaykMxfAE5QHVASfAO6ZrHuY+Ex8ilgRa6IAtnbZ
QIiQoDDlNbyzd9aIRqfETaWZNEK8LW5F2loYApJxOiNp5RTCS9ovcnBw49atbMNMkykFDG8e5TeI
BuyLJ4kyb4m+jxLNGqUfXdIRPdD31KouI+1ueQBB0LbwlL9vswweZFCG6k2Ih3jvonkx3guzT/Or
YrBPyaY5WEj7NxIIZAK4Xy6KJTBhrgWEgyniLaMXvDx/d0CAXAw3Fz4plKVWUVdqLTZnPAEtfWWL
PwyLYWiPcQzeN2kJFI+epquWugqQw3bPrJbKQpNOKFXoFFC1Bi7IbpcCnFT+f03QkLB5hJxF647U
ne20BFkuHIyNHKcaV2Peyc3P4aQHwAAHecTqvYPQYpv+GHozcfuXNEBkf78ODvUxfJ+I4yTempOY
QayaXaC/tRYMzmqSLQpDLhfLLjTosHdaLZEVg2kTeXC2ZDPiuTz1Qza+W7K4kaxVbyGeFypQSPzG
5NEnDNlsnu3z3AVVEZWrCVTsNx+hkK/hZBULbiTMy3VM5EforU8Yx8wFGsohaoj1afuDOcmAzoaj
vj4aOqj4TcTU3+/PWkIYfX5KCSyfQs77ZWVcNVOwqkfEhiHkTh+F2SHEx9FyKXzu122jnBMkQ1ce
lEKyHqmfH5MvSpGe0mZX6nHOHZZEjqM6cyBPekxPE5MuwbRxP3U9YmqLCplxj99sH1DJovOs+iei
GlmE58PLcr0tq7lCt9H+UotKOTDW4MOfm5Gb/BxehgnqXeXDDIBJG9inK0c4CvZZnLaHX0QHOvhR
DSYAxLkwxYT4r12K57RZFZ/WMPshmmryLZ8rlIk7jxmPht5fr85BRbWSSfQSFg93c02Cuxxb4DnT
0Hpkl774LWL1iJFtLXe/nNSTBsl4lkZqW3VzICXhIcASQf86z/Jwv2uAlWCi1T80hx1tejJD8c9W
mExsNvmFjEwyBWwEXynPew6hi5+PphluIgbU4i8mEFF5+flILdKrUS1iWPzCaswi6WjKd6/GFGiV
AxEnlLjp5c820fr6gfXe08z+FLg3ofp+37T9t8t52qMVcL/c7q+cInTiyZrj781o6U54UdHskxXk
kAExSxFYUVbt8J3G6uaXV6yoQNe5obfBmBxMhDSg+MwGRAE10NJrW/g4jm0m/KYpt3dVS45pnS93
SlJ21eHHgm25vYm8hVbDPF7fWcJxJcU5nu0oJf+6oYRVyNePAcOJmJXGaxh8WPd3CAAxKU3wS7qz
lGJofDXJlMoQDmEdu0G58dZaKSpFiqwZMYNz1X4f2R6Q7ddZKHZGHjTtFzoSkrz531niRrY2jC8H
njAgZ9zvvdYo6QqELMV6mEO9FdpgrLuYyj4xNp1BYEfuyKmsh9PSh6SC9hqUdDZ5pRHDiWMvEntP
8TI6EI8EVzw0wVaQXXZAGMlzUq/iUoX3tJqaP15bP+wkBNPxW1Qzct7A6rukazet4GhJIw/XbTH4
BFkAY/tkgA/YbmR/cYemhGR7hnsMbGJPv/BZZyk91KzsuT+yOyB16dPnZxpkyyoTFg2xX1IpKPy2
E+LKyEgGfP+bhHQF9L0WZIyVeas25QyVdKCxwphk/ecxEWqtOPoRQNXjaUFtOsmy2byyeaMgIijx
NZjZs2L+73f5LoimLtUXOgLvDsWh2u2t/RdyHy52QNF7MeI5XORyuJ13+2tu+lwVsBNuKTOFz0sY
I87PHnjd2n4zVYUQdsWx+uOTB6M/O3dWiayoLJq+HG8lTdGTNgGMuV6gupGu3deo0SR5tX4Pp7bR
gD1g0ifOV9qFjof5t9Bw3qXWTkXfiM4/CIQzZEjmNaip3SG4I8xb22N2FxSg+wUGNaA+XOH+Pnmo
dN86HC+cuBf3TyR8Zf6Z/KqSCHq6UfbPP1h7cW3x/9E/YZrw6TrmMgN+rGy8rzceBPJE1j509Dhd
5cLSZEejsE2Rxn7XJd0TV7ZSWa8Uw3salhGKzHCjZE2Jy/tCVoEFPxtsPlgg8cpuQjWMfU6PM1YK
PN4edK6xQJL7b/Zba4yu4KwrGCghtedHxASEAmRp9pJgiOwtqzp2MFMmE6Qkd29JpO5AQ+auUluo
G3kNmHEcQi3FCDhlucKNZs06Y235P4GteOxydRQPBsqpZHgDbiptGDiUCE9Zrvqrvqtca2EIUDfP
UM///lw9qbGZBZUuZUuxFPdmKCxYPa43pkKe1MsOtSfILluhvazJMYo9Q4Bf7mj9JGzLnKFK6xcC
THmOImpy8bKM6MngbPRkIWGCPKDnAFARFExh2oPszarX9jBLLIaEy3NEuQY7HMNQcUATNSztaKuq
ee2xOi1++uAQFLjVNyHhjaFf62h5J9IgJkSwWPnzrEEc/LgpzxgWocGgVjXeTymNj402RXTXCtum
wnwHhrQwcIqtBPuPKWqCot7o7RjX5BwU37wiR1hDCe5GFtarNFtiAZMN3L6PbaGVxs21Drqd67zo
MVEkHIQinEzmHXpke+WnrE3XVr3fkSjJ8vab+RFr+WGKjKQnl3FlfwURWJbcII08mugGtB9+f3sm
PI+AHrQCaEEyum050AhVgTrInzgL9YSvV5mK1eOha8q2A24qmtdr2A+t0LUs8175no+LLo3leQTD
8zH8TyHvugIN/xc1IxNzH5zWYHAx5JU/XDEdOkbGzOAGRikf/088qn37ReXPtX66j+QaPDSPHQqK
0f+Uni+BdgGCIw2ouHHmAJHbatuY9PJHwI01vPTYsNJsdWPeU6NF9GaSuR9td7Z3DsSqQUNivy4R
BZIznqp4FUrVAQdQPocDlv4m7AJIUaSR02ET2vSNnap/b0Sxm98SjA+xcr+Vx/mnHihjc8c7Lkfm
7hdRjpzNXCD6R61RIOs3beehA9kT3Dq4B/Tv4w+3mVLyxfqokwbANiChX5T8QMGrQTkyw9u2QldW
y3AHaZ8eeJHPZil/Fd8nRsoQhH2Slhj6qsesgynL6HolEPY11tO64GycYM5VrF62yg9gqfLYOtns
gi9BgZ1EaZ3/h9dmLO+wlbeJNVON3PaWh3YEgz2miMe5LovxMeunWo+DYDflsMCLu6OrcmCBfEro
OPF9a04Keuw2AHC6wA9BeZ1wmeiM2cwXK8kezSqv6kFNjUGvQfXRVQZV2cmtIXp3wT+FMVN8lBMa
bOO7ZJDiqYZG6tRJKg0/U/QLX3VWGYSdoE2K1MciItouuBCwbEO1HaLl+Y0xUJCgr87jkhQzBipd
PRDV0DFUoohukfWtJBFo+d8W7FIvdV3hhXTP14E1B0jyhe18ucIQkjTzoPjV5EoBigobRHf4xU/g
4x2rYf/KoBolwT+G8cVCq9yjRLIetAChHKuUFSOjI3uH/LBA+siPxP3Q8Wl7D9o567Qn6/qcwYMf
MYCsl91q7hYUG6xct4cIBhdBBgYjkgCqBPIFejhXRCgeri3BVgwD/El1v3Cczan1N9E/PgDOamB4
GX+JC7b45X9XGqok9qHsLBBOgD9X/suj7IX+QyPpQAs1T4+7zE/WNAffu1/lHLqnpidRU5kxZ/16
qlRCqiZzlGWLUpIIB/9yWS1VDOkf7sOMXtNGqq4VSihJiijgr91ElZl0jeiXMCKzRqMc3D+0+hMs
e+1DlE2pcKtdlQ3NEf7lMKXKDOADmn2oHVXThUDPqR8sbhPVaMh8O/M8o8hC7zXheyHlI3IyLQYO
ady4FqrAv047G8lBZYZcB2AvQWpe7lFEz82Fkzubao2ecndE+0MC6SZiO7vMckk5Uo8Ww8RDFXkl
/s7/qxuh+iRAAkzK7ezOKZI2Jguzue302OBX3WxHSV26yLNc9/r8Lmd54esyGw5dju1FrouFe9nx
ppaBf5tt021pE5yE5SKaO2o0RRTP8eWe87uLvi2cQmt7xfum8JZLAEzYXBvJeq8P+BOizClxnu8B
bcGwaBn8SEhDh3/g7RzIgbTuYN1FSPUJM2TiyRUo+X3WVcVFqBZbJGYvNCtpjOeeDSWsWl8lWaGU
akrjWdXHuJauzdN0e/dRzXTl5Ir6hZUXnpyjmxIO8DvpvcVnAFW9flxlBu9eNP2tHUx88VUxTAQp
mzT0aw8Of7xohMotyoS3NfOupC0m5cC4SyXaHJtIEj0iPU7Zo1dUswj/O5b0qIWl1ydTWK+TAECn
qJTROwnwPqYFgB7HglOVaXXW722xVAPmstSSLfkQyh5Ky+JlgplIbdyV8ryu4RRjYT2O4BChUOz0
8sdKLvRkE0WPiWUQ1vcnWDn/jvMaQ1DXjIlKv2n0uWC3c2P93Fj6+bnZigPJzG6/LKH3vkKF/631
glXD+YXJzS5nU+xd6a+LSBy+nzODcvSAFqVqMKPx7aYRV/5V6wfJcVHFIOJylSuGXl7UraLZ0I40
8YJuJfD6SEHQrAvY1CvzMlnLlESRjCOLIfWfalC3/60QZCrujQpAi78V2Onl15VpEJqhoamu8Tvk
LBfDbWRXhP32ZLKdNJcipqAkblmt7kSKEHUYmPuVIsm/LZ+XCTv9X25yVInm6tEdUk4UdsVwaGUg
ceQRtZfdxJw1r6K3/Vvy3m9XlIxszVvueS9Ufb270WO8Zh7VZaRaAwzIUAQ1tQD4t27tqknAXUma
ji8CTzPPCNkWamNG4UxmfiJwHTj9XzUCzDUbbhugSBsZkH+ulb2eDBsBG7llRgDSUhQUHxNGt1Qz
huAGpqYmOJuENYvLHJSkljCvuUkwkLxjr1FrKje541IX8XDIy8lsXkgTqK0iJ3zVXuZ85qSUFSZd
YfH5T+Uzu1AYpAhcjdsg27jOsM1pNGGY3932Qm3AdgcEDJPqNbqzWGZkvRaAhtaGz5wboVlMoVem
yyH19Y1bwXTgtisQxSTucpfoYImVUD5EA+wg8STmzbxzrCZHIltgQeJuIZgVikjgjkd04xN+VyEu
pgIpho2yddklgfT18xAYrLSXodviSX2r/ocdOJYxtiKd5SDCT3Q7s9jYYgGxpZh0mAkyO/pgs/w0
7OxE+nNRXtEuNygcohPjkvntmviiWrseEMxa9k7pM5SiOc/b+R9tXIReDxXXvZIyey56K3jYZdjy
ckPEonii7Tdb5GDOBlMKI9Lt8owlaIElhG0Im8HibHtXmV9FN+KJkHQkdlcK4eV7X9Avxyob3XB6
VVk+i4vX+BCMdaP0iVXcJdAKywjoOJZbUWHAz6kqrP+yWCRKfAI9lW7IMA3f5VlqimeVAj6U1f+8
cxeN8kk5m5RIuq/o5PbakeiBRnCoDhXN9JXyXYuJ3abHP3eIxnCVB8IADLc1fDxDtOzlLD7wsBbi
Rc9ktX3lxjkmplt8hcXGpAU7hYvpCqtVzM6MXqr7zpRQAiZpEXIDUw5EONqigY+CgwWYqsiIB24c
M3XcIoZ/0UJ6IFKSPIh9uEZjEocCcmSezvtQtdrrKXvynyvwJE/X6+w7aSE54c7UZvMzS7TlTACN
xcAryji9EOEi5VgbuF6pPrhMdYocatDjLaVaZ3mL4FSlxh/wVyNVF4WylwhpLGvOy3QDiiaIG1id
HIUw2J6hpalLMMMEPiReZwf2b9aXFMyqccMfG8y/bUMEFt0wrLYnhWxR+oBXvt+T2uuAfvqFDdF+
uzmMowAyzhOX0gyNaL+s6fzq+nVJ2ux6BdswS95fx9Lvl/CNrEJKD2J+K15foUeRH3FWtZGn9a4o
edmumljeiYfYSRbiHE1HopNVXvBMgpk2wR2dfPzxiIyYhcyFlcUQQ5CsLrVbSHz1bS4fsWtm0/Pu
lppMmj4b0BHdIkR1+AB0We8kvra1bZoZowsPrmEPUzEyXKJwehPOz5pO55csY/XTJZZQnIZbxRyi
VG1V9TQzbCpHNn56sIQ7bMYWdJ35yIBI/GAs4A4b97+YPOcnMfp2PDuX6JRdMru6Vo6ZFZMXqEEW
3ZAnW88mK9hf28/L9J1zkjV2HriqejdawLWwx3i4mkvBoPjSQQ9eUmVYP1FgHfbq+vQuMtqm4BTt
hX13KuGYGmddcRHWmytb9r9oQFgPlWjZzM1iMaFB1Xzk1PsIzs/AAj9u/NLM+MNNlcoPg4qhHlgS
HMteKUrEHe9V/vy/iJXmPx05telg0WN1JgLBkdhqxmzZsp3WeS/WA4XfAoZNy93JoB2+y1dYQIH8
KoSVhyOCRuZE75pz3xUqRbsR1g+AvpLEjhoyXAQxLg3bAr8YEKEPZAKCr0ir+7PNtF/sRAZnRJDd
4i13Nf/ZNnd+ob8H1D2IQ/NKyabNdWjb/oLORDCZxkXixBbLY8TwJvDUUOcPzszdod27k2/FytGQ
xNdG37jWTVV6gNuC3z2k48xYayVbYhiKF0+eQktMu0I+bwwru9VLQP+z4+xsXyfycShnk3ywnawN
yA0lev/EABmzhokKQAy5np9sdSGiAS9eyiAmK8P9kIQVjbik26V6Vsl9wqBJ9td479nWYQli0HMt
+B96OkEnoMOaYBNeONTVIYKERyHPz2A01k3fPG+QmiZ3BgKOBU2h/6YF534qrcCbvKsBegR2IH8V
dZrz6XZEX+4tEj+LBw8RHwbphNOzVw0VvCrFonU6FPPDd8tWAZ5RdB0ewcT5vDFDE06JvNux9Ywf
ujNiX6EiwKv6UBY4todU34dx7m+WneX1pYXpnx/VBgl1BobBSbfjYwTVDXuLt0P7fVlflsdJAsv4
Kpsl6EJCU551ZheNnwI0JD4adhMelD4VvyQksP1qYKuiCGE6MiL6vzKyRxZeJSNS7IXAQrN1kwxz
FrMCCw6Lujf1hI6k7lhZotS6W9F+D4qdYaL59hL+pxdZV2kwSS/H5+nFWKLG5sHW3A3Mg1XguptB
7x0Gk5ymwe50aToYLGIYS9Zl1iFOYzZZ6J5mpKkcopg2h8scdLGLUs4n1Xfjtl8zUOTNi0lFg3Nj
mZrcr409Gxb2q9SmnGG2X+wFZAy5xfy7Z9yD7zHPTLqN/fND55L8C8195pBOKPZnA34EwOasIL2U
fQ1D1j0p6hehM9xZqTJJ8fOT7rJfCXbmJDYwiL0u+pgl1lYm3Nsifg3mGK9Gws7wYbaQIfjtMd2/
kPtlIc7+GEihr05ZgDWUUzf+JfQT7VcofUdog4jftUf8l0sUxr7XnGkAW9SG+RBVs/t7M8fW+fBm
HAaxopUQmLJzWxIRcHtkHZ4YM0UXHNWja1L4wKuHtEw5esiNTQzwKwmpZDIiH7CekuTOEg48HCK3
vOIJ44J7URI59UyZH4SPunBdT66idOI9adJ9Yl7nS9fzt9+iZlM0S6WaN1drMoXnIghAoFu6+xhe
QMhbV0LywjUKrLPpcDEP8gam9rhXoAILDXGZqgHzyBy0YOLNcYQQbTG1H3MMJT37J3AWhlFQcVE8
EGGBmNCfPLb1aI++avgDGK3pVhDtbXT8EIOEANFKz03FWTFQCYUDSB8Zf9u8rFcncSmhbGC28abW
e8PlLh1wjVxgP1NJBUMIuyob3k5M0tCi2Lal6MZufTAHlKb+7KwJpasfDuDQHDTuzThWkFD9r0G3
Vly7LbWF0ikgNY2FPDiCTS0Pu1eboPT6xQq+2yG2tvBP/OPpDaa+x0w5SMZkBfuQRolaZcKUWV5y
nxjQw0pOMne7yf4Q4fGCcEJOqIUbhPGKyfX5j7c9SVi7z6vrAXV6AuD0pW63TQKu38mCB8OWJ3dD
Gng2L0Wy2U1i7ECGlyeFu4rbcgEJekBV9pgvti+vvxi61ZW0R2fHZwRtOGOV+2QBYU3A1b/GNAQq
RoWxJrYx1yRO5MDkTd/BoOx/rhgn5OEfr+2uyufS7a9RNhUx2JDBWXAyu6Qp9fOAAHYEnUrdD1Qq
vLo9Jm1pneblA5Jisji2/Kzv9t5ik2+EqQza3gBpzHKlimyRUOVszJ5HCn8UoJucak/S6wKDWDWd
N7hAIirMyD695Zc8QUcogHwp5MixhEAsfvpu94D9+M/b6utmUIqe09DGXFIfGMXrZOdYvWFUmjtB
GEONL6MclOvL4oSkXhPr3rxGdoASzlOBFz71XijRwInubs13N/zW3/unrAKUu4Xx9a8m62pWjf/z
dJss2/q/mUa+rQXGBQNSvlljC6MbETk74sFIe7R8ShXyr5hKRNlp038+oQZTMuJLkJk34k3ppmzJ
kttT11n6AqOQSrxBiHLSBefS0V+ZnyETLrzu6EYUXBZC/ZBS0eaKEUKl8RJVaYhTswFD5Jkaxqw9
Vgf/Zo3TgtUl/63NJgGp8OdER90Kx425OxChpZnIg5cUUItSKsBuUNvbBBoUM2g29GQ0E0E3cpJg
ska+br4tCF5s7XWXkxLNn+CGyUgTcR+fC53Oj1R38Uk8mVuLHJPY36bUrDGD4mhZfv8bfiAHmLTI
W3yvHMX9Z0yyzlq9fvwKOr2pRNEMSeE+oYKTHHeb1BVoXCUlwBpPMlY5+u1CxbMKzAykEv4BaH+G
HEzTmmY3tpU1vB0ypcsgPjJs44DB3RoxPiZzqLqD1uqOD7kavWeXn4NjnrxK3dHSJ7FzNjuUaDYV
aNwRa6I7AdhncZCJlR69RH5zVzNoYWvCRbwL/c+K0AO8jWbgZjOEWX+w8uV3ltNS4Fn+ujcrMbTp
NQCWZYaWExDGQzS9TAllp/XcgI0MWsjnUEyVv0SL8weTTiof4LqAdtSfBXPmuYZ/f69M64PTq8bg
px5ad7U7H2tG7lYlNX6tL+3SUv5CUsL9PQim6UnrEQQTTp8mh0C6PvegrW0P93312cKa99O97TjY
AaTJgfJ38iaDoXkEPIKDVsobq8xC/Jz39SrsVG5Foy2H13C40sGuDVpog7cACDdCfSIJ6oR9pjLx
STeLtqgXW1mAAx0IQtpwuPL9MWWZIJ6M0UatRGPH4OkqaabGknRI61kXYm8ffkrqlnd3/jpQN2fT
XRKS1/+oYLXGyja1svhrH+prcsR3ISTouXBOqfUC3SsuWsoz+ne2iDa4br2NAJwIKzZC1S5xA/oQ
o6llEO8HdT3CPE3V3UbFtynjqehyfPY4Lm6MBm8KwZw74IsAc+IOX5pF3th/GovvBcQS5IKaXWEu
ByVEGMmUzZekN3MkdZZjsGwoDrzNN9PgmdLDE9liOJXhKs8hZXlKVxnXfLXLOzk4fGuWRzo3fOxR
GTRe5rmZRyXUFMCMGnxgCbEbrZi9RYusEoItI8i7KtCLg+mkSM/2/u36MN9h2++7Um59BY1JUrup
xqE6PS9nQosCYPjxu+nQ+32oDF9H4ypTldBKDHnIM4qp+ikuXrZ5i1/pWu10NtNsx5puKT1Zjnfa
jE7xZPyzMdinzUiiubZ1v8D/Ch7n4WiLEWf8tFsgzFLVXeLpbTfTpdt9YldgXDHy5BX4LW1eT58h
0UX4IhNa3L3uriHEGwm31VqnX0TFgqGxc0XychVUqSFFpR5L8ppyyOqLZ7NzjLoMdf+ROXCzTmC9
VXq6lNeQ6LB0QA1K+8ICm/qB3EiKgsK1Ng5G62uMogOKJ9l0K3PyDQH+jgM9PTMZN8nCjRcUD1P7
GmbNvhZfJ1XJswwJiJqzAGVahlJDoNFKrdTBdIlnM2hGGBtIYMkIiaDKiJQk6huRfcnpHyDcvL74
2NN2V49GJWCPEC9dMFu8cVtCb/TEntVlVIj7PGIGUpiP7lg4w/05J25D28GcEh2GrgveS+c8f2Zc
t90sr0d5EVhORLSaGWZ1kb2oUDsuSDGMnU+E8Odl9flYHevKZ/dJi3u6PnRKTnjKrV5bl+KW0wly
gQ+JCDVMS8v6kfl7RgsT/h1+VObH/Walwiq+F+PnyOohE5ynvaHl9nDuUBTOoBEfyezXVCK+kauG
wr7V753xXBfT/T13SJFtEP077k+ukIR3/k3COHR15tvfJwTpXo1HlL+bwSV4tup0UQBkCX6Td0nh
ZtweVPWctcEpLu1qBL+rFxZOEk12Z48rMFeCQb0cAoRiIMfO3yCn8pIq1LhNobf5jLh+MlA30C8d
Ts8kQk2ZLkAMVjJWQnG6s02Y8V6GQm9jA6N6eIMtkrIvhJkh7Ng6riq6vgmElY+QyEFnjFCIL63w
UQarBHv+Vyg0rpyFUngIO52qYZbpl37MmQThWRHsyWq/obhnh3asZrEvutDKWT3g6QXVX19aX/7d
fUMrv8CLkLrrduCXpw65rLgt0M9EAvyFEb7rM/aCv5o03XVSxkFaNHsZYbRFMIgpd7tf4NRPLdtt
2rKCb77WeAGjPBuDQR0dXbp5VAwA94ZUoGZlL4cbl0l//PinjUXfkKzJUXGRjJtlLzqxEAqCRnvd
GP4iDl7Xn65PVBrEdP+/Q9WeY+rYcquhNh7CQMkZYLmD8yxVW/F6qeoFjFGgb5QtH2+YkH9ncvR4
kUJPQQXLf6fzR46NueVLq9osuI7AKfp1fimXe8zv8iWX9BeVsinBMXRhZ4l8YTaLTHQvqqr+9+B4
XruubIbHdjv5wSgRV7lqdeNu9xbc0h/0JtsREMRk2cf11q43yAiFwldtNjg+f6QQh4oW2LWROQjy
/Y26ZP17jFL+TIeF9Vjoehz+WyU3CD3PbXd+rFsBpf1zF51st/s/4rBIwoIjVX+HnI8CHwjCtlp0
5BK0gYQZbJAJoaKxISIXKdvBTKb7pveQiKDpfXRjx0Tv0ojYa3eIYudERjwAbchC+YJalqmclGMo
VuagIl0JA9cojgVEZKUuBOWu/zcee7pjHuBVaN75OOLiCLHmIcHHSOVZgsiNXG2PsodzbJ5u9Yyj
bw0EIGN2nZw3/xX8X2CrzHkEHv4J/5YEdb6/o1miJBt9KknH8Gp8NBAj4uNjmlGOOD7xrWVal5x3
zYl6kmy1Knz0fwfDuRpFvuu5AfOfjxoiNdhxsRADh16brDj9iKB4PkS5wqyS5O0OxiV/VE0lpsxi
Cs6O1IYRFrBDP83Y2lSo5eF9WSfnVumyQvFKlk5kXglP7e2w1rjebUpT/T2kd7NniKrxYbX/k+dE
1lO7J4t1z6o0ZJ9OowtGXEHFEC+Q9zHpwLI2KdiCs+AaoeQgMimY7XPjjGnkYHXoAP/s7i0NXHEh
ZobZE+eMM6qaypXlp6vDOuu/mQWrJM2Ar8Gzr3aB6xJ+H2/lZeD6mMHhUzlcrZZrDCWm6iRS8gdx
Ec9LW5iFQ5vDPaaK59H6CqsNaXSKA8k07oRCUKaRXvPwDrkDwLQS23h9Keoyl/Lzf/ZoTOIHTmq6
t7+bAryY+om55gt8ot/7cVxHqen5HGwhQosvt+7IzgeHlEWahEuGIFkRBfr6HqmCGoCHRHSkNtzX
chvnaXQFHjw4SGlHUhJL3BN9ufsGiMQZuUEpc43OFTWhgm+DEfWtPklCh4BZNCwQiCdeq1sYAfjg
5kUv2g3IUcfCoDbawQMtywQVLlGgR8DmNzd2rsbMzURZwPmeSgiaHNkYLxZRtL2mpDP4lLA9ZlnG
DauZGAgskMN5sEDlZMNe/6ShOgw28+aYjyE0vIHfXDcmpWJaVtGxenWeRuJGjB54keN0OEJXfvqi
tPo+WdPhGJs/8Xx8yofiPKlDoPiFvNHESyD4MHkyUoK8X8+p2F/z5c/xvE7vU45v9cXKmVyMZAsp
1fqPiEK/bfL33s5jXI4SzzC1XudyTL/wKqIoAbmrF0e4oFnBi8oscn8GXIBhOHB6EgbflFQ2Zui/
IYBsy4AxWLyKklHWDTvTwT0mFMHKYNzI2BBszNNdjkiVXYorbxPjVJok8SyGRosxpDZmiC7wVA8R
5Z6bpSWhemYvX+FM1VeF2vFjFGYX1xJ8A6yCD5a2uqpTnw7ge3jEF0LBWJ5fOpltvdd7h3lSYwEM
LE2kv3WGx3h26a00z0K3O8ODH5wYbTkAQ5+Zcm5KL0c2uCGeWxoNw0k1DKHGQ7PM0UcKTUDDY4X/
T/nLEY6ls81otfQuenGexHtm9o23DVC5vL79eRWuiO1LFiVxqDR/X0OFnOhJQHDkXts6yVhB/4x8
cBcz2w42vGGK6VjhmFHCrDOoFlYDlSnnXyeemlH4oLWlFWjAAsXPJRdZo6ZZEvZM2EwG38VgbAqk
3K+cUIbtkrGHHP19ZhqMnhn9Qn4hiIwcm55xAwKPC3FJ4E1aH7+3fnz9tWySKUNNcqrHV2T1/LU4
vF058m2RgFk/2nQ0pKyod21p2wTRhOOv7WQ5Jf1OxU2KFvIZdQd4R+RW9KGjozSbnGxLFtYv+55w
/5PSxcrLvBjbgz6apCqaBAtCO7j/DWMpx9Yeu0ctftEhWwYp1Os5EHe+gO23SDlqzXEDq0B4vOFf
oB60Tu2xuojxeaO+lWPDlWAK6gyCKWnqWs2l+QSeNHGoPbZ1agEwap0xI7NDl+dYcdyWYRTacwd3
rOO5BN9YKbAVwS60bMAuPbpCSJ2+X6aOL7MrddhNjhaTWpohokcRf5Fmc2bA9kIu7gYZTc85HXx5
CEgfqjrI1gAd6zLPR644+3qhSddI1esYjSN+YR0KKBGq8kTUWBjcnliMvJGcqAq5i+6POqreO3Uz
8NSiGv9Y3Azeier+GEtOGBgSEB2EgX9bXbLnhu4NhNetolOfMEuxSglTSAB+Bo1+bVevrp2az3Qo
LSPcRkgR7a9SiyppOgnxBwp4rG3j/0fOE0Ehdvuqbw0dSyy9rq0iBIG5HrkdQ9dz1kA301QBIPXV
ijyPvNp+lib+HuFgGH9hU19FOdtQVb7EPAXejNbOxfAdLRoiHv9CGPUJiUcDK4CKc+kH+8skIVEO
G3J6q7sAmO93rNMC40xnpMNGw/wACnn2JBCzRk7To/bvYzPCzbv+Bj+f6tuohQY2NVQVJ2SccjxV
tDprwDN6vMfUL6bGomYiNfE4pvGMhqvBNgkRntl9Wgz3b/4y69NcOhliTeeejkVCIa0B3zfGbRdb
LDmaWswhK9ETiYNYewcfvz/pWMyBiMzYnoZDHwfrkfnxTjQ8PVpRlC8LQsSaq5c3co9S1U/YZ73q
yF0Ba9PApZNZ2ArTS8LRcHj5BD6mQPQHdxvtOyGhgCfHEmVEo1aioT+bWQEK/r3A5yhEPZPFGp71
U0yLXQ5PbXE7NPZFZm/w1np7vUhTUt3T5TFowdjo3YUww1WnJobUK5bwn1iVdE4Mm5ZOtBzyhaCz
qwXGlS5/1XfYBjfbnqmqqRaQ4gAgkqIYiHsfHfu+mAo1PUgO4+HUmNMBPbZq15d9CYYV4C7crDFz
HMfdeITRSBiHiSt2CbnFoQO8bQBZEyJRoXLAQvEpbNJFhOkbqOX/a0hcxhLcDukrNEOP+WKz+hZl
/IYRcSE5Y1PLZCIXDQdUxHhc6zrnGpEA4JgATuDE8h7EU0kdqzH2CIpn0cTJLBn2IS1tN+AhaBE0
VvVQTmEWrrh5Hs+UP2P8jZJy+Ko3r/DyPjhnYi8YjOaxXfwMaEUst7JDlYDzo5T6/ocFnWLSD/1V
on8Rhj/ILZcB3M0y5wqKHHv/5/Wqlk8TBLo1CaRUrbJyip8ejxBsMjbSH0zja0tHAzuNJBpTexoh
WUOOTC/XeJdIYTmxJaMhYb9voF/4mzhPWyau/qiBzRj8UcWfUZs9cIcW0Ahz7K4GzbN3ixa/ir/+
/8d0z8jb3TtBysP6ecqEPzPeG10hQql2+8ZvdzteP5KPU6peMzXF25a+YJj11BP4lOQ4pW/MzRIf
I90pEkv0POAFTBvgCVSZB6I5lpxJxgg0FHWx4j8CtWkD1S0puJzjwZqBXa6GuXR5+yUAFKT/nP2R
10lUPZAVx+k7TUTpJrJRiRTqz4gA7e0QHzge3dSh1trj3gU+uyp1OhqzuFeNV2scQBYtxWNHthLn
KbdAEbxDc+Y0RIVyRNQ8PTTnp/s/62dzBN0bUjMUq6VdqIjTIlIhuEaPPSkBQLwDhZL5mnJojLmV
Vdr5bFHaSfF+bC0/EM7RiKUSSAS9sLtDdz0jtJjTqry5bUIEgSYdhNeyJaSYkKG0cpShx/Jy1iM0
m+ikgTQMnMIFDoSXpkXHajbHbpKcrjvLDYwh5uTv2Cjf27/F7+GUJiOxCl9bbArHmKTE4ff6Mb1U
+oOrG2jgPj8uqrmJqjOY7RfC0Ts3ikFLPJGuWLesZTvQ0OX3AHaoWhyWrab9bbcjDG4BFESt3PXW
QyAspz1J/ekhQ8bXyaVMfvPZpwXLgn5e6SAJzK9bgccprx9p/FMnOvGAA7mgK9sBxYS50BhpMP+E
kcQ/gISHIf/Gky3tT8lpk05exlr2AvwnHGXo7srhnEfMerj90ILpBTwK49QEJufJtYmGnUoFKgXF
Lgz3xaYQmdif9i1kV0k+DCbnzMVV3iSdFHq8yg13H2nNyMvr8Y1Y8lRuVxc1YThwbH1Xz363mlLj
u9jfQhQI4ddGjEVcnHPUOBx+yGQ9L8Ea01TY7eNzXULiGjdVeE1t1IN7/U3kFedplIh9iCOhKRHn
LpE+8Bobj0VFyFglgYI4EpOkIVArJ8BFZcu58EUciQpW7QDdCE0kyBy4bcGDNdH82dKbzBaHhy9T
njeAjk2/Jrau7Dy6YWAMOXxzk6buEUf5ZQ516FU5Jqge2ojj8W4TzXfDDTyiEaRKGoaZTiwOJfsY
USu+Hd3RwHBMzmFPIJg6yGkOi74H3hKrzBpGIs9tg/hjtKvONdoByo6p2ZHwlthV7MKBu80Axp16
qcU3sH9Fs9GZ82pGoSmLP8CEwLynQM8VAwXRYOVyKpYo+3GGoA/JjDjRmlchvEWIcYXVQD4D4+sC
syI0mE8m3y52f4wY9b6I+7ESfeE2bnLBHShtimKr+ktB0ItstNPAVyqEBricSywPiVB7EqEzzfLL
hLwZBwqYh1U0NgKYgUgvNI/VRgGXyHsHAxY5/2sasKMw0FB35tKuwi8VGDiieJMWSM/8ibvqSDZI
WAp+AhERgZADF2gV9lPbcushjcBnny7q/S4Eg05NiXmWuV26wiQjLiA2tUpxXYhk21A5hhBsliS+
5aYZmWBUBQr7NtV7+8MnSZjDgrNCkVw8JSZi0A/i8XNJXAMV2NchRXKqDVWL9WRQtq9agjjyQaYH
Vrh3mwuTJ8r2g7fNj+CWXKOzbmjnWiRoPOFTvrk1DhOdXoO/v5HZ4oIO79dcSHZld7M4va3KGL1j
cr5+IG4Dmgbc+GIhRt0jnAHu7oyg4j2Lo16drCLxz/eECpO7pMfCEzFH7ttKP+IcutyI5o7YKr6u
jbxAdNrNEiqKi7b1pyqngy9myTS//ZjpAkkkunP4GFC6W2Qw8t8JRxWTDOAoA/c40JGp6ikBbUh7
vMeGO0lXOJZ6da6MSr+Qg7gOrxNdfqW63wtPKHfUliVAjQcJjP94OYCXvcz5mJJTpzYha7z/w15u
S7xQtSSZBaFO6/d1G0xv1Inbv7GA9U+kVQAcyfaJ1bhMDYaU9WnS6uyTAk3dJf14c1FZSxFMj6ID
vY6MxVFN6pSax85sVbTM1fS/1hRfsvvC9Gj/gnzoiOrq9MdBgk7ajEGpTQkBncN9BV4hghqjKzLy
/IWLGcrjR7yA7ArV6FbKAmyqte/JEhYu1y23f4EwCZWdGFNoBenMGOHzrzfAJU5lkzQsRaCQaN6A
/gGqAhPFN3SzimReEQllgjJJG9hQrEm0Cqz/bnh5/s9moD7UeEXwk3i+iYC4+d5JqCTuULVJfgzJ
pYloMqSKuc3e4jy3paX4ZT4s67l/qvtBP8TK2dFLfKicFbysBxRKfQRHamIaWnzToZjp8z0sLS/8
Tx9UwmdiVfLN7avodfHUq2ZgRWbPRdlawxCW9GASQiLCSAj76KuzuXgN0Y945rZVkd8KSf33obsr
3cyaDCbGu4RvHPzNeTIjPQAFf61XnbsKaZXYhJxSD4TPW0cIrm/HnNQTBZZyuH1uElNhI5C6+sdp
xJZLmnR4fzBlw0N0npM3EvBzAlVk6U2mxU3xnapNlMGfvzEKVpLSqYSKpHmw1eh1P7al50C1zHxu
75oq+pj6F0gKpZeUMyyHzBTNYtiKwYpWIVDS+0hhvQ59GjBtSI95T7dFZ7/lYzXaWRgqF9odC8Zd
050+vXXjt9a7zO4QveRmEBr8FgdJAyyVVFLJqTRjekWYMcXaB7A1xab0ZV3z5x+n7nAPMZ0iVIA8
VUrvbxK50DQCBxPpqxSd3eBVc2KDvAlowGXatQHoq840eyPeK5IF3SvrXGQCtaTxuJ0H/3ol1jCn
gAIewnP7sV3Ucfsmtkk3v+D+3tFLVJ1Qo7ZGzwchEe7XHb1wR2nx2F9pqaaXiRDanUQ0w7IRC3VB
kMMeEuBi/MppD7fF1PO7L/y6YBYhrQSmb2wF++DOEUfknl2S+k8Oy9szAUmD/uyqcB2OgHVo/ZyJ
rpwxQQncaD69pD4S0z4wWiGUiLm727ihR47YHTDg0BzF6pNdw+ypRA8+5KNi3QFD9Vzux6XoclPt
91hTdbkdfOWM5/H7xz7+fmgEYEcVw/IvPV72p5bHqooLmvUa/2QtIk0e/EpSRb97y94ywI5qwi5L
KApD2x8GsjG+Ga9Ig3D7on4j8Iav75dzqQM5lBtMDJ+m7cIeW/SsOxxVTkP9lIy8BN11zEYADqUF
guy3JhfgbtMH4zo7eWUhW/kVvR7N0T4V2yyOXUzv1A8+718UAMZNm5HuJeD8IPZUM5MrwizLmOle
dVcFCfm95jj6c9LV127lquFEdG+7ttc60+Hm3dgMA7oiG7SR86WPWWp7Tnyg7CLoiSSEyJXWnQ1n
FA/h7VCQHsbYQqcPfsmdyxzQpZya7ybE5aGG2aZSG6jWNvDzNEZRQfA7x9LsdvwgYXbd8E5wpEbd
/QRZ+Ep1Zv79seJW12sGR8vCoyHe0PaXSPF4fSfAtKOW/BNvWhKEE7UaNqB4nNDoLEUTXufWyNo4
6GzfPU++lkrjrE86QH1WiTYDk33o7xznixmy0wgh80ToI5yFbVvfx+EgcAYQmRjdr4SuK2bpXKn5
57QYCWh6jiDzDXrr7W06Kumc8k/0Z7c2c5mYOEWeol+7G5bMmHj/LRAuuQfxtA6FTeIWswt4un0y
SEmVv+0kewLj9hfAR/vIjWPt1hi/xQ8WktQr4sUKUXsWojbNBfMWNPGK6rGhqnOjiRq8ocTFObef
hn73AgQVhZ/+0LQrfMbxXb8g07iaXRfKL9AcS37y9HzkpY7cVwISkoD6rzMY1rMEZCbI5ntabD6c
Gn1rruoWWWYqPfNnfWjHsqRyC6ffak6mrsJj+GSdKqZPLvM+GUFxEgBeDp4TGEJT0s0rcLP8/hQc
k61/Psueh5smZA118YEtEF/3gMNNNSw9YYdTztSXPAqeM8rnHNtLZBi38CIg+v5/3AzLCcphGwdC
WshywTIoHihMVmX4VMvS4G3jmW/J7U6352p0awLMqjGm75n9FGzC+YT4dFtroUxoYPQ+i0HtAvZj
hdCz91RxDjR98lMW4y9zspr41TYcN7sTeqx0WhY9XXMdcSTTxNmmDvc0j5BT1PrndbFHNKpfn0IM
DgGPrkk0jWMDH6rOG5ogTap4zcpZcPE7R6KNhJHAs6KiZ4T3Taped9FJG1qrtDjBAo8D5jvMVsfP
49FEPAh73jCumWkOLgKf6W1baFkDYwDC4dcXvE/rl4Mq8ytykkYD1pXdf6JjP1/T3qVT/7+Rwq0M
AWQOSuCdZ4oHNjkr6ThMacHtcpQJPY7CbHcxasvw0bf05ctYMS8uTlDSdFuyNI60VeSETN/3e/As
0yfnLTyQmbc7aYk43Wb7FZJLAn2yGCiqrBS2xaeIr8iD78gIuyktneGQ8y46b1Pa8hd3dDmlaWAd
6PL4fffXH8M8nTlNCpzNI5MTA3VThMYQolYpSWzU23KcLA3WFwgq0kOmSqZbL+XrZ0RHXiRqOBr0
tKoqi3Ogzi6IZBy02oLX4alNY89BwSt8crVFww4O90Eie6Be+vmXPx4ITV+GrfthgIuqzK+VSJaZ
vnZmpkJ8mujdq2sBHOCKlIoFO/qIHZjes3TgHeM5DQ5f1xAIEhCwkL8U9Uzt3O/eDgOlnmUat8SX
LrP73Z/ykw5NnBTC23zolDU3LSJr1zVQJO107VGWOSlsPqfnaIut1sfDA7mhVtltY795l51chvxE
qYsMpJ8eww/QG8xd+VzRGGQs1mQbYWRH5NvXbLk2xM24H8gxUOR7kulIFfogdKxOZKkezgkVZZ5e
zeOUSTolGIE37iMswL0sUYu1X6O0iGo3d8BpCWrey+t3Z7ONRL33O2epHTui0U50xRcXQ8FbV1xG
4fqTxOfki30l388WARkYMXttXCygbMmx/VHKHwSiqx5QFZ9HPB76xlzFxgWZu88FnXexpwc6AWTu
83O7VT7M1KOLLQJBZPibHgi2fHze3zo7zZlCYS70lC/9TngkG+p8fr+35EsmTZfLQvsihOTcBEBr
+HPO8HGrWc6tTxxvzbYQKl8sKG4Db0JImxRsEH+1e94/91AgWqXDgm/B3jDpheTBwa6AEMrGu2Pl
Ju73xOr331GdvK0EVIlSLJsG8GfZb1jFwdrlTt/wV1fLlFmv4Ihu/rkiKLpmlXMHyk0uvzVafg+b
X+GcDUkcSyOJEI83ZXvkCzqQwWVP7bC1zg4xWTQI/yFwx1rouZm7dM6PiBDUMUWktZ52rIKZnbXu
HWyrWG5tRE6mOJmKqKWkTYynSUXb1wGgMlPyoQH8K4jHydFo7UYLIfx5iKnBbxG8wGoZarXkw8bw
2eBFJEjjA/yccrCjCnUWAyfsQgSvVlFdYjb6OoQD0peKvMZhalEM25zzLdwC3exmkNwIqlw2Pmff
bLXHKy+7U50GtYc+IO0vXtShIUwtoPFhSVpIzFNiCalpw6jdKL7tCr78UYJKoZeMk5fiRp/eBh4W
kNwa8xYZEesmiVN5yRplrW/Y2pc1gwmp9VQV9gAPdQvPq5i3KyDthNqSZmG2uuGQwnHVR9vJtFtE
PNcf0EzgMirYw5QN4BWWQY7T+92K6z/qMJiSyyP9Qlh3jyszj0zGRKOH22y1EhGNXSmJnaO2EZUq
fQKbg6HyOgOsikGVM/jrhdnKD+L26ypum/S58xUhlat2clyV2Nf5WEHPru9PIseNZP3/FUw7yg/5
vK5/hzJGVaIEotgLCQOpY/vluOyznGSUCPj32PCm2LETqQvNXpyuQ5AhXeIHJ4sIQLurpU+OwDYl
u2KrBLDp4uEaD+aYzrcAHKDlvhd7Nd5Mn6lGlGZcvaRWouOPo3N++MSX1eegx4kSi6qCRKvrB1E/
jlVjGmxHrlqzfIgkpxuzvCB2SFuFFGb8N+KNdjK46qhIhL38qcwf8lASz8lq4wxsrKkgpphFXOL+
Yxj54RnAaslhMPuBcqA3Is2005+tcNE1hi4kE8ig1t5f+Jqw1kYHLdZsI6PC1aOx7IadJUCKr5pI
8xQLpA9lLKjZCk7z80kFXsyvnbD40crPmGH+nn1ZnM38TorrEOMirwHkCdC7SMuM148d5jTIWMxM
WZtKYJcwolQEuOwkeooAvHqEY0POrFSa8DvsXZw1JoupaoaE/FfN3UGSZsWvyIuE/AdB5N6OCNYL
AaoRlbxSgJt5zCsEof55WdNZqZY5gyfLcNZeQbP5cgDvcJkkgVDbyPoCbsCTgFlvaEBJwETSP6B0
lWYC7m0GZVM3+TWnkUFre8c2m91O6hKk3zAOhXrY4s8FkF9vFUBDiBNAkxmAdD/Q7Cy1hdIKsVrS
CN+ocRFtu49lJ1Ww5DpjK8zh3MItlEhJUUwQALVhFtXr7+I5D/pFJF9C2+wi+h4I1x2tnmBgxT1T
f+oX2HVZUSG4KZx6JbnosJYAgyb+x+fOGmTRh3GJjPuf6rqCqTIZYvUdsBvcqJpZtLcP2IqJSnot
52SPdBMpyhiaBouXx2C62e0uGuQartRbb9iIF6Q0dEKM2SYe7P9am3+OqUMRuUR1bfjtDh/4qqwu
30vJ0zAIWqMyyEiJqWAxV803gCjMge28yW6Ysn3BEfSi7H4sIGXbd+Jy4/L3VTZXEuMjy4DP6wxi
BS2x/DIW1hzsszrV44T51R8fS00UwF1c4xwjQExMLARbp3p+3j8G4G/gI4xbWE/2fJUsF9YAR4WP
NIJ9SvBvzjranm/ldg8MtyqGcvDz2HZwd1fSiHXJ9kDzpHutFiWcokEXU8cpNAOj7AWIpqwMV3go
CZBPlcaafIGEBu0wM+03Eu/18nuTtIFqiJvBBOnyH1AH3AaUusY4SwUF3gQf2yXYS1diIhuFdZI4
ywB9KmFLl2CpR6MEJpA2d+hk3UNlNqP+xquF6u7HwVVfnbqjOSSFmZtbppLznaApgfxkat0/zu95
viwzuuYfXoro1tIorRpFziAz1EFI3SMZPirfhXqvxtWFbxc8U3Esqg4YRr3eB+apjuPUDGID9p51
BTB7iuQNwxtI6LsNAMOIppzeWCMVb+K+J4wMHqUU87uqPNhs7+XeRKlsq4hKWb/mFtYFDIBpvs9o
qx+K+/RH0o8XnaeqLJOScxtm1JKIFuE0zO81DVTr7ZpoScdItKNjpQFyx6UWbJaiGNXG5H1NytW7
XZdnM+ftTqFl/cF8H4swsNSdL6/HwWpTOLIkz89wuEIm2ip5YJmvm8Ir8cxhe/mko2LIUWzF9tRA
57dqSWpXr64GlqutI7WMcPNe3d3dYmG9W67sqtp+8puMCnsqllY7qT32Lpg4RH5sebUW0x8qz4yk
5BWOhMFrZzs4udLvT5vIHbmCi7FAv16M2XEOJKd4RPvUtwmGd1pZpL7BuYWRZE4uZU2u1js47och
W4kx3bIRDTzTvdArxForhBRhznnsLnv5Knp/UUFiVNyqKeDvdcjSYVtHq3u1w09Y3dq4udooQHqT
Ze9Z4X9xeyflqM/Gt+R6EC299QK6CPmqhXbtXoQye9U7KyKB5w9VfJMlWNF4qeDfx+/gmzXOcLUB
M01mKCdnQtnPgtbi5SeBILGqSs++GVN1aT4n89pv0HbsG6S2WhSJZ2iBrgDx1c4y3X5QYDM52tyz
o5DvbuOIQTYfm+HQq3CqXFaKlxVJYTZjaR/ReQDviErFZ1rTGG9hmiFCK3isymzBypDyzm94W2pT
cU1LCEQyw1B+x7z7lcy+Ia4MqhmbmE29PO9VbvHIoDnj647bnbngGYDG21x3SGfa/i8ByYtqduX3
mgEMPQ+qdmehrn0+rwf6XcjwQ80msXN833p41dUeW8BL6o6X0i1IoVJTKYmO09GbiIYNTd07sXDJ
4MxykstZG+58Bfuo2Ax/4jzGi5kfxzhTUwcI5WnkQwZ8z7rhvZsURY5eXu1Ea6E2GfvG9+NjcrQ3
knzbuPmh8yX7/TbC6ic4P36WUHYxS0I1OYCDRT0PVrT+NI+g8xzmGsOgk8ud7E2SPSkHpv3hiXYQ
N4IYwVTAwQWcWASHwcR+x1mfyZLSXDGO5j7+CSE+K1B4RYaQPZn+teKKRrsy9nAzWm6Lc3XDM+r/
3IDlSilXgmmQCVAXNiAc+nwhVvBHesUsFWX1Oh2PHbwbIebi7k25eU3UzshLhyGfJNuJ9XgGuv1/
5NJUhZSn/AR3tHDyz8NurcjOUB/lGsPYLyQ7bzdC5vjm19rssc04DYADnQLqfF3kjjaA7yC+GqYx
tXnHZT0i8yrFtVieIePzQKR8GU+eN+cSqTjai7YTN5DTvcwtgvfLVOwLJLSHEksnkzSgsfpO3few
2Pkg3Wz6XQQi/aCfbG4YIoMz6EJDAXX/8BXrio72IKgvR15usB3/nwXJd7Wnl36SOQ4bMoXJV3Ot
WYYFLjUkWmVOrff6yhFn+sMUAj9W+5E46xy9KAULRBSxTOjG7mQqSsW8HOD+ii3dMwpRhEuRZ9yX
nTCZrBxhrLjz8ubMp/fz1gq8b+D1PEX6tdNPWtpOVNgPqt8lPr9Ad4oTOMIKCuGazZWsnp4NwO2Q
pc8FUGYl4fyexLKDe7ZedkswchVEZcANOmlAwbNGUW5Gd6Ype9t5FkHkE2WZyqNc2pthX4If8eRR
fTXb8LxnBIkvn8191povjq8/WIMGs9BDsV74PgFHjNwsKbZbDZB1FujSr7xQjtfB7HwCc6fWO2Xb
O45CU/1VWysqdpIStSD3dvkID9u3Cvyb7DR58szAd655L1YBU5JHO+6POU/clBGCyPxV+p4b8YNE
WWavF6zIKi9wEkVgyk5MCgS2T8sI37icYLw/qyo+rcDb8jQyvZdQfTJjWM96PcRyO5UbO4xXkAR5
kTBwrHN8NwjZ8z+WiTCgOCDfOvG/3fAQYdUzaHQnJn8+EHMJhtutrRkLswdNKOMDyywJglBHsuVF
VZWGVOFnXMeGrGUFUqQ4P1lJ3UNoIPS9apNuZv0ADwTIpvnMxBrJ2SbyAPNUhjscmNaB/LC3qd4Z
omoox/NkWz785yn8mzCJVc/irWK1yIkyy80rxu3EVGXFTiqY1gzF74BIGPmprZEOf/rv2SnYUS33
Zse6ngdyR41Fjwa8S6Lt5ewNsSOZwG9lNLyhE88//uP4tOAgtqCtKthCjdemC/4cIz4mGNtZ8V+W
J0ZEeBRJNFlx9JrrHJ9SRzV/GW/Ysn427fkBDyi66ZHu31mK7Vbi4EhLV+ZYzLZw/5/J7m3jVrMn
EPYn3NqfWPxkvx0PNk+7+l/RJyoAzhAn0z7uqWpxYsS1ZXRPFhhGzJN75W2JJR6dL7n6ScxNQ0cY
oZPkuYJ1SvVmG+nUNcASxGPHxfptnvwokQMaeS7QPZH3qdAjBFh3nNn/OpxIL7boK8fa6KM6x4Ra
+oZEy4z2yhmVrfMYmyU2wgeYSfsju6rG+nyDrjeKW06vDYAHP/474IFSuPbrfn+h7gFoH5bjgmTT
e1kvs1Bxk5jAhNERj76xN3XXKT5pmnw3+qUXU9VkOCCjt367efS5Mt39HmEwb4byK8TWFiakbxdY
qz8wnd0+3Qtd7vP8iK/UKdfyCE1fFI5b4EgqE65N8dfV4lqci/FIFp3PLpsZSnhnElkAk+iJG8Xs
ksj1OZhWycEBeHx9YBCywtndNNWa6enEPiKqcNbTXnC7hrB556oEjVw7nWEkiFWlEFDczdPJxtUJ
6mAp2BDn3MT0M1qEl9LiTtK7wr8RiH7UO5cj8QgIrtcmmGx6hAmW7k+QE1ZTW6icTnT3PCwb6X2B
Ck0bQyNqaVId6i5B6splHYcqX0Yyj9h6Qp6DKjFxl9C3mxnCy62z5+7OmaZMlgA+fy2Y9uTxa4ZY
26LRl4amnDdp5D7CpZvJOXN8AB+gWtYdMvdkeKOCqwVxUOBweRPNOduTCjB9z2rrS5LBSvCGknKs
qqcG6kbh3VYpNb0E3gICnS/v7dDzrOzey19Hhps2HLzIrxvKPjWKYjfzBYn5UKYYlG2Bcxr+MaoV
tywXwpSoT4arIxilKdL24sxSOen02vVd1KCmlldJ2sO3I0lKGcvMDDVtm99FHHozwlo3ecO9QB37
p7d6LIHsE2AvlVuZbEc+Xv3Tm/5ASd8w5rDt30BNViV/XP2OLs1aZCdl6WiVCGyEFuZ39OppK4JM
C3scuT7vGseSpDCQ/FPYjyw6frGuTkScw/DKmnNs0G4UpSdFo95v8FqZGQCTNz8qFpupKIQYPGWW
gt7DEjP/RBU5tIzUgiP1lr13bNh6ko/1Q2uF3xtgNdV6RX87VPdn0Esbhkim+0zB9PJlGv9izZxv
v1JxS9XMzjCRpkoNnkHYH77r6BzuvqjgJrmDtlOJSP4AtfVKfupuuZGy/snfK8+vAJTEnDY05wL1
6d0nhbEuGsqil1T1TLOwwQqFH0NQa2p2ZaFI6JTymO3VOwibsZtYCMkXsNekHF5PT8yFsFEKS6XD
+K8+ypa9h5VwLdRAEck6h7bAk3q3BRmD2KMC+hXSNOL/Yf2RbOWsHxYuQsiqGIxdeoc11sBaZhXq
32arBbff0rot2HNnxUMGZ6pOiJa0A7HYuLSterTklWy2YLnrZs7hh3SJQBSunaTNW5gsz5c0V+gG
go0nGUdv0HfLNOTv/f81Bxn4lix1deNzwCWYqgqZaVJkr5BYQE0OhrWEXsowCad1eeTNRcbK9daa
BPDvVY39wKNx4tb8meh/QTmCOdOe15KznmkaXZlwgHBfZEGmBYiHcN1pPhh5DlbZE4Opzi8Q7t/T
IDKP1ih/pyBJRB9GRsX1UQ8CoQey/eNge6bdmM2Kannj5w9mJLG2/uVao1nPn130pU1JUSuAvHp2
ZhZexUP9Sq/T9cnNszHM4zhpVBxsSZb7vqmXqKKofbR2nkDMD4zxVY19IqEMCJWEM57FvJksAwD2
4Ot3NVGBjKKlCP3t+NqOrC8VpvsIseFQ6rRv9RErAj/MpkxqRORQuQtrJ2U/rxqXmTQOCAGqInJn
4r/ysgKee4OGAz4ki5SxSPN6o453Xxxn+/E0W2bcX66fYd2X+WEdQ0U4WKgfRRcfWct46Yn0qghf
3zGRnae5hgudP2mMx6AeTx/kE0LXp3mSmgZPM1dlNc9fRUdgt9ufygPXYmQ2jWsjpMiuNAnhOm0t
b+sTb1VvQL4LJWhdwxqBtRXRwa4bytY2sz9CI7Yiy4vPgqR3Q+p2yYCKq1p+O57OQXIV1z24OIiS
8DLcakVy8u31ABlkIyoOalZL/0pz7pHHkg9Rh0tggiBX/fnHd3mfCC5zo8YzM2sHeTDXaddoFhZF
pw6Co/uU5ZwZzWmUf3QdZHkJs11/4SjN/NFfyIqqZoZdG4SaXrcV+7bpYq8ZH/YfFV9yE6ivMNgI
xUHdBlW4zoRr88L5qd40RrLK7zxO4XT99W9yNh+ktDWhHGL+kiKQWro6h5mlq7Ptv4Ume1L4M34z
1tuJDQInlTWnGoqIc51RtQDhShv6VnWI78+WuhmdOFT6TKv6vJ5SovQHzfKXKFZyn1pToq4wB/ng
p51+UyIMbIxy4SPve70GCPf64OLo6E3qAXB5FanlXW7ejGAZPZrS7AEnMKDs6QKzCgiJz5EJ8jql
jytRIZ+nWPBH1pmtW0qSMADxFlfFXw7bFQibOTSMBn9a1IA8FcgoRd88OVJpUd7MUzfhoq0fQNEE
vBU8fSUO8Bm+b7Doyzh/XgLQXFzN1fctFIvMbja2S/TwVl2wQ2piXHmuJIkXT3JGR72cXspaLG6Z
1GKHFY54wtUWsRuePCGDC39blUhVswjBKd0tUNIoFZD4RffB2LqK2WidozHaz/5DYz87f4gIBKfe
bBfTZp9rEnTR/RDZI3Oe8Z35l52DF6IKrj67wXe+ZIFtwQLB2iRdagBM0WD7TJSgeGuJ1NsdAN5C
qGOEKriDLEkWkJgw7hR0QuQFntgTSSt9t6R/LxSoHdQoeVaB8tvkcsvWLUwVSaWC8lyMXXcFk5lQ
DaCfJkCqQmBDiYhbVpwNcEkJS/Lworu8FqQL+syqQkaTi4ecYydz5E0n+++TYT55FYU5Tkznsl6p
/F5x/H0RSyvwFLwFvu17eOzoUKLAA1W8NAYZ+GeysyS7rZ9hpraj9yfclSwbn52nwntDZuwMhyNb
sJPZa3UIKzFlBhEuQgK5XWtIR/txz4uSngTlHkgViEBOtYB+05VCyQ4Sc1vKoi1Sae1hs7hWHrA/
ZBK/86Ibg21bYrzunfJ8a3INLZI4DKRG5yuDK9+5Uhq1pZReKRAvxD4rCj86HdYI4tn5yrsSlrUp
H83RHFvP5CZ4MW/3cII5P6HlglXeJMhXv3l+ZpyfmDnbpRv0xV3arv0vaf+tO23ugTG7EL4oxgQe
srkXCmStcSpdZNJrlyN5eYA045uIIoMu0VcQpZnXie00iHNfMCgyzOszl6d2HCp68OrcNvnn12TI
kRo2zIGWYAUkQdiAO885PHWyTVOdVzynNhwYTLina5VUKSexMZnqhSCRg+T56OTqh1E8sGnbyOqc
XbA3CN/7mw6QPjumsOivH4cv3AKRnLODgXukrsW9iLquY7F5EZHattdCBH4C5kTLljK0KFnnfeRf
nsPSzHvYIs22jIKXImXa41qjPrV5caRDRJjuQoMxaXvuPi+gT/p4aw6HVb9TaEX8jBhiflKNn44v
LiTm413Ho58wyCRziPdlWLSS0lFHUqSI3KK3o8/447nkGOyzfGuORFO9I6HMb7oOMPivGwyy2/NV
KBhSHn+skotQhUxXv+477/x+rjNhdDc0dqylxgmg2x9U+cuacegU3T5zqedFkTgeGiipn80QPD3E
ReheHn2UpIrIRTgZBlfhAzmqRpIgJeqFelyBCY8HeGcRZl2d2/PIOnjiB89JPmE0Q4qmuO19bPkR
RTufvVcSAuIvXUe4tMQ3sOtUbZiWdMD4jvG1iKw/htaBSpwDCjI/vyMx4U2yWbu3I4J7siA74Ukq
TH+QsIQu6Tj0xRiYfQrl40yWHclXEentIZ0GpAxnlYsXB/dFbVZN5rbW2DhKbSAldav/yEUw9GY7
kD8+RAeKdOyeRfOu1JxF1EI584LpR1EMXR1U+SLReXvPoNr185s6fz7pJpcBEwD3ymTHcRwpBYD2
eBbAqYHoihXqjYXMGPbPB6pavljagQF62hn8R1vIESN4d5zHFtgET4IVIWysubYXgZNJuRUeteTm
r0I2GjmixdOcgcPD45rXJ3grzPwYAOwCUS1tm050FRFaYPElkDF8TKvo56yvbbk7gApwIdC0TBLI
WZB+ZF3VWlejdUhsictOOC1FN3zdfHxc6GnuUZ82Az8hFX+UU3yD4gzEjmmfkUAtNSgFqQMUcZO7
Z8vtNGV3GpAx8N+VTjBmA+Ib/6CvnKegZH3xMoF6eWEguOZE7wyLyqrRLT2YrvblPnErasb1bemY
fdEYqXs5uihM9ZP+WCcXPvnzBDU7/NNOgegiqDAOMGCD7alM1BR0oHbFRjmu1pX9BsPdxK1KqtGB
+PPqbL+g5SCGiDS6Lg5Q1ykqN37MqZ6OaKOI6vYvsKhGylQoO1WKjpQ6smFAPdBCxakqHpgXb2X7
sg57sRiAPGsZg2PjMDkSn/Lgt2bFt2Zdg6wuG289F2r4SqMOrdc4ajGWdOdBf0EzqNQ50tqYXfbz
MeVEfkzpN8cQrRVR93rfEuW9x/sEgnvX5m4IIGtnF0R/UtrXsBwetCctkZeDXA7e2Ckvlrr/UMD4
HkbFIcRkHNunOfnPE0zgbS2/lZssWYeHdQ7eZRW5F8i0PnA2KO1IK2FfwSdHfK9JldlMLWVizGji
hkZLBvbWMPi0YtK1y0PLPd2Z1be5eCh50DeJ7A7B7ycJgoTP4iZSeRP/5WafNtGpEFZmIUvvM/OG
iRO5SyFLSbGOMMA/LIRxb6DY+2qJORxBT/11TNjAgeO02aGx8USiT/ngPldfnNYz/J9O3zop6YT6
b8ghs1G7EOQ5etHfcT45jpT8XaIEjhXj+DMk+DyV8NVB8/rMvI9wucTmFqGCDZZtxI0n6ENqafaT
riUI7KJUZAl68oz1h2R7cz8Ccr3IhkbsSzuthJshnBUWNWXlV4ZEgIzzCwlaJijzO5aSFl5xTas1
Sod0ZujEd2YFnbLZFs3O7SrKIVkIJ+oi1bSOCoF9/KSf1c/gR1UlO4zqhPs3cYqBnUuype5cOcw/
3TPfqVIbSOIzs/qgZHHtfe9QHniytn6LcHDgrD3T99aHj1iHafzlM2Tv9yfA4gM31JvZGySOx/ik
f+h2LsOTpd4X22F9LA6G2nMp/iFA5x1rMjHhqyhpLeyxO/11kRplx/FIcdH6YoKviJ1I4ehFyQZr
opLioMbqcqxngE5fpECqd8frbpKc5tp5i0kYwPJerafBbFFzaPki/C3H4CpSpURpllNNRS6Tx2/g
tukQDZzyoh86ofOJPx//11zEnC9VetdJxWz9SWSv3LdY9cgg8feRgNQkMfqK3QAdVxefZlrxeaZg
o1yBXFn//F5yp5O8gmze5SXqJqjPIY400Inr5a1cvfpjohutFUT+qjxE4xQDmBOhV983zm2WL0WM
sIvvVlsTQnE8AKNoc9TL2C5aa/g2KiLAAlxHEdHRd1U1bMJFY6puLEnFa08NOcwUSg2M3Z9erwQD
d/fHuQAC3/ASQ2FdxOqMC/iLOxnLyPFDWz5GWgozMS22NDmijrypSG/iEje6wdt3Jnbb88sgM8Ln
HbTeMifA97SDj4RyZ5z9845skGaMAbSELGDtNlfw79yx9Spt3fQgIxlQDSv0/WvvoLA/HEsFgeiM
rGsmfdsxNTyuX4XWucKpxDfyTRJbrJYz//0+QHjUyhubr6zsH3cqXkBjY7/gCL3O1dQGsKyvGTWK
7MdRHFuCh4qgiLRrLK75z2qjvYrVwQftWKZHaydt97v2nVhuI/OM1ydAX8MdJj+YVsP24VTh4UO7
/zHu6twyFo0T+ioNZSQODk4vwvsz/9eizuRUpfSPYKzENRizYO+UHcqvTDdnx8JM8JxtahcajT4n
fRrvW22JFn+UiuV0tSoHkPc97iZZkyn/kX6BJ7lU663mbBwks1fh6mHclBrRguYXH8u+nVG/wyGQ
BFoi418EB9zJrtHmuZCtBdiKF04WF3I7xWS8VeYGWBKEkpM65ca6T47vJEcz9Qu684r84IiVtPAG
foMq7n2a7WQRzP+Kq4Uc5glmB9u2vbEMS9MtXSuQMoRVE0QzXbXU+zKpbt94dl0n/h5kIRCyBBBO
toww64VYXSR8Pt0MOi7vhGuJFBeT4Tw5bwajRumt2ry57srgeBClyIxkoFRrMbQwngLkCDNs7KdL
0RZ8p9ha1wJBLkKhC/dcZhMXHdzafIfdCLqSv9nLy7s7Yov3twQm7wqGZH0VvILwzdlZY+HbcGdb
vjnd/9i/rEh0sUTzmC61tOXufh+3M9V013LXDuJIt/jOqP3NbC1WoOKEU1vCZ35OjCg0Gc80HWOR
6Vrx6Yn6GDqTWvUoG1e8+QZ+TI7P529PQyWueTovgtdEbrpvDgxY352cUTjhXxmF4F9183o12lUq
LykIHEIR17Qzsx/Q3SkYwjSOwgRMZ7wQnd1KHDBlxlHVmf6MwIVMRcf40SqImGPHfIPU8QBWnP30
Y7QBKOddHSs++XeoyapHGTE/qGhkJDrRYDjvP6hq55aTOSgqRES4qx7m9ip/nbcckQLDh72xIpU3
raURffKXvZfBSkRps7Ehy766MZB6h+e/YolU/ra0g3aWuz0NGUTgRHkQ9aOIGexLWRvE4TJDBBlk
HSGcAsujJpwsuqMj3aiKxM9K47lrLzb1ywrgugG1Uv9GtEHLF50c/aF1jz4vypz5wYxamrGmf5wj
8gwQDWiA2VjcuhL9moTJ4cT9f1lMkwSCW6GbOjNNc0rqV2TJtapVfJ6QCEcDyNrlrmDZ5q0MJnVA
wn7tEQbreWERaAkJXEv7KConq5xnhADPN96ef5ApxZG5IiFj1OKKmt2Sd05kr17Q0OwpnaSRPGk7
A6cZdjkMQvdtlnJrhzFQ4st640tYeXeIS9s14esF8P2+j8yrbsF9pwvSNjYK6zxVMqQq46wbxt9g
i5SoBc9liDNiW9SEbcNRLkD7Pi04C7+5F6Q/ztT0TKbhYN5wTvCQFc/ZsvLbZqEUWw6gRyOxFYcK
3xeyYbz1Pu6Bv5/7Sc1jpDsvC9hccM8eMT9NcL3lZfOd2K2Hufif071470XzL60lwU+nHERkUckk
B0kaYIPlv6fLdQ7U9HbaZ0gQlQWhJ399jD/5ClbaBEPSCxLdBfhvb1j5w+X1mF3hwjpl6hGKIkEi
c5omjPOGC3NkQadRLUNC9qmdVy8OSHiYcgMETM2qSFr2b38k/Zuf9jS6h3fnLORlVHlU9+9f0rgJ
pdb/8Z9viqkhqHwvKq7FEGuRYiz2JQ0J8Gh1RNPeVsNq6aOV0f7VEKLEHapevLfj1T8GkkasOciq
FEMP77GmvRz20Fi6iLWve5kL+JVa3OuZ98kglETEXWAz4gMVRIPrEWJ6hwGLRnd1uktDpPsIb78m
DpUZb8YwtSoZIZuvzAQ5rM1ITyoUIjHor8vqq5SUy27VeBHKnbmoT2YcIgM+Y8sRrMEBoFOlF0jH
SqJXV28v/0snlD8X6KcvhbfKxWuPRQrlYgQPHH1+BZfvnxZZAMSOq/wpQR2dqQbCXJgSSK1M0YRe
7Yrd//PW00fB6KrxpJjC79Qh0yT6gF9nulKmFJOLF8AJpaSknLpzzHPvVenzzSgd9WqaNnriv8as
jQJ5H3RsCTa0bYe3meQeTDx7kDiNSBbVzrKevOFeF9w98rvkEQxknbGVgQuOa4itlBuevgzfix/9
Cfrx3hCB+Q+zAwAorAsIq6rpmxVgqc6tJsD2ebFSIejOWYnNn7jL/OG4DOzIGiwLaXiRVCXHFtE5
TJP6QP8i+fU4R25fgk42nITo9YZVPUi2Qo38JJWEaUvvYLRZtc/8HI0y4OuwiNDHAINopEyX52AR
l1w8HR4tuh8w+zONg5xnXnQQ23ZVGCQFB4ceVOxm59qy6Hxtoro1NQvKNfA/UqZT8Uki3VWyXMgw
tdu48piTuYOT2PwG9XXWy52hXjwQv4pGcEPMIbQ+REAOLmbHxlYujTzVdch1U7zH+QKBbvZufXVY
JfU9Qx8vrd4muXk2Ioxs45T9bAeEtMS08fuN2tXuKdaolRrW7r5aV+BohGk6XN7Q3xh5oEX9utZ+
hPiEFWdN6omvUqy92JUS6hrtWejsgVbsq2YrseVD4aFq4NdPBsGqatrysDdAL0QVohOQkFvWAD4b
+GDen9/BV9CzR4dMm6mKoLuJGRpO3kauj5i/aBLdhnC9YRG4JcarwKiG4M3fFj/Wp2kI9G2i9t/5
CsYet+BGrnew7gruo3iuOFmPBxCvR+zJ0R4Ollzv0UMZ67IAILaaLPp7DaKsc8fkJo03yYe6fkGg
tQQHS/QAxIu55RtvaBrFkhN3DBYYvsB7Y/PfKTS6fKmT0xFkdu+hn9BE8blcqMqiw2wtMpRDBti+
tu2FrHBzzppIqkrCcPoC9ctHmAst7wGtHFEkszUw/QFaPGIWyA/zcMT69DaAnoz9hIILhLEme2E6
uSerUUHx1DJ5OfARplQdOqlSYQmsqq49bMD4OjpnzfITb38X9zlwml593FF4qcGmyi1Mwwh0XaxM
rvasEr6M5L6W50sBzOHm1RFfiEkqUdFCpZPcPrxZv2Id90XQ4z6y+R3XuM2oN3pD68tVqhLIQQzJ
mxtiryadubOmhXELdWPU6GDszf9Xg4gfbVcP1d9RXs66Ru42gVCBLlnOJ+TiEx2oU9MZOD+ZpvJF
LSDoVuEBSidWCO5BHtNb1hlQGlKFGM1jkYT7DV17WVIYyTv0xJVHCnDklj6RzVfQIzgshwoXRdWT
42XzYRuDOQ7qrT84JzD0KFf1YwxcS47kN3V/NqFBNvXQf3rAP6Lu2v5keJ1IHhEwZuClTCSxTKvo
5YRwihPd/7hWyHgKRYvF0mDw5Go5o8ywFgIq2fm2XfZjz5+HEuzGjFxxF2y3S5B6SZU3duEluOvz
5ycyH0HPvy7mntw7HzmAYc5jIIvT8vg3RnRBgOlgrbQka7xjVjcRkg5suSw5W8DGba7FRA40be7Q
OtYAecGGJd2xLC/HWsPylcOt04Gh/ugxnZSgUs+VD8/XuqGQgAkMPptKe/5bt65mrlv8c27Q/crQ
+54UDkt21WBjJRhqgPjzN9l6a3eIr4k45oDQjtU/Dwa1hfP30NdWZ8APRGSE5zxJmuxg/vuHWE1P
KDzyiylP5M1MQRAO63fxYaY8nhpex0elms3vzbTv7UQscsZ3el79NW9NobO0fZikT9J4ccl/XJOs
Pyl8Z4B6sYCh5RIV4AnwoxxRnW2EAixnE9hxMDLim46gkVHrBeldITpNNWacbdPMIEumOlUYmlF/
gaSiKVhv7/NyCj7PJH9fGwP0koBbSnZlsoeOnt55RsjgliAFUjYNjm9crc0/eVCApAkd7PtXJorB
ZcOFocQWkaVqObZXp8OXGdw3dc61TdeMEYE6yxItnvFYM6b66Yd1DxrUxj7AbOS3kZvV+cdx8Z7v
+mmmJw6cbzoD2Uo6977kZQZScjOjB0pwZ35gb13bD1oQIIyy31tszofgEm31YbVCIWA+Al5kHtGg
jtNskHbPWwQhcw7OK80bK9rszabQLmG2YYD2de6Ux/TKlgBZBcZmpPkkzXiDcUu2BN7g6z2QTXRe
Z4z4ovYWMsUIPoZvCqZUcfBE1NyguNrGHpertmfQIynvorWl4VcapKcjcAaUBP3UcxFCTI3Ke9u5
jC+2c6Yrt1T7bpmMVAEgCYJ7taMooAq5AP3Mve+ziSEvRM/8yFGLyFU60mLZ75vw3furHh7LBbvm
tZQrwQpMDERPTVwpmWRkxwKGTQv93JoeDhvkdDWngm4SS3oxm+jKjgB8waPoYyM0wfR9yc6ki9BS
HboRQiwSNg1xzdqecaDVNyna3RrR1/u/1/5gy7xM+PSgC308+hhpOWUwoufeNpADhMrjzeetXr8q
+iOa7nScJcAV2/CsDPXMTVesjZjjmeRzGvVOVc6KPOq6Wi85bHBBB+XG1GCxHZmEZx5unDXKYqWw
xouTgxihM4VZWet75jqLxF+lypn60CruP+pEbQ+6UXzcf2/ezT1ujVRhsem9oXFGR429wYCJITNX
ySvfuxhyy0CKRP8CETa90ojmXb5LD18fV5svpqk9lSC6MedjTx7MDG8vJtfdfih+jO8h9961N99Q
VplO5kyX/0ukYjGaTiqn15SPnoP9GXk9GE2lniPvhqp66whZieVWj6UNBTfFUlNM7FN5jVJyx7NU
yQ5a6AZbwlvNRLQRRE5/zYEmYmpO1idMCVXc/dHUSUiVRNYLh02xoycSdmDAmdfTP3pdjhES/UT/
jdKYNGAS7c29h6b8AEc94iQ9sHn/3fM6W1FoEqTE5lVFlcW/uEduFIH6/C1HHdZV4pVlVDk3LARS
xecmmZ2ZMrL5RIEE+1syk/GDSjz1PcEUDuC6syWUCs1ywEesUY0IHQoecQnLmCYOeeEFeK6RJxXJ
5ZWNxXYtv2nEmjO3UgQRyLSB0QIo2mYqzDfC46x8AfW+N2tZPdruZbpwY5nYcjNR6YMpYQ7+eybd
BofOcCJEAW0P75VaZ8rXIHVorppCvVi+IU52nZsK4CntnV+BBae8/TmjUpQnBGpOBh6b78m+tcLq
O1EViGKcosdhvsZVZx4kaP14H25RhNsIENpDOYEg/ddpoqninpYCQn8f+oc3xAOXqBuQRT5Kgk5o
6XjW4x62HAXyUHpLStjDszsY7VgNZ4GZsCCT2Y66E7kVSrFbelS2Io1M19KscoiFcTuO7GsPjUB7
DSjL8bOa9ve2eUr1mFufu5+zinNmXJhkrMWmxbTjMzg1SxWrl/OSBdpAwHLRfESEbpBgbk6bgQ2Z
jpvQIlbosx1L47sFpZsfq9/jz78wzetloU5vsP+I6zZbZ4oFKn8rZAuhzk2PW+aQGT9JA3qQQfFK
/kFDRppvF737uUbYAqDZFWOwmfMTXWto2mb0R6GTCFoHWXywcA/AHyCnNBndORPf+6J1592pdglj
R+qdJ8GeWktErn/RFr9BMe3p85DTc++V99BDMFeDQwCMXJxhFLYV/CGMVyVfL4h1PNG3LFXkdyYc
ZQFwNhdFWlaWDWftpOR940LP+lwBPYRtaVpJxglw5wZrkzQzqi0dYZFpaZU4I21tDikgu+0WNYO0
EnvUOqqmCuhvgOVV0jn2lgNmgKVtphsnxUtfrGCJOj5WXjGXJDiiGPgyzvb7vFhE/Oyu6pSCO6c+
lnsa3PFZRJkYZcjaMc6hKrLXr2F3iKIp2KYVL+iS75sHq6cyFzgUc5a98GnyUVNPUt3hKdu7+iYa
YjLR6ZA7g5i1R/RNAfyIh1V7w3nutfJA62CkA8DF2Hxx9m2uNsI6St2NsrZeINBvFpbUYTO+2TCj
DO7pbG3+JZVEM+LLddCZWYCbCnw8mPYrweKTntfekkvfNLjKNV/OAPz0776eIf3QECjmvArT7DGY
+stj+ri0cFWT2ip6sk77L12ylmh73kbaiOUYlTMBoUbwnq9dDa+xYbggtmDF0hszLb5YPjcAq5Vr
Qn0QMM3n1scN5XsuVYNsfpkOUkN/Jy/r6JTIINS2LBIuxVF8BxKZozppMLtfKDWw3x6a33jh7Cmb
rSXAEYFkFUaA//7w/n6Iw5pchXhnkaZVd/S5yAE/o9FckJ3IZdDI1rQamyaue6aLpRe3oldzaE4A
PuoOvPtZX2S6FDvmX/WDSxMoG6CinMcvCFbAbPattQM9Qsi/vCTRVOEecwXskt96sD5u9IVO/Lov
5W+QZ91McZFj/LjRv0fDGDeXhPPgBKQ0P/0wG2zlnedfFBRrMfv6Sf6WMTrW5EJJWqsyssM3noTo
cG80G5YNdTdL+DBs36KAfojtLSt0tYR1U38zVIuaeW3n7lqVRpcrQ2KtsQtUxIoPpqVIVOZ/ZjRB
I0FtR/9Tm+o9U5TSFfSuZ/A34ipLK1+O0N2S9tVkSLMb/a3nqk/mGUvTluU19PfCFfYGwwj3W3iu
1dczWiqEXMe6zuv07WRJyn39w6TIRH1s5Wa570kaCymLvnaRcnKZKsewyyGrN4mYJOjeogDPQ5qe
ATCTiSvyKZftIFu89CDH/P2n3kVWRR6rKF2cI07aKYicN7HWzWJwMKfmUNLyL/99Xkb4ahuFE5KP
7CI17leu1tTF0DCARNC+5KqC0iO5sPyWugXJYYsbFvnuVLf0Rv8QgIoQFgch5ZJAtldbwSj9ehy1
tyVM22h939CYUJXKUAjXG1vjYg4mNaZCWtJrtLtmuWl6JJotJ+wHcrdKeUBrX/PX7CnVcpORP2K7
EFVLgQTIP9Ygzx+YIfqF+bKr1ITQRZKJEpdwmmPKAw04ofUsP6I8qwXGohpoOWYxMLcIG+IMIkCw
DPGxAaoKKi+SCavEt5jmmmCds9sbiS0xtzYDv5/SYLMUi9vM9hm4JP14OngqYiwxHoO7mP2oRvDf
h/SgPxVHZo3ehpZSikxgpo3KyCi6uyLUGWmq3CHxs262D4LTiLhSrSOEKHoqfEx1Bc5pi8LqT/3e
JBoYO9arheX/V3PVlXh0IjHNx+SGJrFBod0zoH1cvLLDDIjb2xW0Tbnag+Ld+xj82DujD5rTdaha
DKVdXOpwsDWDDXT6AtpQResEd7//ID0Gp0875CSdPNvFMY3MHBK1BHY2eW4lg5fEsNAIrpHrPxDO
WHOktcg9id+GuQXH2NsFHHJ8NPez9wYdcry7NiOzSsngkmu1/kyuYDXD4j53P7jhrLCqSl6yE9BA
lHRAHQhgPIV6EWu9sJLqRjMhJM20Ppp+sQv8eiNicWcuKd+gW1OGi9O9qdWzTSksnSn/gJzPhz83
YfrFMqEoJIJptTJCARWkEq6QHe30MN6udQ1RPQxiVehf7nWS8geyPDqjxmsSjj0UDNzoYsRIe+no
mLJJ07weCHkqPYwCkGe6ywnw8J87vUb6ZtSZWXbXuuMSDV+FhGz/gn7ehDYNwp9gwueMv78t4WOP
i9oy0V3YadnO1JyHuuV9W99cDl6zSWjwa+d9pamVbKb5hVq8rTLq+C4EZfi690XHeBtAJzdAA7P9
/0D4OARfUz7Gol2mqcpmb+jSfD5QP/PygPjG+wOuU4m17YpcyUTHTDwAE7Wu06XcIIIGRZRbz3ni
TG+NF7O0g+giRUdIagKeiSBwqyG7brouaYcJ7qNXxpm2DqQoTGpPFX6kUTNaV+almANCthDHHq5n
BAU/pElQfhCGevAQ5U4SVgGv0hx1hJ/N7UAoV7mcpftTIQKpvY5yxuTmVYENg4FcXK5FmHLbzY6A
hdbn1r3WlRBIBN1de8pu566twhtYb5SxBKeGLHQDypOI63+WHOWMq8yGI7JIIBrBDGZ5MhT7bLjR
ViPKMJDR1l4x4Ny5L2AD8NxvtYR8lrP9fvd3LctyDEtkUvn8BZ7A2J8BSs2195DarjnkqMkMuz3f
/yKJ7Yt3Ouv3j2oxJD6Qm/MtDMR9mqBzqi+NYcwXVRRAvHl+AgfJ1GKhrZ7kUwTaGqk9iRgFe3o4
kXhDvA9/nnCM1+nzZWXsLkZ5G3nZ1ZbOqiy9OaR11WQwZ/p6D3YQKm9rJ5VtywOIMX/tJ79zdPG0
OcOCVC+Y252pdDRmxk8Wc4khJQef+usfJ8PidIQ/gp3Pi0pOZq6ryAm3Kh5wT70ZZN6e0YrTv1ua
A/BhaYv5ApRMsUcEx7QGNSOQW3Y1gBIE5Fz89KP7YJulGl7m15w3NPL1WX7jD9wMtPc+q+vAKBIU
ptp+3k4MQ0D2puXcSS7akEpSmH4iII9EAhcLLH5bZhvlAZmcPSawamCHK9piGkm+BkEvC738wg1N
IEytBQHYwExtIazSFw/ZA26BbsylSiLjkmkfvg6BktGYhkonE20JV47wJJKyVpQuzAIgQik0pduB
tR6jdpDq6R5XJf9NPbXZHwIzlZfI0J940Qwfy03wNEHJd/YChMmlBlsf5yuc8PmBh6sYeh8bEesR
K2pDsDhKw39egGewLFM3RbMYV1VqX1OMKau9BCQy+2pnV2AZ5jRH6G0ir6xNy6aNXWsrykmbRdJl
uiOvQ6KxCHkvHI3X75m3KGyjO0wA7qbJV7gL9oZZv3RmxwXnJW96FZ+hRZ5WNixVmJHXBIJipTLI
sG421RTaN6xdsA6Ol0WBBYOpeKe8kh+VQlzOg6izsEDQKhJPaJlvhL02Jotd42iAjCbW3OqOwips
ZltEp99kOjLPwWGoW6YMJWcCJdjrfucHUqB42Z9Dv+8k18aWoHCUoaVQMAvorzNZBf6AxLzSOiMq
XTxXdcqkhrAgsGAkHRVhfTPs4XJuU0A0KleKiGdboQJyM/HcSaDo9a8bb7eFLko1BzrfHOEDx7MA
v3tTO15zViUUsPId0zqsV6sDXFU0ZrTJz48pCWrKlfvyAFdUZ978hTnOooPB/mhSNh3+dM5APoCH
jTNg1WfUeqlHVLGxJGK5NQCRMmg89CK0bCLbRgVs9tUoBqPTHPpqXuiMxGM5Dp3Xa96gXESsJGT4
P+9/HW4lNwVMA7L1EjrkltaW5zZBNq91+/vyOiposR3+y6VRyTiFuDnHe2fpIjbSjLEhaA+8/J4f
1sM6tPIFRkypCxiZc4A206q/tsBIogKfDmX7188xeLwJ0mZP868rQkxQyJfJOFk3bVUja+9DwUy9
Q5zGUaO7oYeLS+88wsUxj+sNHRRqhvO7PMjle7KwWBUe6bFhx/RDnnkJZyHfLaZZ0jOHqq15hdNg
g4TswDJoYY/b6n+ylp7yNZqdnBJ+22QdKumD5AB/3gvJoYfSS6/TBBgBJeYz7X6anDSjXQnkJXpX
dIvezKAOOWFG/hHgJSTdK5LTDpRkzgUQP89+frcKsEDU/7C3Z2awrUqFXwDKxbMPGzOf5o3prjIK
HXJoJx0H9TwL7VQdzHkIAUVef+DKffSARVlkgmWHdmjHeVzSA5+mcd97mMdTA2yF8JJz2hOxwZdf
WjgviDdLTeMnSiXMgEtQoED4MGR3z5dXNHWNbofEymBQgoUIQaD47LRdxkh+CMl0kUJ079CpIT5v
Eh/AkynrL+m+YChGzwaXvHPo5DxW7S29Hw1KHdhtmiNKykCVdFrDGSUCe6apBQr67KSJzcrNjivp
qjm31sihaY0MfDW6Mps5BesJfXJ/N6FvG0sWT3R1f9nBkD/kjkbZ7vFEM/w5NDXFRZp50r5ZZFy3
xL62dlH3DS6wsWM0gjVysB2/8yzSBakOhL/GgU6dut+YZM35iGX4THx04hm20OhTi4LndjBPxWgB
+xp+HrTbZL/U3ZVoYkcnVQz+Q3bcZYmm00o0mTvpETLbXdMepuDJVF6w5awLBlq0skoOg32EOoZA
5BLMc0bBlwecKbLY4lAF9r/As2RTN5AQIjldjKWdb5JOIDaJ5T+/ilHATRvot16sZ896r92Y5vzk
9bdF4MRH2RRqNL+cvlVzVWf9AhLqBCZofW4NJZ+4LuSiQBpzi5u9MvahO0uhJ+1C1Ej+bTrL9Nl0
l/gJ2QxLqkGATVfCElWNLcmGPr3caOfJN3DKMf08FSgpb6SEJudHebkiMf2pO4/99bmvVghmvoLN
q4WEIZMjg+zouvKPDqNDbnWakVfBbG5mUs80CPPQi0BsKkC686LAsW8/Geb/hngGmqN+eN9UTXFP
2un6h06RL+kvm4gTcifQEm06wwy9nMVvtNGycLC046WfqacY4Sei0FlMStymbr6mmEIxBdE4MPvj
6/3yITj4z2wQKOUnH0I91EQ5ATRrQkiN4dl0eGY3hHxRlBNhWltUCGZjjR4sO0SPjO9ke4QBn5UI
S+2V73DCvxZEXpY5cUIUfNkPg15KPIvlGIry/wU4zPRArvyoNEtu7U1DDhOLpJgukm+8NQPfGHpQ
KOyK1W9upPEG0tE1AslKlSsXCJtoowo56eF4KPH54uafCKb+t2X7Onlwvz6FzQiN/zwSrPXezyxL
Gwh9YV6hhhG49HXCrObJgoCBTAopL2O7uhYXcVYE3qqWelTAs3+1baUT7dBJEBGixBxVWP6xW9Fb
BV0TPUDSXEINqv7W9WvW4KiTwtWW8PapYWcPH0ZSZCZX4qtXTsIFDul72SpBqbqiRx5zOcjBxAEr
8YOzzAR62KtdzkWau/A+yNlzfLa0VSqyQgSvNpOe3XTlj7ma7lHcjDshkvHwXmrpBtRtG39HoZZC
3EIoZcjUpKQ3zfp2y/D1hhnwbPKeQQeYB85TcwfigZK63NKpBwJ08/c4wKBuPJyipaf/O1JCEcl/
6WtMUWpEwKWotdphNrcEssx3DDkQea9qL+QElKsjgKMS5xS43I/FmBcnnP8a3XqPFAO6R+nL8Zfz
REsG/rnvMUh8Mk7t7SDggH7ncqxY+uGLrXfRU1xcRP7SoUwq0SW1SmFWN0ZL/aGaRBnFnIQODJgi
1697dwv817Po5nA3SD3onNe3vg5otkAGjuHkFLDYHP0XQy5X8DYVmF+wfQ+J+D6SfIbir5+AkR8v
dM2bVRQjBIjtKctJ5sQ0VioVkNTBvflrzF84BykHcrl7uVL3cpZsAdpQO4bbWpLny9bHvhmJDXDe
zaW8+yx6LY3rrs3GOrEkl+/pEyxMV2AnEXE27aV7ZrLhn1MrywNi8GSamqRAPQ20JZy3+SXi53AB
u6pdDM3ZIEGGV9aLwgUrWGZzFd8Gu34WA7MZyBEJWqgzzWQRaGc5I4NvCD3NhFR1/VAyoNv9rJcr
89snCKsf5M+Tz1B4aSSsxngEwdYRkLwAE/S7RHrqdqmBaXcb8Co09oInNoMRCxtY9yznNNTaMWQc
JP48t9XEXEvul1s1/iy8nm/GVCyUc8+7LLizGP0UjkfSM/AWYRLPijBBWFNe/nDGDXMZl2M5SOBe
KRdUY/BzpEALW5K5HzggEYN+IBPdbBegzoclnOklyN2J3oj/URn4Q9e58r0/9FCNOZ68pARyl0VY
SDsl3GZS6p6gsxmpC1bH2ADMuIZQy/hpcdyPRmFXTFc7pjT4JAcpSDou24Ntm5urHs4ViY4uk3nf
7kjjQDRCIvXmKavxMVjk61SUx+Sajkt+q+zUswCHt3+lXooMe912p6pzHPRDJ5TcEXXfDLgBMD6i
IDG9v0mP9vbL1V3qU7eJNTW5/3EIMLfYebB4nc3DsKfpk9XlGRrRzbTrrB2HyXazCdxti382Pb9u
1n+w50HqYbxjZNpLYXXnJ6AA+e9KHjzyRGZiOKy8N37Gq3gggAE3fAKGjNwCFHZ0xBd1JSIBM/2c
tvYAUnkjagMvOvHUlJe/iMkRF02PdtXuTiw5GY/aHw1HL2RGYgydlRDLcGgLki152UkMLxc0OyLZ
2XQh4HNfIE37Ue0xA3Nl4mD+IYWx1aErs6DsQh6SrntSsVpTBBBicF6Ar/LC7DAklo0wGkzeymWc
UC9Ma/rujcytsNevOLY6YFMmGhQkVjhHW/NCZHbZubixH/apL05shQGcqO53d9KJuJNdLtF1iir5
KqC6O5UmymPZEB51CXrKDDG73+OF2xzj0FCB5Wuo8SvJe8OmcczOKzAjYSV57+Akx+SHmKVMd4tw
GzAg9Wnx1ID5pJiD4D9yC0QpSH5/H0h1gYNzjAI/LmOrLAc5GxEkPvAZL183xHCE4fcQs+NeCG8S
ffAE3n0G4mBo7mA2nFR9XNLwTRMji7ag4evf0jdeTw8bPukrL11rtGuhfrs+bOxrE/8EUHJhvGj9
KVI4ULYr3HKV22yAbcYy2wkT+LNf20esFleuwQf0tpAUPHyli2vdxrvCFG4GstT+LAjRVHoiptUG
YJnFFlY7td0zGlptC1Onf4ELbW+yuL/AQLFnuXXlRNvSiSw9rkHLxNS21CP+kX0sUIf/n2oyq0TR
n89ecZw2wFM4zBr9SOpB+Qu0x6FPrNoT38V6pn6Ce5XVdBMmaZsRgo83XTVX/iyJyn5Ln3oQtB3f
+Rf/xTrl7VEB55uYteVfTkVVOB2WRPf00Su0PpVXmcodjcHw68PPv61glr82mH///XhCvcHj0rQE
zVhhRP7jSO3R7QiKZ9rZemkuabHcZgFnRSHY/U9wYl5gAHm8qvgjvKUN8CxWwlD8L3QCYvSciRdq
48wBW/kDcoBzZ2ozBoHxp/SOo4ijQjbSS1jRkRdgXXp4yP1czeT2DwFysZMVUT15VVvb4J5P/a7k
+vd1spoI3/R14AioUpAdk0BMELh8ip9OlM43ardh4/Jul/fIz7+dhfJ0wjFij9fPcEZMmaffPNxU
qfVlgQoawwVJr2RiBkdR9BruWD9bSwKZ7Bjxs+snLlyDkdE9qgic8x3bx7SRrCRgCCi829KX9YrH
JT4uz9ihL5VVs5v2KU2zvpQG7Vlq58Yk/x5zitnye6pJUml4zWz4W+vRpSlqm4Fjn15byUdGqJHL
l9H7hMnydytEjh7uCvGrAE468RG7LYeePaD9Fhq1bGHPUYUSr0m3glK29UzO7rDrIDlsUMrfR2BE
qdABBx4yqVhto+SP7qND4L9wNRh3DY/AlYJz4m+vDKo3lLCB1TNs1fuYVMv7oiekCYggdrq9t8ri
QNUQ0npVc/oZh2m5Vw3k3kO8aQpILTgZOcRFABXQr6O4vYnqVx+1nbhryd80/TBZ+wJhThOXBRnh
021puPZFQhcvt5bejvjb5gJ4X3x6CVuNizqEQkJ2AjpIj+dtYQF9DrRqacfhFd9PXYNQ97ZRS3cU
NYY8gR7GmdVOoHHlhAzAzkFacTlJG6YYyzwokC8bJH8u3MNjFnvxR8IXOR0iLnEaVbU4hZgu67oe
NqDB8PUGDeIPbQsPC6eKkh7ZKFcIvmKT0GAQ833xDeLt3Z6VeOkPsD5aWVqR8vO/NbhaU/Ts44Zy
+2UnbpT0zH6PF901BO7xCQoWdKnbhbOWoG6tBoXtECVQ7BmuPr/4v15kGpUichuv9ISZaG2xOuwL
6QI/9d2hAVaAPv9GXs4dh/byNdp33hkmIRyl3PItI/45VJ80c7IQyA94ac9Dny2gCTECgSVuIM+K
m+12ETSAojVr5OnoH9Q/4sUhHYffiowDnKkdcp/q+JbaAS8HdGjrn03Ilq+nu5zpSOeVUpUCSZXy
B+xO3JD9HOMuZZWCw29E4+KyA9BmzRBtT6J0pfCw5N58Fg0umCuQarl2XcpcZVdEjd3xjcJAwzD1
HCBH/mJu2KnFy+w5JJSfMHqfX8+YLcjWSpFTqlTvDRET9Rs/AC1idosJryoZEB2nSbS8FaUCvgzZ
92FmlXQO0Tmrzsp5ZfB2QxkrY3E37pe7Cz5ahltdbQpDhFXW13FyTfSdS6cF+AWkBLbDkNnZ3VW3
UxChVKJp4bLbeT448O2v3hhIcvXHei5412u9aR9B0wiX8LGQPIFQAENS1y4NWj7mDEwYxGDPNVjI
atpJYgKmGwXLA8CZ5CB/mUVcz4lh0/b4kKL+BG9Ia8cMn9L6SavXb+Noygh4XMJ8Wpx61XnZL8cp
P81hdOAPtI5DEWRahsud9lNTKxG+wGiJRokZw9EWAsxsCb1sdMaz0+TN55npuAr2dx6rqRDAnpVk
8Rf6ZOvVLkUTbwpSyms76Nu7iiRmIX2CuFo4nYXUUzOSX/dQkxBHLEiYQ23ZT1T4geCweLDg8Un2
R1YSh8DiYdxi598vAPSb53mqbDjMP2aJiHqwi8u1huaueGB12yP9uysYk6WPjzPA4zrjZha/ahkz
BVybR09dyoY9M1Tf8OdYzDN7xNRMF/rVwTk7BlQCckKD+13U9dKKanvYs693IMHiZDvkAL1cgPI9
79TDB57xZbCYi5+XFa6kquj0NZCFbjWVU/5k2o9CGuUefJfiLPjtf9L7vUpmBZ0z3NPjz36j5Tte
MYNgCKKkv/00if09So8fV0CUg2pKfEWplCdCmCewF2D1t10zFGPpL2t9Bt/ojRXIJlwh2Q9uupdO
Ohhh7XUknc9bKAeXY/+SC98aVPyVnlXldQZzv+Xn/Y8RXT1+KyttjKREXCDZYdYZKlVPWgN6MY5I
KDmDDwIqQxDyMrTtJMOn41R7soML43eOuzBLXFobSdAeaddnBi+Q6Vnu1WwftN5EFoX1LaH8MGca
Zx5idmsy1NswSEIwvsorHdjoydvY8FTSdFTI55jq+TJ86zgUh/x8t72vdrJ1FLAn2WJslSIdGXdk
sMCM62g+jGU9tWA6N/8j39ooEoQ3Jt/Et9xcF+hGQwXlx63aYrVOGBZnl3cMJO5qnYbq+AQE9BB2
pHfmGRE1zEa2yWkfrSzuhql+D9vxoL6Hq6gd93LIViII+4HRrGbtoM513UL5Wh8jxXi9wvkXgfFE
IieHgNFT+squWyc5esDoNhpQ3ViWHYVhBn8gxz/JdM/IIUMHlr0W66ZK2m0sAO/pgw/j/VipxKxt
K+G1MEmoA8OwM1bEyMyyaWvH02T40jf9yxIyy+CqWnDonOiDyDkTiJ8nV0d/2UIXKLpGEea30VHb
BO2hoQr+3itv35gsFetxFvwyUa08/P/BCMctfk1JwdASJbMTo7PGma4GrmUjGVD80RuQswvKcIM/
HwSdL/kaDvVcxranIIu5zaGIWERT9Tyka0raJ+iFWobHJHHrHmCQDW4HbDvdn/FzZmejdkEZdNl1
I585hPx2u0ZIs+3wnUgeWCjk1cXSuTRQRUbKdwHSN9NEmtNd5pAaAkcoea1A7zggHdRrVYlhUcfD
8kMJTjRhwol+LM8iD/inH7/5r6gYKg3FPU5b9PYkmH5DEjELKgm277K6/L7gU4XoQQVUGMNAWHQ+
QTYcOhO1PG8TLjz7UcOAiIg1OToWAvsWFIKZznUGz+izD6wweL/b8dmrpYtqHVHRl7jXv8tX/+gV
pGRe9736UIn+juYA5UYivIA8vtYOqzSI8hAAta7uad+ERqkqEHyD9aBWtBHyaOWXJjcycwPjPjdx
1Jxi416o2xnsO+l+IBVcrHlzfzm8eW4alKUJyKtHa+4nqMBG/wlMYHeHNoVB/BvoLOf5yKnDNCzI
MckvRjCpAnUO8yUbUHWc7qha2vRzJZI882LmgTg8S9qRbKXrv3A/rVFMw0dRX4SQ1YKG0NKogkPQ
j9hvhr9PZ8tfV8OlhWUbvQW9mO2vBC9NsZULOBVNnI0j0vvrCWxesI1UK5XPBAX54Ls/oViLarUV
vY/SpBpT2qyKMqZ1SC2it1k2w7okdYdM2/KLNIKyU4kSWnaeDFB9i2mLse+QiT6+V18fHlfhQ4gJ
3Js95eGWbUKqU3JQBaw4dyPR2At+ZicmGZzdI5WHMK23AIuHz73kTthnMKQU35Hv6pv17reTn5cx
hzHJQn/khQpofdjg1PzjbaP11+t3qXaIFLRbbpA/Kr5egPkUHiMGN1hWS8R2wp62aIq6lGKS+/G8
1/SRH2AIbNOAMZZB9X/0fk/Kz9n1T7hKv53JtZy28bXWpssL1wdtV2LMGGOxAHbpeaWur/1w1uye
kIf01EcPBmDlcVnHKwwGpqv3K12mIBjDyd4lct9jblz4zr9MIHMWtjy8azcOQ+b5cDImLYBoPOE1
zdfXZ5UC7XrROo4dNVaq3AzIlemCMWxHQ+WayisVcAPDv+QCkYGr8Mb96JvPk8eGx/cTmvBkS5lT
4/qpVbRdxF9LXz96agCvttG8ocqZYlQ6ZQ3Vo/yxlrozpdv3lkwOVgMtQyJrLmhPsBbLBKSnEe2h
OCXkiV6cb4UzAwqrSLPgVrYAgUeUEdF8IBkV//3hRgLa7gNYMPNdLrN837d4f0JAH93T4AOpkuoP
Ujs54YTPn8Q3pjvaVJ8wKJt1iIxiUSe8QnZuyIB12DdcqZgZKwVTJzLUnEniCL/ITEHvxcmRiA8M
b0tSEaahiiieKvLlbTZKdDuA2eN3Abb+4lQAmbv5/Bq4hUuP+r0jD6hLCK0gdPE5YglQafm6GS7X
Djfk4QUoPK2oSosa2du8MjCeeaYqy9l+ZrseSmtHp+e5kU2A4I8rjjE9ufWDGAtTzWks/Vcebd9o
BE9tSFxF3ctcYSnOtFK1GeOyCTViIQ//dRYbjuRU9AefY4RN50f6zbYbePKMdPLoPnlTnEWPeiZV
vFFxoayXq1e8x4WKiXbJbgXsdNLDLcSUsJ+KAWePGQvG7Cd3OrlJhoCj73j950+D7XrgpgGoARsm
MIMoH62tHSttrYNA8Pdy/BppNIry3+hxWa49aNHh36xZJTf+kvQ7kmGF0xTyiN5LpAZHgOuwrpvb
9ndb/CtXBQ8NH8hgCQzJiLYHwmQnhxeHnXZAPyV2i4N4hrR1rcxoj5qpOJeMj1R9gTGTc3dzeAdL
dVi1SbSIQiuJKexxyYDt/FsBiF7A1o/FgsvernySRukP190nr/uOT7L7CUv30Lm0/8MY7Y8vSnHX
Ju+S6ScInpwNaZiLvSzPthf/h2b5sPq1jrFN9sGWG61EvxLBTxV079GvgMwAG3G52zxKnlKgduVF
DUtinrTv9TNhHFmFYIZ7YNk1lfedHtAFpCM+tyFBuE08dj5Xid4ui3M9MkUInE/RUAWRVcX6G02D
KlWhM3Q2Acn9lARTxFX4xMRVFZDiRUalkusebZ7Bnnub0+HZZAsUsdjTf/SOcz7KMydwfUNgLyOw
AM8kPx8G9cWept985I+OwmJnwWfO03qfHuT/siCC9a64oWptr8si+EBMa25uG0nH5OwJAMw4lpXl
Hj1QYg+/zYcm75oXQ2csmKdszebsqXD71uhsl/nvpTxI0S8rofljJm5j11stwhfYCBSjZ4Eob88P
8R4JFSjfaZQ6+gUf/slH9DTT0A2dMGcbzpaG+/kV+nc4YlzoxjX6OD2put93axUueVCqS86A5MVu
NPqFNFwGkQTcDzzBVNW/S0SnBR+Ft/mwYL/KZpDSIEp+wliUBM1hzJ0MpqBhpiHj3OYGOJQeW23u
MTY8FNtCjp31sht2H++KnqaWEq/3UiZrX9uelYYk4u/YI9Wx+jt+BAHozgD5dXJ4KK+IBV+c/J0x
e9jzeseH4K6ER8/1Vz8OeOFZGABGPgplK8ZDK7lWcKzI6aqx55+GnTemQg83yDf+RW4YUGPZN7xN
801oAljadlKgOXRRjQlg50Z/DRlgftvqBT79lWMDhA08kRsyPArD1y6UnD4TO+f3+m9wsxRh3fie
v4yh7mDy8RjnttMyx5iTjKebGlm1R1VIbxXOZM7uB9DQkreO/T+pYBKoZo0lR10ThZHe2eyIzfTm
6Oy654lKb2oyisMzbjv4VJEAk6c0HqPjsbFh8gxZCcbPSic/0BK/e+e6pRaOqysXNEtfoTJrWHCr
v6BfE4WTOL0wcMXEnO1RnkEVaS3sQwCpbK66LHFiHDgOU7jlHjNAoQ0bzdpK06n/UF0Yp9eGpNKi
OBmF8KqZ1aBIzmYv6Z9jWAejPRTXZTyy7BAWhFpp4xbMdHCGmPPA9ZSg3CIeFF4B0f4HV2QaDChq
lhCrG1JcsvylpU0IIo/EIEBWJeQ+9daYo/IVBhfzgYoTmORsYmd9CjcQ4VyFdFeup19Hw2IEacro
armwS7Mr89zZNRVKVVn1zhO8CxsWVhpOTwqwl59IyCVfXwB8n2KXa4kPM4xUTY2HosBWhJ1e/Vzv
7AvGmvX+h+l4MegYfWdkt5BvMDGgCIa4CvuMjRd7dRSRww60vPnizt3dK5BHNyP7BX+MOIomgXLB
GyljDW3tToLG+CSfKqSLWr9t4XcBD7Mej1RtUv0ZwNZhLtg5OQb7FEdcWOc2Xo7+jkKn35HKMm/o
46RgdElHWzWQGMYCG0PzFeA3mAGGcrjCWq4udJSRmGO2IF1d/NHRYZKcNzfvEsoz//IVjNBdVGxn
Da0nXt0e5noqAq/CvHH5Kw5f4HsMr6heEpF6sZq+Er+j4T1/I6UcsSEo/WU2HeoT5kRp6vjTSRES
YPPQlV8KvPerQpF730I+gczC2vMuB7SoOs0tD+OINBrPql2SJ5mL8ijeCMonTXxn1Y0kz1tfzLk4
TEGyegyLYrR6hUGxvRx62IRCAlF7HTOq8DDVWE6ODCrPHr0Anb0zgy9QMOLY/AjLkEb6zMSGuH/0
wZBaXRHQLfboOk3Ov1kHy3bHV7C9T7biR8dSs1kqd5O7o0gwAG+okLI1mzCjDSrRV/bJbpsFB+ob
a9cyycfdm9A5gquQOkM5UUARtlrlOGal4nn/pOUeWe78hqKC5iHbb626L0z/nS/0kfeFbRUIQ1At
zyxJXqaolzG2mVrWPSslZq6SFGMexaCRG5j5+7ANyXFu9sdvevH5g19AyDRetz02mUD21c7rPi2t
Us8x1qnuqSktNKAe8ttS5n3eq9WpriRXXipWcNqBSYIqNhGmHksJ92LmNic61zueDhPX+5jsrkRi
7vwadJvmc1egggh33826k6qvAvju2h2YyJdtcrgziinf9nezpebeaEPyDUcdH0lpcFmRScgj5eG7
O63Cx72KXWv2phriRKB71F9C6Eej5dHlt5cf+lKezZA2mwoVSAfBaOy72Y2SdEkBXVxmBYFTuQ5d
yI+AuYs7Zrtq6uyOe0Aqcy/04uJScrFpYhbyPuBwwCAmtxva2V494t/GNrnqRgRLJA9MRvPlsLVu
O+WwYFN+7dp3mTeY9UE8JuHDSxykGFlTdq+mogHUw7PJqxR4diK5yHs77wANl6WC4BKUenRqfvDp
TT0NnzyBTkEyN4VYp5Radvh346asM3pUo8E7ayF7QnY8/qpsB+5v8l0ACjzeQllF+xlifBVISUEu
5dLluhtFBC3pqazWFJ4bFarLcXMcGbMep+QnqCzyrtEfeD8geJd118OI+kSDKgMJ9cLSAOBtdatd
CT3SuejX99DKdgyTUZsNM8+uVAwKLAUg5RwB8GGw6LgiGiJpbouXCUlebIRMF59xfljxCVNjvrcc
oXFVxHu/kA6PJemJtaVGIVA9eZRNYSLpOt+SV2GdP4kEc2I1VBW/JqXuZuunJ9tqVA0n2LNwud+7
g0c5aw/dqY6+RsRodiz1mdGKWtbPXTXBMOHhPlkoyTOxGMak46WdCjvLju0nUPW9IEtksBwTLan8
BGzCZgua8yE3rOxm6GQTkQxfstS7NVy+xzVO1C/wBPWWO4y1a84vYtKKqpr8ehij9WTlSYYIAMxl
grH5BahoURpNGd8xqqDhgeUaOFIYxQN9czkoT31l+xKcNaC+K005pWEtsdzmbwWF/+JpV5VDCLiO
eQ7DTchy8NdtbINZFEvCKQnuGEZR6YozaUcKi/cCUqC4lwwpoVDMdoN5E+d7sFLtxgsyR8G/Oxbd
C7pJP6SVlU0TNE7LU5LWnvnilDXtWH9PTNanE1/qvH4bsU9CjGzNZnlSSt10s5WLlhXw6P8yjsWW
PcHvyDXK2sWe77two9vo5O4NyPyewsKe8pLrgoGQeTlTT4h+cYbMU3VH8l5V6GT69WThnFACv9Ep
+klCe2dVt7b8Mw+CCyWn4ukmS8Lwa6ww8j9nPu7uc/y6wlJyGrUl/YyadpJhIfM6m1EdZE9svvOj
uC49BURw86ZAXQnwYT6KF21enOgnxf64C4A+U1Z+QdVeebavUZ6qgKvAyNFBXlxRhEMddMiJ1fYN
12H0reX2DvULiyzEfKI2LbAR2RKq7mFgW0vUEf2qUIR2KGs2/luA78821XQRuixDWGu9cTgHfs10
SA79XHrN/T92bkfgrxvHHrnP51cPjHWTMaCIoSMx69ZOsHOjzhKDiZ2UymRp9qU5ZFodV37mofnF
0NvAYVFgWVd82i6czC0pPWpaiaIM6MpwcyZbdmTWcVoc0tCyP1q7505INaFw3tsz9w7/PYDxm4xH
8mn+oyxAGARgsJxFBxBIcn/2tzYTGiXpl+Zb8AhwJBU8irWA7DJdYPJMTAMhlbDpRKU3xB4pfi9p
JBpMbEC8yYE72Sqe8++dClBLtCjTKoGYV96IGVQMUtTDGc9CiTDIrMzs2Hj17pdAevnTzBnnLvj2
upiXKa0oapcK0+ZAP04oobRZkfe0X5226Ja/sFB/M4KvrnMDZtusNymYrF8SxCYtAg7FbS93xNZV
2Puan9ZzSqaWz7dEbYryTSWgUXzQyZTjoZN6Rpn66ck0ZgsGBqULouu2QXpu3wcMP80llLlmtAnL
3JctDTZ5T+6xdTR/xf+zgFN2uQqXb5kxNpTsiVFONWvwYglNtP/oMVTsPNnz1t7/lSqyAoTPr1gy
acUKGM4knyxrbbcKhzTKOQ4YWauhw26y+svRrTzNtI0hfbSsn0eGcm3p7pjoAyp/sW4T+bEPpnLM
2hSA6Eme2Vtt3a0e9cD/roIZN1B86LLVxmOM5SU2Kdhkb5bXfTOQp5PGaTr7V1YGpj+LfKGMGfwz
vNFSCC77+YZP2emU7GA0YEykzGrlXnAHIrJ3SLAGxdeFgsgrZNq0i88IOfwGXcw+4saYTuuX5s2A
qSmc08G4j56MyfGpStyPUJbNRe/3VSXeGZKigWG69FFvxMjCbqfE1j6AO/wujYE+mYxioI7VBbTM
g2v5pBT8LJXctCrGqkmSN21Qt5DUSH+IxFx4xqWxRy7+Pxu1pYN/uLeus/6ffCTC11xVpVW9ZHT+
Kb25E7/zDOJU6Bo5LyRRmn8jJH/EP8oD8q7mBMk0spWAfn3whma/SFIYgCmSO7X9w89/zo/BOj5r
FVnBPWpaZU0nr4w/jLhnvH3yvxXY4/I3dE27xwg0uAGFZX4xfzO12DHDSexzZJrIQbpLxMdt9tjg
9e7p8CjRWTtnMcZyJPw6UL7sKcNs4T+N5mNikftO2EYfYV0rhVlGgnUFeIHk165Dp2hjkSJ2aa8g
/fgtkCN/5QkBQaKR3MtuturV8IlOLRqy1s+eLjfacfk66Bxjps5xTwz1Lmh31gpTZJjsPs109dBY
u1Byzj8srkqK8UPrpl4QgvWtu8JkKJDme+J0XLdstvetTRkGerR7mZADpKCoeP51zKv/Ar0/FHug
Dl3zLwiSegzoY0XvlFGGIqn3R4fpxXXih/ZcKoOh5c11k600+uu4BJZJjtCNMZ1OTA7up6qRs6PO
8fCfgjFrilTJU16NVi/0hLxhSlXtBuLAHlAJJFVb1tobcd4lWIc8uL/07/mlXVhucdJLpzY4HHVI
UzaT7laIbk2SuCmMbL4HV5qoeElSOkQ8IDydYdwpUSsKamICquD6Nz9TWfIqS7u35WFB8fKSqf+d
VJiM13cPbYifVs0eS8TYvSfd89K2KHy2srDJf5NESF8u2q87QyTciEiRCcv1+HJ0KUJ+vpPz/93F
UCQijJcG4uTYrj960gcol6JUyLz0ngji5UJ60R4RFlhHOOenMehZGgLQzqvNamkQ9gS8vb85X9Xv
Fy/1WOmKGccO6cjUJ1llj5Ewox8+FSkeobKiEA2KdvyJcpyxfKppj3byG8+A9BYfPyxB8h5+gYnR
adHSy87Q7q63lS/kbbBZBNIZ35/Dag9UcFEyZaji+Nwlo2Dh/JtbX9o4RRueCdhtpTXcinq2GgEA
ju2sYZSuRHp2EZlgfI/zN0u7rxCprqZTmxR2ozOGvY9aEyUVspMDdTkBeMCiQTHEQ5bXXlA3kRZA
qURnfMbgpFsKnN44BnUvImoyOPO7nZqvcJc+WGZ9CR37Nbe0HCQQiPfAmRRWKOHNm5T9tVavoyDP
6jWfIrAa1p038aJ/3afC3ZJ48lw44BASlkyGJQnYabT+CPneuPK3aNuG/U27gy4oc4J61zHsdDrf
yJh7sZCoZsZe3ObZmQGYdLltmBDqdLI9iyYQdUT93ZEVdXBNtFflIRlfgpZqJSBHjgvGSb1cOp9k
yBMosGHQ7256WDNqpGU+MlAIiqiEbMtKdB/F971n0kD5jUWWGq+GsEVX2mCsqELYxAeFVKp3SfGZ
iO2mTLLd/3/RsawuUMnenFhoeDgV4dMsMVFPGRHC/Kwb10YUgmUp9eEOWG+8ox3VLV8HmoOYkK9I
cHhlgDu5h9YZaYl3K4i7rWDiGbSczetx9ebZVVSZVfyfWkMGKtYfbANXkdB0Mi3jA/30Z3i/RY3O
u/TOQZWri8WvR9UjHCrcBoJ0HOcK3PR0+9DX9DUtbWDrdiBIPubTFsZJqusy/fEnm1SpzWS1yGhR
0SxINj6LL0Et3/MmOUC0EtwoOpWcHFZnpX/01lhFIJ9qa/qMEpTclisOVhcHQSm8n4xAshYS+qeP
6r4IT4tngtGfkGMBAQ7ucHUZFW2zRDu3150e7HTs47vMfTGMYxhENwhUJ5dbKd0nSFUpeDvzgzCx
jbZgXpxYCEK/m1/2iGZjdHOFaxpE6oLAwx81fpaL0YVOvhY5NNW+s9fQcY+38/wgfBbA7FwaMyXW
kK+3pUpGQk4TXikSNDWq/nFzlT7kQIPL4G2Yf36nNHt6ps4LJXobdb85lkPPRJSdLnbo3/4BXqPQ
h5AtvcNLOzXNaPYmY3N8Z30OwkFaF4uLVwsecevDtodTNXEKZT+zLFKKpgPUPsyJzys75EGtuHAX
kkDheXH2YLh4w5Qum58aAsKram0OjbW7cRD9mSTIHBnyZLkdmHIIb1uBEJWsjJMlN98uZBGKB7yS
O7OoCSDLaek18lMlnM/NGREfvmKGW8aoDZQr/Xopo6aRTE2kHqcCpfL8jM31nIZdU5lQpGpDkrjX
nVOu9GioyXYrBwmnkDx0DtdN9wB80Nx7qZXiF+kUaA+8+x+kIA7BbXzUY1HEjb+yfUnlESrma62v
qUwy33inQUGaE5vXhPr4XU/0/aO7x20iiynagjz6jYN6tXe5EkIyDR5kgWcdtNrosyzB67DKVlWv
g7YPb+QT7xbjrBOubYGHDZMMJZEQ45BPDEdn2qEQ0GnTl2JwBPdG6nHjow7ISlmZcDSl5omVwGyZ
OfA/0peHrc2S5iHJscU7zlSw5feRBxy2KnP9992cNA+d92PL+c/+XrWVtQFR4oSTLwobUkWm8syq
yjYpr9CcgX6GmhL0RksR1xAYn77LLsUmxt/Q95w4vkQxJNdjRU/zoQN+6J2tjuk3JLDF4L3Xu3yh
spR3RooohLUZfYYHRIFcEPXx598r37+W9vjiaOI3Gf0bfA5ew2adiRNq+Mq/VJDnuY4qZLxQPXl9
bGJjZxIczu5KyYF9JEWFj+VDv3Rwh8oNHctA7Y+89rGSE6Yw+KDPuiBsY+qGkBsNMAudbuhJYb9k
VCA7bocYZ7A9r4ml31q+qGH7sOs7U/BlrGtlRgFjRWCdW9fcFZ+EKYMfmtlyww6alnH33TDvREGy
GvAsMhimPIlT73KZlwrF+XP3Af/urTjbDr/FGJYGPdW87bkT1CdicfU744IpK8r2FRs+5tUVN7O7
IkFI41r952l5y3huKll0DmdK2fYuMDRbALYmV4haGtWX5XVDo5IbD2DT3EZkAwVHYum5Nf7QBiAj
dHLEjHSea0ksddV6E76yFLnXhEKPg3pJ61XjFMt4lvBlYmA2HRP2Xhv6LZBF20mllCCNV43vO/Z7
Z559nlfdYtmyQDT13AmnS33RBD/drJz+p37jRdDLOamKbRLS5GwtIwMFQlg4otsWA8kEi6n3tsl6
qxTiN+Y2wL/+kVtBljiLUOqbXzE7nEX5WTDYJdLgiXirDYT4j3JpGhNv/hLZHYkN7Wx7Go/zupYo
lJoK6GVgZSB7MOGAYfFQk9CK84ice4XLGsPJKj0OjtH5HxavirJFzU347kClEiJ4x6QN99bdd9lX
d5zbQHxOQ4cGYxoQdSk63bM8myluVMaRHxeQNpdJrOgnNXy/F4EYHjRcrOPa3GTiHby/MrR7W8tM
AXhwz783mkGbftSvEQBpecxAo6k9M26654BPK1pawb71+Rdmeu1MT/Wyel387lUiGXrqKGlctg0J
+Cggwwgs0CM2+vxW01dss0Rhs+vQ8aL3nfaM4c/tuwqksR74pcT9pyTgYE8LB3FFDZY5jbRiDjQW
/HXiLOHROWr+C5sSLgYYlwso0wpWegJWCfRcJYFVoUjKnLIERXgy8DX+Vx3y5yJW0kKegb4ZExCt
D1TBav2o5zZFBicYMIuq8fSDoN9Yu1Bv2GmB6MUBwFTth1zrOBZ7mhyw/hDvlmkIJtKrerQMdOM9
iT7bpfBReXwCM5+ZcARs2JwY23fC+b7ABwUtGfqcVIXr5gGi7Y/+bmIHmQ91d2rfzAVZ/RClcdAm
hzCMrlvpbcPVnQx652Tatuh9pT1UJwz6RdrfjpAicOcwAjy+GHzUXdCh9EebD1EYc7SJe8AKFuo7
ybVwX7/wEWCzzUoQmD/r1Nc83ji6qhFkHirxHYc4RgPibY/c+UQr9l1d6IZHZ7mgDqn9qXNIiXfs
zM7V4slfBjPGIoqFAfV3iYEdH2DOR6ZIb1/oeMn6YHRCplRmDh71W4F9NC9XNA1aXNEwPvMPQgq3
WHZO/I4zang81K3RHAQ9gnWZEjCfamE6xOrmIn8V6zSK2xmArTw4/7E8+pOHp543vHIQ4FZSBxVR
ZNvEM4cAmjVQVPm74XY/wx8HPlVKQLLNYj5j4cW49GCwzTXgj5XIt/2v6DNRpj7aIGwc2pWkP0RT
rJQ+aaeh5mnkoY8yWntaeDwMaFio0PQmw7BKvYcqfC6/dVGL/m0rS/pghSjOLv16o6RXdn+sYWO5
OPrFjdHPwSUnZ/6Jxuelg6YTAaodoLfPbF3aTL7ckzjXG2dO/dCzKgnZAqI7TxWEXl/ZhLbC5FrQ
mkh1K4TLrkX47FuCmrNGXOPc7vhrv0V+tGBqIf7NN8tkfxyj5MOY6VeRS6siq7m6gBnljNxPu2tz
8q28GvK75AjO9/VwCxDpUZYzXZ3/q74mD7W3JOfHVmKXPBCSdBCbA49AUdPs7x96FYkvv2hRf+Z+
EodrKEbE+Jpkrhpuk+T07lAa4OiQbaKQapYBNckuRxZuz9bDyIksnqbo9a5lDWud37iATJQaPgL9
Pw5uuG2y5eyF5JDn6qa+MoIeKW142l+swTFf2XULB5Jp5GaaF0MrgB2MvDRJA0Os7CyXX6oHke05
ZEW6n6/+pVp3JvXqfVca4QycNNAcqoNxadezqlZG8q0dAZZ/b4vFzyrKcFaJs36PvIFxpCMoCPJd
TiXxGUKp/+zy8+pnyuUFNpIOw1Y4z/3RxujrCumYweR9EaeQYlTb/uzNAkRkTcg6L4dCDl2LPL9R
ZKES60/EMd2ET5cSxkJ1xWuTM7H6A0dmPRjPch2waRuHJSODaHmhAyNEc/a6PXkL4TkS/M0AA59p
QJR4Jzs1+FGT1KbKDmx2KxdK6rBuuDZcpmvbYyxqw6Gnx0g9giQXBBQOq/VQn6WX4JKY0pU1uDYp
bkyB/rkruKbIuv6TiG6UUWzq081KvzFUsZKpskri3AIv4/dJW6rtdCi1l0VY4JVJFU+7DMdLnSv6
zhvJOfl51iIw2Lh2uSrMe6btlwYCPzv3mO32LtFY0EKPAYzjVMH1kr3TovV+oDLqspFV0NgeS2BE
14y7AoibXWePHe6tuh007hiYfUCLGaOSKtTP26/YakCRqsf9tl/2t1M8RZvKSfdtj6qCHPkbw03u
RDfyTjz+GvFg6FfMa6gmeVhopmCM9/oLa74zvjbna6vmC/mIGzWl8U/ALIsSGe9l/AYi1CAYSx8K
yPAg05pVuHmLSNG9+jyi/ihzGAhQTAY58VI5gRoCJQ/Mm+6Auhx7CGzqhMFWoLJFNbTOMtpV1pYm
tVA14QKPx7Sv7bZI9x4qtdCTFojQXrqJdTKFb4mAL4ATKPXCM+HHJ4XXYKYCJiClEaToh9WJx4ne
FGWK6Eixrhi467oW8ajIHHkO2/UE4Vf3iWrT2ozr6Hb0ZcvgJLBL9jHMeWofBWfyI3dK6J4ELbEd
bWP9Cy9xlm0ZW8wO/qDIPMcsRBY1dIVfsbcELq68yn/u5JeLwdSpSeyhtCRux7z7On3WJm9DKPZh
Daz2zvqEYtx58uKSvscyYuYmWSWeIRE1bRgdoL10Bp+6IjtEfmP0rI5FXpbXiLjhujEQf3K4Cns9
QmP/foRjpE/xpxMsZ5ztN5vsSlw0y2x/6j6Zvw9fEhlc7N0SG2AM5ZX+cuBjBSiqFHHZ+koKf91h
IiqsN6lB9j2MaysT2Wzm1Rw33tB7ybknskSGtMbkb+YKpQyTZHa1HchpZkJZNASIqn8ORvNUgZ7S
iME4ODk/c8wqMTCLuB2eEZfBf4/QQHZEbi8Bew6ImPJ8ebwYgmbbrzL3h5bF0ZJE7HxM7AG0ryOp
zWUjrmQHCgEkGXnxfRh/TUnAL8An6oyXLaLWuZTkc6/Je3hu+dwME5bGpX1Bj+M0OiFhWT1qc24Z
Ry9imwpUA1wYcDz1HhBH7u807nayeZuCzKhkwTzpRUEy5LnY/+J5hwvEno0Gh/LKvdgNfIRf49z/
LUymZ7z5fm6+2XnP4kMAaIZIGoeLWhd3HzqQSCDRkiI4z1MpLfO+Rg7CnpGDgMXNMN3hGxPYnUkl
m+ot/BhJC7kdtuI2mU2mNDJQXqZLYfztlOiQeGWxNI1gOOSmBZmq1GxHnISn2eamQte38YFEdTCm
CSULIVNXgNnqb3CH1cXQV/udSOhmUoxzhNTjTlA0AGBlGPBcO9BQu7eV4TUJhbhz869RZ4I6pDhM
wrWoyWDHiKYIYTWJfPPkt68dpC1mgKeM0+CnwfdrLmxwRHPkJNvXVKBx2pT8PMXyv3SYdaUomKcO
tmb5Ry7j4apuy9xMKtDdDAdyX7z3/Jd5CwTQEXR6fe2Xc3xabWGnML/1KG8aVkyBcUfTlF8mlB+k
lWbet2+QO1bjEQ65ZgawXbwhMh4WlsjlwQuWmUKarcOVwo3ZtkLHbsFeQYbV4sBe8WzAUz+D/8vM
MpDQc1nywxCX0WDif+y5n7NMYF6qSHEiE4i67gal9u6aogMblV0IRbIKBCfqBPzQ2pDMWMe7tDLI
v9qYAOSGGJye8iNPtyJYwABti+0ML1Nz/l0vcYyhVFMAPAvjkS6Hj/9XMY6j/olUEeY3MCixVWP3
s2ouY6dd9hQLlKA5TZ+470vOG2yo3KNi/DmRFvC4trwdAm+A6eNQZJcE0t2FD4+fxEbTlbv7EoGG
jSKgBruoeuvyIc2Slvx/RiPMdlzbEuyisvZUufl09gPGF5YecxQu5WK6MBIonbg/zDIWGtBkEOwV
9R7sbDcdlaiRtruDH3ihYnvBpzQF8KW7bguZJHLnP0JXDYI5kwN/yROAJv5d/ND+shbOAPvMUz6D
bzrg2WcQEH+UhoaIi4Q1Kmt4ooWTCqVl4K/Co4nzjFVgxc/rryZ44pvFhSQWkB6Z+2c3EoO9ZUZa
Ecpy6xbeQxxWuPR2fdoQMoE0syZwSliKuWHmNaxFMXvPZzSl708690593ezkVECNWetc2pO0kKRd
Ae4kggqP7PewpvyIgEBWMkkqBziqKxgPA+MQ8WRF25OVQI2R0JvN9PdVtacFlmbfpxNj/yQWXTUl
lFrBiSPaxxZtYQ1vXBzGjfoIPbu7IoiV05X9PaIoZCJjubLAZ4Sd0JKSP9nqwIxrNsoCSFze8IpJ
pYG11e2dSvBDEerjBDY5VUk8ik7fCX6NVFR8dDZyqxilVjzt3O0UEjqn9sqj7CsYAPlssSAmC9GE
3zd4NOopOie5yRiVqacg7tL0VfNqtjtvecTqKdIz5t0mPGVSYGFmrVD1fCiwyAyJD9HqEbVjgKmC
2f2rrr0KQvC9OyJFv6kSzYO37DUNf6/r/q4AkVWjFhNQ2Fyu5cka+pdb2+V9BpJmWcmhEimiyDFm
vfMBy85zRbpxzd4A9EWb+EuNYLcBTdJogQNYA4L3EOV+s8/boykttQ9dtgR1b+Dr0/flmq+IxMJg
YdS23Bk7zyEaVm4n7zcn5cgOEvXsEgoLLdlk3JdPOrxUFxfi07FfWCqDbmrpQWbRAlMWV+Yn+bEj
G72QNSad2IyKYEuUNINFEvoEos0htGvZeM6/Buh8SboJqsnFgh9XTcIepRF+UBvMQmzxE7yIxpje
O7QNnv9FjG0ChVkUmn6M6qXtORCfMU1DzjECD3uA545c3TVJd7OZ1CcUTXsVXsUcISzZGaS0eCui
IkWw05iDbb1B4NXrkUaACBNboOoDqcGGopsY0/u5kJIYvSSiBtOHW2CEQvYtZ/GrnEDNtgDa6RIH
rb8AL05/tIV4Om7ScT4l/Ajk7Un18Pk91M93+VwekCgSiiJu40p5Ggg6P0efPlqjJhPKCch6Adgl
mpfqWID1zjWgnSyWnRbtOLpUMXYEiAzDDdyhsPgOSMJn0NbEI5pGLOv8MBDRwsDRZtQFxyMpIlOY
2DtVu9JyDidGhUGoS+ZpOXnG7T0BSbISd8qKJLsO0IlVAxrvbeGJ48MQubVTOa7ywL2Cx+MZcD21
QcXckZSUx2r85nQGo6v25mZKiZ6WFFJOHnQ+NKQ3lSUEX/xkeJfpGIsOaRNtJ61eNe8/PTRtTS9z
ts/ak80ln8uXVGpvH57fz8Rr/HY83w7f/VXZBlLzKme+3thQCCmrqVcp670nQ4qTbKWJrzwzIJof
BVHLytOJdHwwt9OoKhLMcizHnjuokiP4880V3fmkkRT3qM3XxQP+DhTgX4mt7eeTCel1JtPvhHdo
L+wfY5ud/nEdm1CzziB9xgfzrNqSZodlgOnEHQFLKTY5h/QA+gg7Xmft9cw5J9rRFa6q/m7xOkYu
oxu4Ak9Oz2ZZLwM5WRRGPDlD6jEnGZtL0EcOT6KyhiEGhxWFZwfja6G0MdSZjPcFZgNdxhNL8Fdj
eNggT9iaA+mxPPGk7Nbm4GanPxVeV93Ebx8fy/q+ngMaoS4OXU0LdRaUxGyAaPq+CaeLQZcFj0NY
nd2TyOBeGNMIUopL7DLDecuBhSX6c3tKo29KaIaopgPUsPSWbewNJmrMkBF2CNiTQRTvMEqCNY1Q
Irx6hnGxHzNH45hJdlVVnbNjYcr7bls+WbtEdolJck+99G9AuPCM8fX6BJR3QBMO7miWvVsGz4Vl
9O1AM3kDmJ92IY4ID9vKnrpvWdhPBjTwRzX9D72ep0R5OzE8y8X3LvN5KnKJvIrCeYzE6hWGoviF
XZ7RYd/1SUk8e4jRH+6mjMZVZSF0po9bHMmTL74e8CTJDsh2yxoyPGB3888oFRWmlz8FETSHYTst
3M8Dzf2c6hrohnTUeBGx5Q+xjtCOceVUFGY3yDWgnuz1tFZjru9ZKsSkErsVkcrjrWbxyPbAfWSC
DRnr5jEi3+cP9kHo3sJ5TpeXOQ7tm1JRNTRGyhhFB4pxv1XsmU4EXqBWBXEHhEoqdPlhBktho/YB
t+KHNAtNIGXblUi1X5R6GXgWJHnM+JPx93+mG/gq7RjdaLrUNUN5njRWfNWzSItrL2aFoamyv2pt
AWuRh8kPGehBsvAbEwfSBRJX+PYjYlK7XoLm8rEacCdX8qDwqqzIewcO6+r/Cj7NJpz+n6I2fpzp
y6D37+8ecFojzD1w2Sm0K+OdkgWBRk4lZRzdNtpb34WJ3jtstNs2MzM+pLf9mRoFdtow7XN0JFa1
vGc+VK2u5MV5t9mcw3HnCEop0Ohuvmr2ONpVsFW4EkouTVYEUdpFA472l1Z3qoRGywv5LcQ+ZDo5
gtNBrmAEdKuz/tDyFJ0WED/WW3wGWCAsGMYwsobSJ4xNuJcYJLa19XNscb9YxoM1LxYcrcpJOiVe
CXejoMbBpRll6ffRHxln/4goor6cWnLRHjtXyFBMkkiLhrRTkjerwu7lb+k56ZRJ0ajSU4wCDHVP
jKbxWGhQxBo0KgjGFUKb5SVyjI2YcGx8LlQYBH9MtM7py6DWSpomgJnr9SNi7w0nomq4s+nYOHbN
3bnV66OdZtHA4of/clto2xDc2+WooJFg2Ydqkg3bsE4w80caLxdpMLUSR8t8LQT3u5G/0lWxpHYk
9s8tbilVoNHH6sGHf9UJwJaDqHcoLG6NesaB4FcrV9BW7nqdSjn7AdCCazLz2sAlfAyLcHueh7zc
ePnY6TgQ1bAcPsuyX9kpVqExx9EAWT+2Qkz62G+Ng/fyUxjNg6GCi2kgol9yWATaQNsalWnixVOJ
7bO905P19Il8JcjyaoE4C8U0vqAIWwQZ1TLfQaKtXRrwpqiccm6IVTP08WTNYjy4GJMIKag9bWBC
1qV0hfixfjdR/Weei7Uz2QwTsOcXRDlr0lNqxl74q5pV4yuGvqpQmj1bIEa+22NAKRbPUjsHJ8t5
qhQRMiS3EgC9mUEUp6S6AZUCAGqY09VjnDB5wvGF90Ho6Up/vBoF8PU2iSXQWuDb6NekyJkT3e3B
Ex2S5O073Vh000bGNW33UuCAr8WwYQtJpfCwaAaB6gmhMtw344ZG3cDgZin+6oVipD8IV0OFvRpW
oPHsVRhjulQO/3vKc1GF4QnQwiIgxPWgEgkr1tu3s419eRbzAA7zN/pmDVk0xHD7Zrfssv+34ckd
8TfrirVF7418iMVMm5t1TWvpKv8tacq8zYOQTVNIEP2VPBBJCkIpFyFqsziUDx/XukTomNbaZe5x
9LazdJM7Mf5Kvju+hiHrii6aByZ5bLMfCM1z9wcSKKap6TO3oML+g+PJ1OGGVqmSDsjZ6k3+Yk0k
6P6Mui335OzN9BJ2t6WxnxVogVrW5O9JC8Eb9yxmtrOQjEdmMNCEABWwdXy3q9gTcAuyquz8mGV2
k6JtrYut+sXRdqK5vpIx8yIUEL+4xampvniiurB58VZlC7NKDT7iBxoVXHG89PLJxGodY7uCaw7w
hXnAWzVoEVv92pfO+mBs6tQkWJklo2FDh6PolEJnLmvSUVu2+0duaIYjNt285Qnzqol6L6Zv867l
QEJSSvJnqzGmP4vuXEAY8Thgj1V56+g4EguztwI0UNtJvte8lkLFYCae8qReZcjuVKHxXVhjoAsq
9G0yzgTVW+EIVKx9mjYqApCh1hrQ+CDCJkO9GBSllOpL+oV08ABdl24of0UpZgAoPbRVZqfDzS2H
gDgiplwpyGATFPJ9pAq1RDIF3BvaadptqlmpSsChiBTu01I4nld+VynBhXaoCmFuAKuKHw5rF0UK
fGX25J3RU3eaBQpmqbFqAt+JbvovNoeuwFD8axyFBriPLhVVrdXFa/+noFVvrBTdnpH01lopr8O5
BF33d86HSHczzVe926/anZ/c3wRHw7e5K5Xlg4k0H4SYpPh4cd0T4+jrUMKZqFXoQ1AZMJvkHTcw
1WjqF4KbtZw/AUqycO+uHogdASH21NGPyDom21E4sUTLpIzEK8KV3ss9JlMcfPsIRJ7suXglKFPR
uTD5SfqM0icrMjt+JrEb3lI2c48lf34n2RLaJj1l2JR5oTFEkEeWJqupZ9ZAYe7+LPq15Ypddnab
EyeArVxW7cVU4IfJuiB1Kjhbqbs30ZdSF5MhsCwlpfA38CX+l03TFkMDnyk+ojcvQfNTB6hgGyP8
Qbm3Zbv0GkTkoCVpL2lyVrmw8GRW4IzkgxaaXafQNeoLJmvdCSItrggg15oGBUJbA+vCs4mgjfkj
dcQfKANkzC8V0bedFx+EAeJ3MdPeWgwloun3R8R7Ffb91D+n1eAdEh4fOXBKE8DsOF9esdoJH+y/
FUbGB+juiu1thHycjW7AbPVc6IN9j3mbU0pe6vfStPHEjaxFtiQL0BtkciPWzmBu1FN+EKJI0bYg
//Logc6xuqqBElSbMAgtSUTzIsOhU/ZpTh4bUnBlP+onYKfkk49ZpOY0XB8XItRSXWI1kgRGTMUi
SAj3G3I3ykZpAjDMlNM9h08il5IaMIrD1uWpOpzYNZ/GYzdyyG3Z7jaia5hBJrTC+eXyWX9GRkHz
u9gPclqn238tNP+CQg7KgTHZAeFkUiFPDSauzIb2Q2Q44FpsJzRKH7pJZ/l5rSeWLRksE0n3o5nW
8RlgEY3yz/nICnsiOyOEEiuUPhu5W/iPGzHpvt1KLtf3DuXoIAE3k+jP8m6R24zwWRqMF5nanqfU
rMIXAkaYO/+GlssVtNt6rfPBPrNluqzEecAz11rZYce5G5IXfxVZ6vhbDmhPhn25HqcnFQ2V55UF
+oImN46iR6RMAIrbBbFn8Dx3QaXBq99WOavb6ifXgEW1mLX4ht+kW6Z6Bc8H12wa3FQJcZ2j0p4W
48MhSBBdhEm1eijb6KIUok4/z8EdjWtXaZiNJOcCdrdL5FGdHu68VVs1bih7EAjR/8W0IZ+aMj+I
YWhZRcXno2/3W4OpClvTgD2hRpYt5VKeC8JitaegQqDSEMA+9BNFivIIC7ZVnNAQa/MVd9PeVHmt
O7tZlB2EMoTwsOwQ9fDHaV8i0H1YdwqG8PzKVFLZuToBzGt+ahKek1S6lkQmY15/+cIGDj7hhX6Y
t9nlnn6np65HkWhuW80u6OiTyy2F05r01flimXI5iJx6Lqa+Ww3JfINzh3CrJLhaE5tpEWbc2MmV
S/CaPFvRMDKukOTMTV4MPipak8VvCd+ml71iqkZurAUmz4DgAEQT8CyxtxnVGdGKTL+eRJtemsCQ
dIin+dWV0MfCx6ezitX0L9ihzQsM9cvkMh+YRRqFqw8tpqJPxnyxruCPlBVZFqQqTsrPuXK6AAoy
3ECncuhxGlfZ3408P8hgcL5HHGNtmxxPtUrTpFNEdX1B24vzjcTUhQzb7hjqhLocGRuHtlohY2nP
DXyLOk7IxDfE4oYRT8jh3d5x+40HYmzwoYYTK88tmRJJ/TfVS9qn1Tz9omnS77NwLvdhglg/jGqc
Tc6Ub4SMllikAq1mXRshFzQp3FaJqs53q2TIgLLSGZM+EAqDz8iertizJEAJ1LimbGgiDSCiRa0E
2gv3ikqM2DHoidO+pKVxNQpM748li5WUoKHzdRmi2EgY+mczJ69MDYmaBGmw/lre7uaWr8XFBEBL
gw38gZeiWPZMQbjzcv6FqujdWc73pDsIaBn9nFilct8FOoFnKHqGG/Jnhei2iEKMjirneoj8WvJ6
2Wc4RZtshU4rfuthuMPNlYiysuM2P7tTZT3zKNPMsu0P+/D6SAQ14vhNnA/g8Br9024H7wtu/ITV
QaALl5aIX0CKcer+shtc3l982K8/gEZ3sV3QzTGwUa+d2S8hyIQmZ8viw5kNkfTH51AD7PaswzcP
kz6YTK2Zqq6iP+j91Il/pzOO0lMgUkiBjvC0RCRNzafjsHxXrq7wDP3h+CroN2eTRe5WkL62qIdk
CKHrahk7nz0fRyhF9/W/mwiIIlRxEO/WbJmhYKCQ6mQgZ7UGPxpDo9qhHCs1mDbVzv9yNZ4BicFh
nC7GzqSNXZVLMnJ4ktr/OlKRwnlwzpCuZo43yh1YiTUu16pKeuj/rvgJbabo8cUxKW8Suqzs2jV/
JJBpOtZbB1UVkSJqwrsEFJjhWQC3sBDE/gjzJUAAt8RSgVw9P0CHUOYbiPTbyjYOlrZRYukXB88W
tB2mfC0YfPPqtWzI2fIcmlwfVvtZxuZgmCV8aa5nQKj4Q9O52cRrya0st5sJzFue7xNNbzgHgQVR
zOia4dr1biSSOrdNsvsc4v1cXL/G8LccyWTvQZGlBlpYoJoeO3Fvw4qiC4AFrP2diUiMwAEqrW2n
IjZBSLlBdVkhS0WhsakYFHOTQLHrCb9AxpHxkxqyvxjgQnol4XW0gd7mwih+AnNOO06paoExvZkJ
gmWOWSTqoF1evhrUcgI8ntNQ8t7ZwkcSrwBvWL7eMtTg9LYp7ia4MFfM9iExoZbpHx7tXhtia1cJ
fmdlvH/ld6sZEVqEqE1x5lYjVIUK+9+xFwGcgRL3ISPUGMSoXro3KK7Osg0Os5TVAZKeYYpRsQuh
I4Dedabu5UVVr6d5XmhysRqzBNnWCOacujS/h8rupsDTfaMQoW66kQ1Z/24yHsINovfQQ9Yb8MQG
23dNBnsdNMzRR1I7Idg7G4gd501TpS1hoY9qapRW9Xbf3D6AwR5AmhbiZmvAKB3qhy40fIZJ8fze
JJwNXoVen7xyI4w7ygRopXlC4qIHKDfHsQ9bhJJDWMxTeep51BrPK1FZffAyjjFXxwam0WxE9R+X
R0jgHdsgH9sxU/1ZblSmxpUO7m46CT4LnB87lK+OxgLSuhJRg2f+OJUdl90EhA3TU1KXAYgaulXa
BYVBQBfYYUuecui9+IwIM7iN5qRrINab79xxeL8KYX6ExOfkq9IJKRAnkXwqDddNwx9x89O5bJ2s
jnpNRHl4uK4fRac/1EXNDKEglQjiyAe3CfcYX/Ywiqowukp1D8zv5SawCtIKKrbgpMUES6UuegYN
jRo7OLVokpMRGDjJ5MlQs/pkKTFnZfbl3ZKT3eoRCiqfZpk8A1z4OnC6mwrFbTj2JKh6YCEhq9Ff
fligXwHuh6KttZd/oeGx1RhcpUX5Q12yw/FxxFWKLbFqviTDSkfd30dtvr0SPhWZyZxLnFdevTPL
osGWPDnEGsq4HcEbS5Xzbox47OuMEN6276SzMq5T1RFc79vvOeKJsKOMjbUIBrkE+GGzeFomVdtF
vdyYpDWZuHHq4XlgUF2s7bttQ2vFa/erxn4Jcq27H9FFlIs3aAsltO3QelmQJIPWF3S3fa5fwHGq
0Tz03yoTNhubJuqqF30byNtiHvVoAVCOH1TMMGwnpPgscVSol2Lv6d2+ca4/dh4GcFo120nAU+0Q
ieitNxT3v4hLNyfjL+aXU4wvRMY1tVdWxxWxQ11g5S59zVtEA7ZUtQVLtJaq12D9tNit2Yt0esqj
4fWLHqne7LYzt9WuWL9SfC5ULleCWoLi5TzULHDaAeq9tUGGQrmVo43JDLo16AMu5cAVHFja4oqF
Z0yRdbvnDcZvjs33lYF/zfpn+BXJRDNIiPDk+TuU69AqR52lXxaLQQnJHlcteAHAYFGwuXR7VJNM
2pFZ9qpDh2EwM4q55OCgCtuT3poEcy14/IICx3OGvMnv5hUq5dV4UG0t5ua3wqLHVCGBPmXtK74P
l2hHMKpm7GH1mLU51cgeWXnBnwnH9a2+ogoOc8i1VnFD8hYomo2r7EF/C2XIr09gSO8K2j8lfpr8
Z9xaz0mnAy1j0ul7HQt6HVX80reK11DU6VekoPHyUBGehYo05pBO2ADylpsiWYP7darWEW3qWOaZ
FMDoGYcj3QkgKQenr5nHqfoI5u74DIa6pgOKjSx4jYbMX+7QsCOuRoVXLyaJiJlsKG1VQl8EfVRo
3cw42gpUFumpU2FVYB8pVG+qPKxXKNabBou0tLVPqY4HoTWkdEkRBxeW0AHsHGY4V2MMtsStCjpK
UNotz56qFY1EKHVzRVrr8Mo/PDKSmAUrhp18HwsMen2z3WtdskGgqS7zh+NvJ+N8i4u1cheJtxAZ
4NbvB5PPFdvaI9tPa5jvCFC1DxumK52BZ9FZ9A22p2b27gV+6srfV7cKxY1lKfPzHxWMYqhAnaqh
DuSetPSMcurkMVrgTt6CQXBAUY+2wRukNmPGXmL/wiISnuSXE6RynZZgThE4lQnxJbYf32DfcaQM
aZKuqKExRHHjg5YG83NgyDIkJKgmtAGezOQhFXeJJ/K+mgi0bxDZB0O+bc98x3Xw/cVEjrAY4Pmz
aC8n29vqls+9HSPkWH90Z9RkOU9tG4Wlic8/uKXXU2SnyNXR30rTUzXz34VWgwzAcWQsIsr4zbkI
rSxW7BGak4M3NLRdbwyGjMAJkG3CtNNiMD+nFlOj/P55K1AJ6XiBeU1MrKnkzjBRdw5Hi0hxXrFY
9VQRNOejCj7ydEeXRHXgkaMi+qWFNZELH2sHjAfZISgdH4Dj9qYB62yYkb76EpiY3gvLhFePurAD
Mm41bVf+KOO1hDBxcY/XprYRbpRwTDnJOeP7nzs1BBA2irvsimwpqayvU24KCb+EXGrbdeOESg+6
2ktS7OETyve2Gvbm4Io0fg93VEBCyBsXw5by+LeNFU4vGBLcX6i1ErDHUyxQzcSkaUNmqELaQoWQ
GdWhPDBzQvq8CmZCgpzgtUOSEs5eu7zlIsPCoSntEAzmGuUjCPQ5k9VIJznf+IZNAifPuXO6lKMA
Py1QA5UK267fKWbfFGQW0Yctcp+89gNxuNyQLmBSOIMUgOapapsmRKjyiZTNhfRbhE+dokerMLjU
CoxMx7weJOZvrRdH/bp12WkeMaHClnDZotJxB5K2IJ9KBb2APlv6wuYXdVTcGezc+ysEe5bRBGm/
jDeZlyaSm8iZ2PMp2qzeKSuDLoABn9HWv0mwGN3ECZB7csLNH6k9tuljZfYluxLueAexK2Th+La2
LK2a8Y6ydbizu1rRAc0/xoDsF8GdvPjFUI7xO7W3+JLYLy45RW90ZvW8kUuTIyxo18TqKzlXME5c
NcyAswuff0UHpKhVO65KW+tHZ6AEETUNG9zrKUn3B/tia2sckidZHOdNeRvRXk+OsqKAuIuOuUY9
WQaUwuSpLzXE7rMhOIKyM4Ay4DJP/HuucGU8iG1bhg2JFq9zLrz8VBzBHcgFD3Yz9pv/TTe42Ymz
pRWnQqHAyhweuj3LZ/ldP8zC8+CRXXIaKlsodVPclWl+XsDsncEzxvaQN5QX0j6zYwuyR1JWwKAa
7nQxSP0vn0/SsOr012ERZkGlK6Pp9Gixr4+FRzyRBaJiJfvr5Ck+MQ+uvkKT6uEK+y7nmDHh0Kxc
LpCRxcTgWI2a9pujO5ppGWUnkzWPilJ//YZr8Jncb5ahNNMT9ya+RQIAZOXYK5HTkH/h4wmbwggK
VznstDWbK3PMnqo5KjOxzvnsMbctX0u4AimYW7U/y9VLciL/W6GIAs/TANceAr/UijpvRpXczfRU
zp+grbRgZ7afvFDc2TXhaW/zREStW/9EvUzECpGPtsBeAj69doIYayyRTygRmeslOVPJFqwdjTA5
/Jkjom6wdB9neSqqTMJzbgi3ZzP9awgFTy/A3ravMVkKT45KyZ7p0oQyVq4+Qb0FuKMmI2K3Jkdk
OoiKVQcZ6xLHNk/FCXREfd7GfNYeNhPMfrjhTMLzRCT1GvXXpilJ6kLGyYGDc3FHhtKlJZaL4Cf4
208LYqb80kMJ2iofq1ivhSgPEsVMemP/qE6rDQf2+70GcYR0xI1rY6feQI0iitItakr7on9xvhW9
2VLFyLlYJjpCm1E2Q5mLTr2pe/RAGogSmXu8y4EvTVglZ9Ht5OcjzagRMfEYB8m9S2CXZamRswI1
cAyMYsBPFYqUPhpUhhyzrYlTYlI7iAg/DfGMFUkEN6X3waEWYPn4yY7KqFM3OUZp8S5+nQuMswdO
o3mgsq1KCOo53UFSXqB8hWESDrJbW0G3uHKPJrkaO6HMF13i5qjxIX7Q8XnY05zKOmEixp0raos3
b3uUcX4vAngnp5wPioPT28y4hh/kjj/FzlNW57pRuZLcNDIO34439Fl7IVhF/naubk0HUg2qVPTQ
yn3p8l5b2v6y2iCu2jH//JZ6FIJIeb6yoTwzV9SFM+88E1L8ONuxXDzyQT4tYK2uL0cpwaTGpMc5
Cl1q5ZBzMoeQXGGL76tOFk7J+ziVDacLVR22e5xhXAgek+/Bis+1VFxOVvLZ9AUBCTDqhffm7XXW
SvBe3j1uvG6YuBvmRXFc8R3vQWP9dx2SvV4BftTroOYNBB3jdCKKjkIy/SpN51JoPwfEwoWJI0sc
iAFLiraGAb/diMtzxVQ6HSoWAguFratlsW8Hs4eTF0dnNwSYSQ0uB/lYYpW/ZE7buTg9Djyl2sC4
+0wGMfI8L48ZT4Q/d0/OR+Y7/WKqVkGJ1EgKwFagDaNYNwNaph1JDfiLA294vQJF+kqAFOkY08TU
9f6bjfBV4HD/lpgsCGRKcglHzbq6egsqtMA/K2kEDEerGGviLMb2vhCkpzQ2qDBZQlMPMDoFl4a+
uUbhqaNcdIakxt/FDnwPxwSiTmLx8mY587S20nPor1bcwAtdx/8Nl3r6pzMhNXWHczizwSRvbcRI
bamtplD/gaMQYu2S2oyQycAY3OEemj4cl2V2uvCrEORSzFQYUoxF9Jr7h5ynX3d9GWZTckXuaLfI
LdZJntJTr0PJL9LKaDw6EEuH+LM4N5ZRekO+ewulbkvbv0z/DU6zDUPgSpK19AwvZb2GVzLfpIij
tohK5Zg0tbExJLSGpyfu8Kfv09y/b4l+CQ3t3bYMrje1bU8YYQYGQBjzJ8cfaHzJyGNHXPcT0m4b
zU9NnzY4boFshMvGJydZeTQSBtdeXKa6Aez9uQfjwNBffkOe9TaVI9i96Idbkf8nhFmE2m/+iqu0
CVniqoeFg2Jbf9hYkfmwWza6RACplnM0pCtkEICyy+7/MjOwoMY1Ilo8ncfV1NmspvqenfKJVZhZ
9ffRC447eIPenBTmL9edCgFAU7zPeBdXBtH36TT8OMbNjQ7G8K+XpdhAwIp1p0LVybsuw05HjnOL
ym87o+Dl+jgAU5YN3EW1GFDFquayWXv/OZ5+Kuln3VpDW8pxmTuT+1hnB5to42FYT4A6uelVuz2Q
AsAgQy8TGIMv18scshnmVHI2k2ByONV6L+w6tng9bB19epA8Jn4fpf+gp7LlJGHMiM4cXznJ8Yjh
BKbbp2gWYhbP6+j91wz+A4YambN0rttSLYSHGg900RJ5//cyiyz3b7Yyt7DEF0uGDZGkeiw/XSmv
YLJYfjKq/aQWddVwpQ/5q4Pa+S/KZ8ktf5SXYE33IHxzApSPWqO7MWieXb9xT3VyxW7epGB9waqQ
CZuZbOhysog/qhJi2n2ixG3MNr4mJcfB/ZfTXg8FhegFa12afZpkGldjsLTnpZTRI3e0fITV1QkQ
ay0e5EE+jR7E5fMRFoyiTAnV+rIIkVhs39ANS/w+RXws2DGNyQMYp4WcC/KFFH76ahdOqOzP7Gnd
xKAfXnJN01a5bP1gIdjv3fKui8ApjWPUv/F/PoxIf+sNGx+dY7VzdQnJXFtUAi2x/C41cDjfGu7P
kTapJoCT9isFCYDFOwH+R8nZobErMEShPPbVfPl6d3X4Q6Sanqw2K+n7ZE+TjIp3betH3ar5zSRH
zoUk/cMt3UVtMUSe8+FWnrd80yqMLKjs20O845M9aEEiG03XUHmgHMXkLyYt/g0sDLUWrB9ueZhu
yJ9+XPhgxeIXLvLQuz0jzO+C0H7RJT3o+n+aAlGD/BDb5IWjtHEzD35tXcXTORSsBu2bNVCtM2eB
H9dxdaCvDxc5D0Sa+FH/vM5cqco8/rtS50RItjjuh5wS8sRoLW5x3BrWQzofF5R/niVze6WYiWIA
VByRt9d59Zczoi5rwkyAUygCxWzxPHBoGQDUFOLTIrSiznfTBBvghczyi08wvNptX3CvHPBgUyw5
meDYspI2YKwNe5Z4p2JJHSXrK6w65dvxeadR6z4gungEs//pJMDBZHBdiv0wBVYV8zzDTGIP7IQn
EAnCzEHWUWIT/d0wKictFddWYItp4ZUOCnD0mZY/1VBmq+Wgl82Iz4/Xy5K54kKDJEb20XbyU5N7
33qAAmGUpK4RZ0+iySKihb/hMvV7N5pdqGVcLndoi/CvZpU6FznqBZNdN46L/ZzgMd6A1/7aiBcW
JraFxd517Gblw8nJux/R3gedt33hTZZJdArdv+5WFp37XZ/S10s9m61Mx+hhZ9cG02ze8awJH7Vv
HCF/UXu9SGD4oGJMxqQJaWCXf5Zxc7yDhnyYPNeTIgCw+g6N3TyHpXUTRL3lzLkVEMGUjnwB/pnn
Eic46EunhjkJKY41CByiJESE/JZ19/BIi1CrflMkYkUXvz9fa0lDooO8ovmp9Tguqi8wpAeGj7P3
czr9z1f79uiVAPccYoemGA7STpTkzrD+RndZo8O3ooauOlZQmW6SqrVbCJ5P/NJVZopPmnZ5hl1H
i63t4V7lBwvZ1U4ZOILqlawjijfYT+bqiu8wFQYDVRg7TbMAV0ZsbA+bvIoR0ctcDUdiOB68RLzx
AsOurWF9Zq7vK1vpyTfWz+PdsYHEKJ2OzoF9yGbOMiFbIQ3IVPVU/lsoEOQezODlk6Eys/jkyBHq
PcLAWdIeNczBxtMgzAnZk0N+54dZq9khDdo9bkzNaS9HFBZqvhJAj7WsJjw0ZlCfQZRdXdq8eWeY
QeYs7G13ZlZNjsXgTG6qBYUqBgwERXuPE4YuqkWZ2WH1v9MuMD2jM/e50kExZrPC3ihGXFeVDUvW
2UlszmRInVcrIrDBuckOvMY8lXVsbIrwnU7Q/yDKLw2YUD9ek/PGzgyHUvxnZezmW5VCL0s/xsYa
r2YCWvh7JlQoddXThzWMuqr8MzbxnXWwGr7rj9G9IdLfGqY+P8+oqKDnHY7P5Dp95+DmRWEWTKrZ
CFbumQ7YKnf3pWhByK1LplKG3n2qvrgmU3FU84aIFbbgwryERKb5wDrmJsN54gsb9tB+E3Ge3A5d
yjyvUjQrx+l0mQzB9cKdM7OPPSrUnumyKMqjKfJbxgr7oACBDJdsP0XjOqNK8oSolCxWHnyTg8Xi
t2GhGFCk8DtWXk/w8Y2VT7UAcjgII1N2iDJTpduhXFGbw4cklY+tgKtWItOkFbyVm6yjKFzDzYjw
peYqROXDVuh1Ii5JJNzWLaoL3glvAaY8ZV5azuY+z9f4GWhvplzMl+OY+czNMdS19oMepyX6u4nS
1aJp9NTB9ETFdGI5WDcRSe+t5E7AIDXXVpO2isfpvOXDzBJLJKsxqjIy0FXp2b4OTkgSDsr91zoF
TyuGStbpokICz00njXhCy5EJyoXwztrD9WLC5rJFH3CUCYTf4nl/lC0GJR+8r2cR9HBxE81fwwRJ
shDdQ2Tgc+0FugGytg9v9JTPdMpcxWYVwEORr9GLjqiVEfw3JNkTIViJ98wfqAtMr0Txq1W10b5M
gnS4dzOLt+t7e45v8J9zQURb7/toQJkZRSCP7I2ovfbQxZNY4FzQCuPH9AHpuwGgIAOX77jN/EoC
NmX+brnkUDFbkZfKEyCXih9gULWheCMd9pOAoynoVaXMKmsvznLIPM3v4OR4bsT5mmKuo2RNqKRx
Ar+54zDG4wR+any2EmTTnM1u+x/hikhanHjaYVhNI7l0yo343ohxDa9qnm6RdrZn8ZW/wFWvNHcW
CmgQ7KjwNv13dLq/OjUG1zC/Nnk6eFYm/oVpJGtlCnB/Ur73bJFHBbgS724qRsKldobS1RgdQSkN
n+aeXKOXXUx/Mo9N03aghBkQuzBTiPF1gadAmRckfTxR4Z2yAgupZAjqZuzWgtV/XKegk0m+Ynp4
F32dXp+lRG4UEJ262nJftqLmLRBtBnaM3G4ylrH05uMQq0/XnYVECu5uMb4lGY7sDdG/7EFK9cuc
lg7zH2EYDYL2foWYHX3Dx4ltw0M+2Jny8gMLI2N4LPv84VT8aOdCIvJ3+2eeSHYXpXdyEM0ouMsG
6VLaC1rFcQCJm3AcKbmzezT1vCXgEMOm0/M1jav03CWRjn234IgJAwH2yJJ2voCK+r6dZfnePSof
GuXZNsC7hyByVBfaZ1EagwU00nANKoA0lS3Tt/ckYT5hZapYATbhzOAes2UHGqvZFgNTweNhb4ul
ggVtxexVECtn7cF3qD/6zzTSWbUN6AJu1Dh1ZCL3ijdaW5tQkIrdBdf2cJ2cz6nb10Ys0FK+N6OL
FD72KVU0OOp9ndAfX/OPoVXjYP9dTWdjOFW9uzgzKgryaCN9d7A7Y3Lgtf/UqvhjaYmXINbJf5Tt
L9RZgzA5buZRhfv/QZqTgAZ5OR3SAOgcLApGhcK4z+MmvqSgx888HBQtLlLMl2xljD8OYCulpeCv
sRKw1FH0CM6OA5VIMYwZkxrvYDmZIIDSCdFQZ6Lx2zdjgBanQvbZD/EMCqVUZCdqib8snk43eh89
agfqvzFdInYc7VEMaqGvAMPrNM0XqNqTUr21YDCx4TXWOt0Xahbs9CAVQZVSc6kdyrkDmJePrWHE
+ho64nYhidm0BlVFnXVbJPbXjxjx7xqkdZA1pu0dMM6x8PUm87pRkbr4nY262g3DAPyKlCkIuDU5
xpxB0+rrTs7MzjImlxdX/Arp5mvMvWRXWZpTuIKLJ7KzJ3aVyrdt7uN/JUtc3DELnPpGV1zi9B7W
S/wRU/3E/8gaieANuYDuZ78Jdq6GDFICIg2+kTGW5lasX8DrNjru8TmwszWVCGPIv/YCeMbbT9N1
SXRUdNgccuFBxGS4EPhM1pmcYSUl2+5+qiWRdkihyJ06m6YbByG5SNyn35L7nWIv6zJfXK1y+NIo
UFIIifc5l8bXAzJ0inruOQ1/4LLbOTMLoKsirI2E+kmVynJaDMTUVEVEdyPC9jX6wc2F6Qotdv3P
qOVAJ1iC0DfK+XbMP3p7S5nz09/fO9StQb/P2O1XHjcJwYCFQCoQXf1wft5dyLjCVCYI92PSsMi4
O/B/CLU+fsHpF2OVTR6YFzXOVx0ITSjbl9v15Ze5HPi9rzol/XHKHHCueDSBtzRpJWYVNL4znWQa
VtdWAxCjE3pwU0mMMYzr6Za30lSyQF2fQJO5sf7l3497oXqc8fYaJIvS6IgiAmAN74CHJBgLblLl
ftqHAunfv/WqTlddhBwBqjfNX7ptjQ3mkY+1NPuIoqAoaubug5hI+E0FKRI2iZF/6uvFDGVwn8Ol
72jKfSkGgC2sFDa6fv/zUMzU1p42CWyBrD4c21DiI9asRz/feufHsTtLlJ4Bl2roG+Ye+mMI+tLK
8QLr+SeAf7xHYao75s9jM7peVoWAJrJ9XESbQpAzotxihqvZ9ZAIaw8crVXZ/gp8FIWvTjm/xHTM
Yg1teJd5y1KO+KfETTvEeKUIBOtYudxAzX5oTNGzQADOBkIX1LED05IepU+yCfNyTOsf1qI7cPZJ
95HQ+2yUYcE/wrzhoOIshaixYee4NfeCQ26+xrosAwgCTfd9CuqDzP8BzyYinoCHAc6UqiwS+/jU
1uOKo/sci18aQ232YQsRleFeUlmHGwD0fmaxnhOsX6eylDs1uJQLgHXpqEDId7ivza4+Iuk6GdY1
9Ay0SMl0TcRp7DI4/f06bMUPCQzD5rhhbmu2l3tOCsAA8p3hUV6/kaLkzFNXjmtvf6zVjk3PTS1k
Mn0Yosp/i7D/dOhKwtCIKpTOTteA0Wo4NiL28mLPtvJXNIPSA3FTkQlJBff/pyFSj/WAC+axFT5M
nteZlRvPBfjT2A1Mj0n5Ict0MM522Enbjz5nGZjLTZ1kmnOal1EfA1Uy+GqRMco4WIp8s7/x6Sx+
CLVx1HjZZ0uB+k7uraSR7RYAwZsAxBPFDGK61he4fRtL/A8JI4i2vdvvITSosC4ubB1d7Uow7yec
9zLbVbgoHhSvzh+fKrx+5y6ziReRjpvpZGIVW+CrjCW5OL39s5rCQqmYcLAw32gdlKYrpM/2oCRg
/hIbZ++7QSpJKN3tJFgmol1KHlBdkut2cJsHrywgZLG69NcRTRjq4uaXxj/Jy+eIwlozTxFz66vz
Y5r+zcQEwJxUJN3dHFE9e/IL1MVE2plu4e0oBhTWjjsLsQJFtsu5SomWdTG5IMmMEJbYrTru+yX1
90ehawl+HquuBpPsw6dH9xU2lO4q6qqUjrs9CiRB8twZdzbNgl5WKXP0q424f7lEijTRHoFELyke
l51r6BUxyXqYHiHGwC54XUjEaX9VM9rViIA5DgW1CQ4bkhe19UJ/rK03DDkpMyxHN45Y3EyYXq7m
IPMON0NsKT6o+16QufsjfZuiq4ysxsOKOBnwu/ADsc5pX9uRlb02WBCs+UZddzVSB9imm9gorwhE
qCq5y5eQ/AUALGCTqpm8PdDlSDXfTPMFa8NHrpu8WQnHBxYFJcGgjci2kf3TuK3TrQu/QjYD/ODX
coHsOBsBtYauuN61SnSyh1meWkZE3gOWjVkDlCXXLdufKtO01A7HkSt7bN0FJAUQa7POK3/M9Pzg
O17aHoUZb6bGMk2oZcXzYV7mXaSveaqSz48/DBmtGlTl9mTLRU0lv8aFmr5RIYPFo/CXOOVlAjaK
Ot1KqdzAbq6vT/G18PXbMPmsEoqSGLamPSXf5S9e2IDISob/DgBITez6OHxlD7RhEXM2E0TAs3G6
zSAevdEgs7qffXlXJ+MTJsE7cwmbHMiOmunSQ8ekGR32r4+mKhZsdVQqYR6SVXYHh5bDtPQGpu9h
gcgyNEcC6FX4Jk3XiV8eQKwc057+Pf72pFHYEv/29LZ0rg0Agw7EFUcNSns5UOaNbybWIbssmu4y
USziy/GZtb2lvuLRMxo9O58zjkGF1VegK8/nvPen7ACF4tyJbNLiwFSxCFjkEVEvpQRvIU4mMJnE
yIn7Qg2OeIZ6mw4ME0tJdb2/xgFuVUubDS767k3yUomdlob9SlWJ3dwH1PH1wSsFkORaMFNIADaI
iNojtHe/44yzvYwTdE45dKtla8mM7W4hIl78wJxNVd4xJ4Cf2hFVVvwZallzQ6xukYtd4tiyWO7E
unPh2S7XLrhZ1rb4vD/Cmqtqn4V/jNGBaGYgci6jB3yzliR6PljrsC9GK1ibSgYU6V3iP2DphIyd
g6RfaQjbZQ3vfKDRGaoRVrhbidyR3CoD5HNRZ0sx7rV4ajo0XXMTT/i/QebjP/9ZobDN+oapNEXY
oCnVXgMYf/c9C40PqrfwUxUzRVQSSQs1rFpC/ALfwZKfEBn8QM++JkHrQmvqtCU6/Wzfb3ryB0L5
n4W/r3TAkvzztrrbyWDKHQxi971V/HOIam7csBuE7n6+ICsWJ15acOMLVD0NjPgncxSgkr4Gyroa
IytQKjWyMxECYdX3azoWZrZ2E9QxGCDQimCGdNeaw3efGUN3G8hi+BK+2skU7xXKI1kAFa994U1k
aWr1Frp77M+fCkl4MSnv9CWJ6kjWH1lXv6vf656y59cGvdvhIYy0aQ4WAUL5CzySiIgdX/n54+Lv
joUD+xUZCWHMSDi1m+FZA53QhQ3ghhKIEsc3C224hQse3dPe2mY5SyUcHG/Av9PvqAnSjiS8ZzJf
iCCUz8zDjJ4lSCGPwwnnP6o4XRpwppHA3jiuMrLWblmlcSubJtXOPJ+Qqo3cEmlfjIKcDo8TM+kR
XqOzrE9hzz4ypI4EsjaHA+Q9xI/oiJdGTImZey5m3w6CGQxBoEb3BAOJH+0K4CNBzeTbcF9ubFIh
ccv2rCK6sZhGwou2/08gzqaUq8YeRCQ0BMOckOxzj6ZyvOmZIJ1Bs+ym7A3qE6xKofc0Audcfaw6
TxX4CNmNhGGkvWWsUQ3Ycci3GyoPXtXoloYEQ9zof979lQ8BkGLyrShN7Ti4gSGtJScirZBs6f8Y
qu7IcnATJ9CY38IfIzArUPTv7xS5G4wnTR3tlzI7dcA6HOj2+ty3xnrLTij+aOqBGyEdcUtggq0T
Q4jVk14j6EN82iUYO7SF7qfP66VrqJgpsYDI3SjAAqJ1squINijZQd6BylinVAdSuxGdmuX7rea/
6ACVTaKeR1xPDAXgvVR7hkA4aSzMoTrk8YM1jsrkO0LJ3uRoaC05hJAsibDFEb24hV5ZhdsQZ6q+
Nn+jeOmUukSeTilE0ekFtwm60nmjSgdSTm6+rwBILfbURcYCBapmAr86tfQ9E4oo0oQ5GiCd+gQj
imSvPrCxxnhMgrtW2pUfvy/SZS3Tj6KB86o7fLissET53zbVokzoERRLstAq7yp8Dk57dkZpucEl
1x5NCDcDvO5nhuMlz3SYqrqWtsJbwsXA9QGqaaVx1IQtkZZ2xcSaDpDs4AntDvt3u947ZaZEDode
xO2OuPgfBXurn8YXiZ98thMxNBTEa0jQn1AkSE3OjtQ+tiup1MKjfh9SrHw8oXqETjuNA5gBj//Y
9YkTJALfk3HMEYiWhtKnM35pZwT9YLsv3cJdo4W4tWRVyxri6ABG+ocYk5FNMjmhQN1RSibKbmkc
f/OGHYZ1ZAJwDuV2fqQHUM1Vih4Tw20l/KncFpXoxHp5CHUcZLTIOL+ppGGhwHONgy45wPBktRU1
OnRuF3uMKyhGxWtV55AzwFHmDybU343V8qer8UFMRjireRCiBKZM6Z6EP1rmRAr3+jypW7D4rK5K
PHTf3/cJFs4C6wEvdI44tqxvE6wak3frjvkqapcqHtKUDKL6u+FNkF069nr/350+oYMy+QQGCoS/
xlInbgYycS/ghLFaudZKWn1XxDg6muo8F/SgFZyB/y6Q+cKCJs2NeHb7hOpwMHW7Roj4me6uPFWG
1Dr4KmNB54UjJhwzOapUosTA2CLHfcHBuGZCfGSRR/D+n7mj4Ld46EXbvrqhSLqp29CVi+x6ZOju
uxMz/e/GvmyB1fnAhDK4YAA05jeWqOiad28mQWsACJfFwmDTP+dYG/M4PQP6tHGmGeSit+eAoYMv
/n0/xhI+dtnwzoNfTnPJygy5kFUqbrChAzz0BaBIcKF7CpXupGbaO2LGlLLmGMBMfeXciATTxhvz
qKJWfhRX1S0/OJ8A3fYjZk046tYRdE/TuAU31Lo9FdgCuneqfL532Dnj022QdKVV2FA0WBiQU7hF
KfA5FhWjVQJ/s7/atg+kKwF40ro+cOtsUzTvvyaf1hbaqmjGE2rZ2yditZluckBEwntWuUHgh8Rp
w+QOG6INWi7skM74hQhv09b+9aCT0/D5ytDuHqR0x0emnDZ2jGXOwXg6S5wp30/o1MUtKv26CApa
7Y7ICkr4tk/738hQJ7fROw/LSp/RlPyQA2Q8CqSLSBMTl7NvLKCVFT9XzKO3TAcs2Img4zLVZiAJ
J2ccfTMsx8Guty+TMVdj8Rts5xLZ30DAQjPMEhVP5/5DvoSX7hWnPQCUMSX2FrRKt8Nh61tb6o3p
h58YKxDDi5V84S5diDaMJsfszlMQ1iA27gmjDoWIkVUVww2kic/75FeRdGFItiHK2bihfezievZV
93JHDGDO0f2DNP9ILFCQWb7ziBxd1G0cqlqgEOk3CKPig3XjiiCR0FfBWOwNfWQY3SnI6jp+1A18
ZwHokIvPjFaTo5/no9zF46FDNw1QaO0br28snoIPahQI4GAsshAvdavClcbiC30rQX2xSnx7c+18
XbsdVSHBbBGqc7SaIP4wQGuVy1aWM7h6kHdvzsx0vW+Ap0miA0DG5PWPGMKcJP/6vhGfHI/C56WP
2GVwOMOa9MpRaUbBaJbLoQjF6X4wYHFUwonC3n3N909J+skJxEi09oEXu5BrjS7dpKTxWdvD6R62
7N83r476wZ3ZC1t2vx8TtvE5RDTUS9Mmekv5O5xofi7A9SQhtIaMNV4fVV6GRjw1SN+hEC4CChAb
F4DMonLA3Eus/vDhiSvirW/gBZHrMN3YXVVXXpcqRN7rvJfgbpWSSXMAjnm4tgVGjhl+YoKi2mJ2
LzfwV0CAkkpJsoP0GIKvo4KEszNZ/eYHDlhlZy7JKyOc+HIhkRGCu7fhDrIErE9JwDl8b+zYywE3
1ByO09WGnWz8KaBkz/zMk76Ph248aXgWnSuvMzhrPfNiUUtb0K2xEpvTAhOqpP5in/0dD1roEiRH
mV7kdCVWlAFTobM+XyhhgXfx5qkwMV2UrOzNCHf/toE5OZuDPtIB1JMqsPwi+QxVgqSl9VPTnLgW
DoQnoOPtsQMJCsbtN+GQxbyeLRSnPknWjzrEgmoFOwDJetfN9LEL2IvaNtwIDu8RbMD611ap1hbu
xXE5xKc18Aj3YDiCVzRlv6cbx24YSBObeK7PPkhgaPiiWs3rzeMb7sAvF82+a9rMQZuNZv3Rz0zF
QK7WrB8BgW5daabgr41QkPY2FW27o65A8QpWSDnAwOaYHyJLSEr8z17MweEsHnSjWXGtWlQuWgMC
L9mNqkNionj6r6th9bKoBnK8LY3PfYdCU8bLqTjcjvdwkzA1pF6OtLERr9Kiwp51U62q9yggL/nh
0+hPjBYtsRMIPC2Z63tZyCA7UuAM9mOtMz3OddV9SjMDGJxzYs5ZbvWdGle/+sSoEfFEDDV6xUtS
8vPlWtCfCw4MK/BpqHrGFLFI4uRkT9JiHPMqP7Z+Zaj1+vKmUSktNQaj6Fe28Rl5WmjXsaYQWTyA
ZVdl/GP7Fa0NYZ9WFcJWTGtVss/xzogeeoPba2pePYDwxC0Ipi1NwnBTfcP+DTXMcJmvTueeMGHq
q+NbW76VTStFsiWKEeA1bW/HEo4u1fNrLCt5IPA9I7RsMDna8HF6jcQcEDIC9MreZ0oiXUHx0qE6
ZmCFEHFOnquTmISpId/VvNBUVoe0L5zh00G7bXPF+WxGdxVoX71S6XdeFcxd6rEv9G0hVcVeixWe
wIcM4QqchBl1l8p4cA4Sba7tAuoQBW+RbPrXDRpj8Y7rK1bafV1QZwFxoHYThW8At8P+1PDGxmLs
rBbx1hVVQKSjO/rFTVQ5bhXVhNPy/wDPcubbTiy0WTgzFZQS/iJOB3oCDGyJ1F1HzCn1y5Ul0Exa
Y3o9CFlzJHMtrmpGHzDp+wr8CUDB+f0aqH43sXPCKulNLQZ7YWfhzZzJtVxPJ/vMCSuevKMJ7yDi
RNivitRQho3adBPh0xaf6VwO4SLD5dfGvH7qgt8Ue1LS+fqzhS68ht6ctL0/UehnSFQBASZ5559e
u6nfyWh+L3OyYMS5kovgXL75B2v79kbj6ovuUEEh06d5ul6k022kyOgJembU/irLJL7mhqARcgRF
GZDtPBOTeO+S1YwoUlpqlTEOFl3ShKXRaw0z5VojGcINopuZFh89fLhmRPoCCiW6Vg1kbrzkQtAh
92/na1EqOJx/xttJ2Kc1sLl05gYS99v17BWGTVmjGtNCDvgfVk51jSmukj7Po+Kau5WsY/tb8taD
JPWq1rWHMhrNzez/UCayLA0AEpxqTTU88JHnRjhXmK+tpD6KxGuD5cRKfGLKGZyMqI1pgBpTnffW
gciR6rwowy0+rOTkQ8zHV96JDfiylo9gP+kLtZd+xd7uywEtA/HpEu6bzEaSXexnAuaMhK1eSOR6
qhAUPoj3GxLO3bjMBSErvQPebw37ClwMtKqrVhpUeZpMAgUysNvKUMJBjryOJM+o4jQeTjNzRBQ5
Lj3YI4XhvWL0Exlp3PxCag4Q7e8dAIxEZF85FzppIYuxj7ZfyGs4We2Cr7tWLeO72H1XToL1yKRi
7FLx/tmXvv3H0RdsMmqnmZqvnlej04OwryGNWXMvfa5NYMzZ1m40U+QDGY8K23vD8jyHpEi/8joh
YPMO//geHaJ2b+YI4O5r2egkqKVZ2GzJlHwdU5xI1Kow60elFBAZYHFc7CGexO8Efn5+0LJMlDHL
j7RECJF5FIJS7vD+mG6pxqiJvTqPb4Gwmwsns61aw8umCn8FR2m3t3L/4jH2uxPN01H8sZmbfCdy
oGVtT5HVP3ooWiqSCklSrGdPfIaa3btyriRBsXlRuPyVCkWDlE5Ig2euHbn+ELBUxAEushlVzNrJ
HPuRAt2HwzeH6M+ep0UGLQvBflH26iP4Zm2gSRhSW8WiiW4ddfyZIRfwuHg+z6ZO7b8syjqlWMTj
u2vfYcOVVhJiLBn9wvQg6E7vqyIPEAF39zYG0qs/c228WF+0ATgfnbCx5yPiFlrvcugBqpUmWqSA
A0eY4hdZuLmgThMuGQeNA68j0Phl7XuweYd8NGaI6s2tN3OvkjykEbyG9ziRTGi6TrSMzSfP+ivX
XbbJGL5LBr9ixra3yg1gf/3RRNS/EXjJAb3Rrj9s+5pqknKhXeEdOOEru8NQ/Y4qsjhVvfVbU9yS
nDt8HlJYNOIxNSHm01uvCzM/+Z1XjsYE1vz7MbwLOpYVUNQSIm6l5pmXto+iemuoM7YbS4P8SApd
NLnPf4bJztKYerKdmr12S+92Zx1WdJuNLQREoQPLxAWp5YTzsdqYPzfSeX2mpZ088vXxtPB60QzE
uGNUtnY5+ZrNeLKs6y9fhuOxDaXpwHiaFjt0N3CPqCTY6LWliauQ2B32q7aAUfve4Xwdw5SEfh4p
q61IciMyAWo/m+xfO5p+V/RdnTxOEw1HrS35qSxm/3DbY/QSPtHU+1Rq2F2/8IRgdcnQpEOJev7K
YsSK0655hNH94IHYOGq8QmpxawbGLuLE4HVDPl03ELioYY/h/kByrSHJeEnBP3UnhegcLSlFSUKR
pz/PrpHxdinKnji1tjyGlL30uvkPOjdPHpEWpMr+UlsMIdUJP+WSkiaymexPgcQchbPmYFU9k+U8
dEjW6yB9DOfTbmY2q8FQpjYUD1PiP95aNYb+57oWsSZBnvW63gbF1bWaAclddsxs0sRIZ9IZOcnW
UIwTpQjpecLIh8jV/ogRv4H7pidfCwK/dv4w2ARmgK8ZAn2X+sZrtfWDa/Pfx2H0G3Hw9BN45Qbn
r4iZc7lIjLJMlQJ0sIC6jfsgLkKfX1q/ujeCMzxBPvmquc3kgm5D6nXUzuFQjoB0GqSbfPeQIaSN
6f6zUsfw5kDv+bU0Gzg7ItAb5VDGanW/UztnDapHNa3cTgfowyxg8qXJxeB3Nx1DmQNyvVmmdHxx
LrfEFZZwCv3lzSRaUbnPkHgMbCsfbLAZiQ5V+fKxnIuaUTTokiL4wXfOLcMMMfUN6R01kRK4OoLO
+f5tBwpp145MgEDHeLR1ZfGaPwSe5vnaCBy4r01JgFw6QIgCwIwGwnAT1ZWlInHQYwX4miY8iilx
3VmAQeL81ZtvNi9AtrdQfjrO33zbg9+Iqnw9pKMuODlIHMv/LmX1IkWW+HJ6R6aaS/pQ5lliMHbG
tjpAulUENQo5+52jSXcrUhrI3uEXbfBpw+WYQpFULwFJl50OP8/p19CU81f12MmMS60Yp7zGGMDT
GmU2IRj9Jp2n2ZMha6naMi+ly3m7HX0cZW1S6lYZ/RrTVfOVaOkNCtfnNmtV/fWGlRCnG2of56DZ
D+0H5QJO37VlXHhlj+iMFDzKtviUR6USIl8L5tqInUDlatOQnCNV4vy7EsQJCazPdymlJYf913he
2udh7MjotQ8qkrJLYZDswJE/wpnQyJsqzpoGd0w7tSzpe+J+h2P4X6V/HHO6un+fkgm/Z6MzCsWO
TQm+2PY/r3wV1mNTphlu2mQQAAWKNd+sBW7uHqHEmwb1/NXwJC51eY2SbjzmnzPik8rEDsQvUUxp
D+JMC0+ZqZQ78UvmbIyIAZRMUuLFo46cGXXZvC0JHLnUkR4t32efmHMFsB3xFyKMk6q3MGM4a2iu
6j4oQN3LRvU74TRmQUiiT5MO3DrY0HQAMS7xUdeznubnBvAJa1tnX1k70S2Y7e+s/yZ2cXlePn/+
pzenVcsxbXRvQzGeB0FsfmajGeylz7weI5T3tpHK5dQLqUuBc0RlWQtMDjW4Vo0gZnufzgkqCfbG
VEjZDuttRNWw7tcqQymkNqYiEBaT/otf3aHgqQEScKUJ9SJYARN9JxHZwMQKpIrpp3hw+8zyXN8g
hzqTmtUibQm58v9RVuF3XL9dIwvl5vhgO+JnEm/pjIKc3mGc08o3KM5TUmj7+HF7GX30ZSWWi/mL
b2K+keUaySDYn1W/tqhNSCez79lvmjKz/+a9DJQlCgHZhvopQ0EcfX/UJctMAv9fWs7yudekoYDI
SNbJZjaukJpIhW8jn3/CEy44PBlWD49wyLSt+LDTCTtjTlgJJ7ESxtJrTx/9+L4Ks9SIJa6Om1Ug
xCZGuACjm0WWa82OZdAWEut/2z8jl9UV1+dcgr67oTJ7ofVKZ+S6OGpKBeVSsB2KvjZbRn7kn8OX
oHntJ4bo5RQUpZ7CIDY3VQnhneYtFuVs3XjrL8ScooJz0KarvhBikh4NFa4hcMIILfy/pLRSLQxd
10zBYkcyoyxwrOJQSfyCQFwTueNmSZXyWbM/wyn3+riwwD1HHQcFzL4USQ5j70+LGgXH91SEEh4A
fKLVOYMiGslq6F6HV4jIrmbS3rZYsYgbPpw+ivnDK7YgMVEkwuGfgO4ffp2BD7HGJn7IEveu5AGz
214q8WstXFvdBBGbHqRc4Tu7171d8zvfvgvc9JNsv4g2qVa/qwpg9ATn8aXKhcVHqKD+Db2DNJPC
Ol0OrmeEnaOIGTj1WmzR26DYBR3ToAUqolI+olCMXvcWrRle17Of7bj3mp603a2s5ns8nR8nTFKx
VPOIQFu12WCZmFCSrhSjqMMrXX/iXKZK8haBC9X+NtZHOJm4MwV68msOEn1PVrGhHCFNAkdSfQ4B
Wlljv5JHIN53Xmo/lgqCwjCA3bLA3ZPHa/S0qXm3vpT5Fd/YhZwRYAp2kfvLk+cJsfS9zl2OmjUB
vl0lxDK8Tar/zD/41sd8H5mNebr6W+SQn4rdFnGVHgLksA8sqGkB+xAIgIWElnLAPdqzXMWeBp6w
sPJghlN4BXPC+anU+ZvbFjwfKhhRDTdUFI8IQ7uWjI8g2bdGwQIwf85Q+Kfg6HiwZKp8Vj/E+Max
9tLUfI6voEgatsC0t/XCVRUwDUaPmBViqU5dX7yo706TE5fNinkB4uppBKnbAboDa9EYfpXN0OTe
p6DHqI6j9KyFz2WKAsLbwOF1EuzLSDgmqiO8jKYHPBzL7wPC/JciUB3E79OZgsiJX3sIqvQ8pWYm
K33aXDgS0LQW4XQTLMTs+rCKAG3qhQgemZ+hmDXbp/E98MxE/jMBSXgaXcZ2yuSunx0gl5Icybi0
1FnsP7UIjEYsm7I7RAfcuqms/BkpoeJ9weoepXm2rt04P9oO54J8khdV+fX2XcyQUD9T5NG0pzJf
+nF23Za80nPFP08LxOFiecyTMsS2FUbcolewCspmUBb0MQvqxTyGZ2CsVvOPx7PifYoIXiMxQ2gq
dqk7DxRZXpO9jR2E32CqmYAH961w0MsRBSbuQFYD34KifAYSRbnGJ/gW7a/AAhN1K1q0a7Dwp+za
fxzeHGpF0urpN0Bjb6AvcG8pRKsA/I6fGhEC6uRg8otQlqTUv7Vqp69xO5JJEeV6w6dJ8f1p3Qb1
MsoPfaesi0uKXprbrRxQlpBBi8SmP2CEkCMnitbYmxdzTlY8H/B0zQS+UrLTQIOYDsdLS1UZWqKd
kHpItlFVipco/FVxPAAygOIt1vIe+7l0JiDGSSwTbyGXXgVcbwbI3mXyV2d58KxTWkETcYnmBHHX
FzF8BNLZLXqxkDpJFeXulEFZCQXVSQ++4d/BQIoV13CcjmkYaQVUhiSr3ev9kqavRzyE+kfPEWxJ
bLQHaaGaubmjAXbhYchCoVLsl4JzM50z9YOkOMuBOmOw/l+gMHO9KEQ5TvZpNp3nvyktXphttsaE
mA/CQawS2JNZuO9jAyS4rQxmdjbZRnwz2wU//K6ySAe/TigolHfAe3pYA8Rb9KEpARuwlh+CkK/t
1A89pVO0M/QLc3ReXTmDxSwxXSVk5zx1U4eWY+fCtWMVOt3oQic9eqYGNP++g6z0QzY+6Z9dJqQx
TRibMjsT7C2qPko+3EF0sfYMGyS/+d0jxfeYhLqNOfcD0lxvNgFJ/SDx7eq8iwDUnqxFUS97h3Ut
j29KkSBAIRjHWmYKmsldwAYXb2BQzGAewduK/QjETITmLpu4yrpGv1QT1PaNzucsSYT5vnDYs15q
L4ZiDcRP6kDu9EDyPvmf5X7Fx4KhSZubyMDwgI/txfZ4OYOxwr+a8MoWFRozbL17fYv2n8ZLu8gS
627pcWb0zL6U/oqq28k4qyj2GbUl3bZLpqpeHrWbhCJgEV31iwA6zGLu/IE03F77U5BYfYhGqhzu
RM7lFW+pxjmnZLocroNnsHKdS+9GjObF90HFoA9sPAAWZfc1HRBG9rQLO12ct4vUcM2yraG0fLiR
datXzUeCHbL3dWYCE60WAf83YfoOeCIH2cQwBul3lOM1LyiyjwKIE9K0wOMlvENfjHejNLsLg+VX
fynjPnL8TiemeCPoTT5N7+YW6IdbLvVaTGuHHnJLSPVvE+2YbIXwzTC4/fRdELe2D+s3kKiIJFc6
bpLg+picQf/inINY9+Ejb4rbAR5QJelfMHiz7RqMceLLB3KqdN9ijJ2gsaw8LZYKG8niR2Xd23kk
suc3jc7LZ/Mdr/ZUsLHzB13rU74D3jD5dp4+2QQBlNWKhXnMDWNOSj+AYcTcovoGwWK+QZi6R92R
p+VoXLJeh+f/zYL8Jx5NDLigkbQJxQ0ceMqpwQK8LTXEnMB35EtKNa8SCoCxdTYvYz1fv0U8RVAp
uZx6jvs5NsPnb41+1gCfc7K/K7qypAbvUEEe1fBhuYZGN7zOPuns62gcTZG6RL6dzJerHiG0JVlh
JqqSYPjtXbXKCiEVuRufqjRmeKMeMsNkKhkKaX9VpaNl6wnSm3TmgaCDgTtaPbQb4yUknXbDayjN
aokMykIDT+aGxk8IFLeGhE3LRdAB1rM6eeGVIUauq8Vhh/1E4uhZH1LmwaMcSuu1wf6R48njEGSM
158Fe6J/+oaYu5DAZ6cQVizIoKy8SKpY4cIZoo+X6apANOfhoXJKfxc89eYlOwkvy9rsCbrRIt0h
+YN6UVRzh9fB8zWHnNRGHJgWDYouOkDkXE67axEsH+xN8EzRJChWzryIVnDzrQTyL5Vcm/eb54We
3OrkNdM1SiUzO42ZDrnMIOE8snMSQbE1H/pSwdzEV091KmQUM00ByJ0mUA3jruxBEV3SvQLJx45T
HULXoA0lZc/eALKawA93ALfS0KrliJHDBfyRNcLPH1Fe0x0uYbKManohybpxH59GgsK1S74JQlRW
qQR86uyl4BHsNu1uoMT4UeJ2i5PEnfljzt5OYhaj4bBkd6OAygxfJi7tLM/a5HieGj7Pce+3u+fT
sWlicp6Zt3wudyx8Ur0Tz8PCGzKS9d+WXnXxKjv7AdnsNK+pnCu/cGlGlaE3ngDdKwNK4umnXDnd
/oF9D348os0QPbKQGboWy8EHBfDd8HjRJ5Pp59hHo4GnTh1vc4C2ARxj/rBv1miBJKRBJhie+8fc
D0RoXDq6OdMWD5dAZCmcUAiYXFX7kJj+YJCoQU4Yln+xf1rpCeoYG20DHmI5vlySBtQIFGyc8cm4
gu5l0d8lO+9WmA6WQRxuCeiC/TOMlHlmtfVBsCFMGddb9bHbgH2JAPeiePuhjli0SMK4QvWYeQzk
gl4RHCfj+z/UNZgNpuXmHyyX/13X1XOyTNVtitgjnyi0Cy+UYiUAlotELQ0oxKFZ71Wpn/sgNzJE
5Wwp+Md7NZdNFoMbk6TQ3jvIoGU0PWYK9yNkyVn/LAoTdsT2bpMCJIiZRBJgJVnYWaB/QvLWNGSu
7/MgrfFyTA638bqcwVN+BwtMRkJ0W3UmsuaTL5ZkHW4zEU9dqJqV6TNeP6MUWIqRT5T4WPETVvSQ
TOdfQuBQ4SVkfEf6gUffx37ZuniPtFTZhTKs6JArKsuarwR4kZ1yYpLCZKuKx6Err8I9jpxukWtu
Kv5cCEiO6kFPN6kxexzSkhbQBpp5mfIuF/7umg7vEJA+0q1bziweKB7g1QwvXDKWWd9MxE3qcigI
bE1/IQBFWpvShvE+X9AnQE4pD9cIj6vEzb6HjqebZyGd85vg+Ws/mwxT+xQzPN2uxCIm2pKinPjs
RoT+mJOEdaWLKihFMOI1I6rweESeVUjYBARbIIafaNywb0yxaGKvA2bh147NeO2bw/EKyAaPns3x
/8gnsBWXA8LrZ1ItPyaxpNBHeLVTj6VXKykzG3xE34Za4//2NsVfo+RPxUjmz15VLxG632sBJG1C
58cBlvKqDM9uNDxpGDpiQ8x7uf3/sJ3mZGuorf1ThH+bjjOcTKheMAwd3p7obQUyqvPjCH7RKVS4
31nsI204ocSNTRmPzxFvW6S1TmjUqnMW90bLmmUD8aybfJ5Q2AF6TVX872puiLX00cF3GtHIkVr+
nh6bUQIY4GBDY3wgR9posvyy/FjAlo8SLS+TLOda6YvgiGB4pJ0QZVt5PtVTh6hbfZwYGDJdTlTv
hlExu15ex4GwaVCj75+AYTrvUZ9ks0QAaIfI4bNnqT+f0ky8dYGNQgcJyXhLWyfGmpvzq1JfY5kj
DAWfmPqXpmiT94sZwX8mJT9gZPJp1Q4BKVJtRwm/kafypHHM/760owZB58fAmu4AjdklVXfROUSu
6kz2uV9K1kbHtyxEGkiIp3rAa/UyxtMIQeG+yprowwo/4Z0vwUS9RbdB1ffWeEUHxSdegjk2YZN8
bOaDu6jRFGuiQDb5hfZuuQCemOXqBAx3sV3m7clVFyQlgCYZdkrCAajammx+X4DEYnGDTfNj5Wpo
4Ns+P52+Us4vLW7NLmbeoOrc8VuR0njNOHYVxKW3HDUXhTQN3b0jX7f9Y5QSCiFzbS+MV98F4vR/
9DVA9lKSU8hmKPMGxgZ1NsG4aX9STDUqZGyeYVIJsBjpIRcXi0MLG7Y250Ep5KjNtnIqVnNr7AXI
Ta/CwLv4drUjjl1BqCk0U7fEugn2Bvz4SeYj48MgYnrMQW2uKiEy89Dtjq91GsGY0wBhuNVniSgg
4ekPWxNUxbmlrdIT5eeVcAtgeFBN+Zh8u5aFMTIIM2xWFyZMPbJxDWnil6hfyMGpcfphh0J5UwKm
rAJ6++jDCJwh2OUJDAGYXsXZ+FUp9Zbu6oV20ETFDHXo1IU1ypDWXvCyOWKAHV/Yy8JEJ5gvdy0O
HjSAAGs2boJC4Mqy2+AyM5rcc4ZjUk3gzk5dmLkX4xEKGGR+xpcUB9lkO0FDUooaE7w95vmoJ9z6
8GhPQmj1aLrJElURQFB7EGcYcWAXEDu6KvodD+RIft1SMQW3YIeamrLJsznyg7PRoFVBxe1mm3U1
ycRyl8VT1guqt9bTUKbBcQxfz3TeBbUE4FdCUbJ/QvFhDXcr2qlWYrmrh5LLQU3bCiKAv1Jpzhvo
dZTjfv6Wq9b861/FBHJF+G8l4sg7zBU0uPD/0kdz+JfwiUyeejWN6wg+OFfDn2Y++Qvw+wbdzwa+
cg75uHAx3QKhrlKDxV0aivuqN7d6KV0P0VKUInrtLOMzi+giiLPC3aQNk5FhHAHcgVOvc8j+qW06
Th+iGCgHk1ILiz5/bzoNU407eYa/yT1KnzpD2QCC0CuJGK7ZIR8JgNf+OGUEeczUyTvkpa4WgRlI
LU/xwTRkixH0IjJjUBPrigcSsTnfZHhY5RhB0036Al1ZRHXoTDSCyGLfDDcaA8Gs0/byk2mQHHoH
Yda778NbDQIrbtO3yfnL+CT67GKBUkXCcjESlowNFPUOy2mzT/HhKDozfdFcjwO6Bn2Ox+c4f6kG
y+avKNwleOMZqj4eKvjhe6Rv/0Ss9ESc2VuT7i+d088ZPcNxO9v7C+lfxyb01urJyY6MF19v1IMZ
MqyiG2dIz55HJs7nc3Qc7wn2xKN4Q+ucLxvRKzLoeKSAZOZKt5/e8wAsG+mgNih8toVMeu0IZWmR
DpI5iX+DF4oZF+qAhjT4C6lupqjra7lkjimlQUFzc9v9fZg2g5Aff9dxgapa3COwXMKzS2Ec/rl0
HS3gUNlIwBrn3YciGmQm1psZyvl06LP1DTcgA759nEkaduloc3/vtm3ofmhMK5nKYwya/Y6G3O46
FmC6lAqiBQrcbedm07ualltTlfhJHW5aZo1yzwqMJBcru0wbvN235e74O2uKruzWrCsNA7a/ivBd
pCG6WeoKsTSPmFYjV4sv5tSyGWs34LKZ0DBljJzKFiwPB7vJ/OU1CudLQsIYhWEHkqwZUJQ+EmgS
aFzfPsTCq4OC8h+sobGuskDbu+xbDKb6dXyYdJ8SDI8Q52zCB6UffZ36JtRYTJwhMgd7uvbCY1iU
udTAAHd6TZfnj0EyB20H/ZVgUyA4h9kB793R3dBreLPuF5VEvJLTUpf9zMEITNZDKdpqzJrcMXd8
Ufu8meZv223zy1WjUajYmuyOWLIR1CAl1h0bAaPEv83grjUn2ysY3I2LJtfJ8dAFHEMJGt8eH4P8
tTE3F4lhpOLgWnS2yS3csR585jO6+lC3IcUhKoYdvOj3GVt/WpFZMrQgVTCuPOiyqDXyORBFcK5Q
PBXWBTxhIe/xKtrymE1D5bkgFRL6gZ4v/6usmUXhNv8djjxDs3d6Tu36sC478LXRk7A8divlJkSV
gAN/7dvoiXidrYrzvnG1iO9dzzBPEv7DOmITKVQBKRgesYu7fYpFDltS4v0VTs2KGlY4qIJhyBnW
1i5KuwXSdZGM2+pbR5MfAZ41/v9ARx6Lv8c2zmsoWKizCKudPYRn7x/PI8fv9Z9IuOSzRzT0udy7
KRHGoEgEhyfATnKtjFhjR9cXyaJs7P+JeA89fJbrnJXGWGrcGUa8l6OozlMV1AmalzmxBPHddxs0
HolragS1ZiRf+gaIyE03uOjtER647pAGUMiZ1Q3dQ8i1c7AnZ0wQ74Rvna9ngosgIJl+BgScGhIY
T0FdojVTkDYBT0HKem0e791TTomJUZNwKb6dOsyj9st6vaadA8kFgc0XUfDU0Fy8V6WDQKDJX27R
jgo5Uiw0h3G1YISFoQKNrKrETkxWlOEOrFTSltm+/bhXH5uZUV+Xg/tL5GVCROxnV/7uoxwp85GG
8EL/5Vi3AVmJ/nTHQU4e1rJZhJkgs/T5VX1L0HvuLfovuFJhtTKFpuRiElcV0TzO9I4OLzlM7m2K
MeJKy2ErM3mewZtqRAGChAYpyL5OQZNtsaxtswJgyO0o7HJhpVcuz+7Pi/njqdA991GMA0J0ktW8
zw7Pk3+CXl82gS00GmB+GzuqkvDvSF8fme0hotyYmWtk0EgvsqPPiwRIQ58YDeIEesriC4agKQXn
N5eFNs5IPfR7R849qar0Juva8jNnNEQ3EzEephOLIZ+XvTnA+mPWuz+zy7ZCBeSqlXr8mBXQYHJy
wDEOfdUZxg+pQFXAx0k5+YH9sPX5woT0hx9czH1GEf+xUKdCYT1GklZFsa8X7ldIMKqf++dDv9vQ
acfWlYSEUe/Z2ocOQJ0q6G38EnPaku4spYZ0Sb0GT8uX1lHl1AzuPjucQ9EFWDSVanWmiwQ7VILE
/r09r18H/7KNGALoD6tJ6znrhHxZwQEjT4WYnsDyUTR+R6GR58Hgr+PUhULtIIpD0kWYqMq+MWnP
TnnnHUqIx4m0piZo1eTSvlyP+uxJR5Yq8/masgd06ZEPD9PhFYYzfD1iVUaEZWNGSSYGTNpjPmcC
WSAKabwA74tNgGlNpPxEZsHEOoHIJlwxUg6+1isWUF9ZrdAZCBPIb8PQRTxdYf/QFqOeUg/H+UfU
HsVZiykHzeg7lH6S+GgoROhnmkxvHM0VCaL1iATdAqt7r5k5jCASKFOITeal/9JQbcVSvGR1wXbk
+fDG0cF1gAq9XwN3AvwtPyPtZZixw609UXt2DFNDStKXFn/4vGR+8t94Xkezw8mH0KwSqF7IyKMJ
amM1RSxu0DQw/hsaAkiaq/oL3CmpM06PDDHkETTIkEExqYyR2buiuOz+2NKkxwhK13jTmlHIcuf5
jDJ02LW1xgD6e+jJ4Sf1P1R6uz4g+1CIUPW1vxGnrNEgXwb5+Zpmb1p4OKzsdWHZekPMqT2DjCRp
0OR6iQkzoFLz+L9UDV1RCACo/pmjtc/hQtObLcqKX41ztCfz1jCjpDVEeOPuMmyIbhsjJClTTN3V
/CZXQljg2fclfXKsMVzU0ztwguap9FG6jARKTVus4/3hxnEfXDWpK2CqdbLFL170vCa6VnnMzR3P
Kr84te7ol3oq6ZNgOWeOCvu9c9hNsDhfNkEPFNk3Vs60gmMenP+vnhLMaa+XlEH6XMda4WPFQLrm
X21pf8ubVLniJwP81txDA5LV+iqoAGlwsVY+wu6+XHRhccnU05aUVhvurHqojsaXcOXhVnXaulUF
8lMBgcRa6idtjJPjW8aJ6/cVCC1gzCYgnZjDDWNn+sfdoKQ+9oI1fIA9gT3O3JqKUaQtobkVNIvL
cCoDTwrq2XmWeh3NyWUM7fCrSXg7SaelhSiBeecLHZ3TYnBGgzw8VkQiN6wPJeFmC0pDeup+7fJt
3gHvcOHqnmYYYHi2dxCsz/sKl8kzCATVApoqYhojyyHhW+sOILX5RRb3O/wkMyOsHtWKxJuMU/1G
mIxXjtcuUPFlzp5MyHpfgLUMxJ9p6tZ77XKFpe0WJztNtZH500CoQ+tGoo3QxqN5ACEy2bL0nsX5
Nwiqzp7yg/PC/sI9kggpCqQvMsfvU2OU/nktVsUy3Igg/DjBuHbcPEXsfyCCmMAsO90WZweWwEbG
FargzeIGt4P/WcXX5KgNdUVg5vIyjTDGlvc+mmw8KReGsQbl6saUwki3TaiByHjcKYNH2P+QFjAh
y/Gc2YQxR7UwWnCD1/u8YMJ4c0EAL5X5byhK2auU4MJDAjzwcqb+nhsW6w1ojasdOZahl4er1KxC
9cGWKiEq440lkSy+/3lJ7RFfdb4ViZQIQ3NLhDah1xrYaFAkWHSHTDLdrY4G/25i/zUsSRTZ6aLn
ZcgmxRNG0iT2mXztlTBek2OwTpHNXTnjCPfPvLMO2LbSZnN5oQ0nTgryUFrpDXhkDLNzFn8Y8N+1
OFohpyBsynAK6BC5jOs3knE31n2QNLveLqB2pMPW5FcU15VHbNtszqjPMSnckBh4ACVDjJ74bxrd
at/B8ObIysZOipSBW6D4gqkJTuz0U42ECqtLGtlvQY9xQyjOhEjyPVO4vAhaec5XQc1zuMImMxPE
HyAEM7dGf4qef5TiVkI5vtdCK7Wd2jXMXg+ZcsxtV62Pfed2gvfGQEOGId45p6K/hLpeql4jSLUO
op0c3WrZZWtAHukJIQzSaDbd3Ne79+xWEmg7jmcrHi5thjkEhPqzjbDUWG7SutAXUrwN4L6AT+FP
IXl4nvplm0lJOEtGIiXeJ9SQm4j7acKGmaVP1yTvwvKJcL/MM2iNhURi4TQvm+hDXdrO1XfohKin
L+XPeW8CIzLxH5tbj+aRmdYSytu5DKQ0dT33wWVDTKYoSDT2rV/dosAkKIryREZgZT3CZ0xHrNVE
z8dNNhmJiEjOiSp0cgu7HuOKrQ5gk80mL21KjgnzY0WgfvpYp3IaVzcc4SZ3dLAwZhecFIVoIHEX
NbEE+yZ6h3VYOfKx0AUh0HPqOiwj3eYj3ddGvp706BylrTJeg+i+vEl5dTwdePAvGbzyCGJcciF2
3PQUVRoDB2P/x0XzpQftOQqXflPEGd789sxNnsMoJ6KAsUlNJTbJpTRi6qMBq5yi+Na1yHxzwt2H
MiNtMXMFEPFrTRLGQBXG/t2ltmXywFD3oDVZAl6kcF+qsYu+xbgsTHtEK3PfFeZaqhoXEqqD5Rev
zuEGqcQbgtlM4wZLHF91otEEzLm7QVxsFtjiC0DjKDyMyjLUJ9BZndnRfs6udWSwycWfL0B0ggjY
d8XCdmnE97xnRO+TCfxsXn1l0ofxspFQAzGCzsl+EWNQ8rvKT7tjo3vTlewi0ZBQFmi1JTc8zxQO
RXKnKWxG9wfl4d65OuWK7dwtx55eWilqtJNhL3SsBqiK6H3yz26dYXKFDrgc2ZiVZxWCxxXCQ2Zn
Poy4YrqQMjJgeVAsVbAaW1zc/ig2y2ov7Ra9srbmz/KrO1cDtdj8qQZufy0oWboufSR23QbkAXp1
+A1EqVpLmr26WpUa3aVxRICrjVNM5Zv62X5+XJ8qISRiJi4xLmfM0F5Jp/Zo8j7NvbxBP08Fqg4W
/dntU43ulayPFRdvVbxYzENI3Q5Z0RpA+M9d//Ihtga3b8X/HYrXKI/2cVBxwxusMlUvBA+sEq9m
RiQojoZ+C7XKbZXXZ/JTt+ElTYExSxTAD3jh1jhA9dqpWIA1ypx+Y5SBgM3RYsaLL0KxSvr6d9N4
BB9zXUBoFlCZULRPtMhggMkDO4m3R5V4GuU1g18P2ozm+1v0XI65koKohBAlAzYpxURgzxE3oxZk
so1xLkYv2HzsY0JheOCbprONIWcx+bd7V7gpdFMFUtTmgjfTt92bgYkglWXh/oCnlgFAi1xlBrNM
Jtc9JZWy/ExRfzewbBbAtB6uQUMgQhOPkYyuU25FmaS1uqi8kgK6ZYdwlNK4DJn+hlOMW7toD7VR
2SpRPkakvHVuK7OAJoKIBGWhx4/AW+0kg4CzwibFcpI9tTseB+8TeRA26/fFP+84cS1MqQzyvH9g
TPjoZdsEtXj0zwonNzuTksZfU5PXV/bfCKLhEw83m8VdZgTL/NKgtXgWMkQxVoDb3EY7CF9HgS6y
iftuU8Rk9HYwPeX3qbc689CpqMP0f6/qgJnY7u1L4NfrcpTF8IGcB7SREfC4EAmJtKbScRheYOyp
0/CezCGPNlNrhfum6GxlK5jeZfO/gkUyGn7a1vRgvZk+jkDFMqVQSCcItlSmZpeYOyX8VhbtYc0A
/VXGM2mqCCyPF1KhfNcZKJlMFq4BeZxk+icblMbqbj2jDPHs77gaVBAQqyIsYvhmcsXardcRD6u8
JP8ANG95oJtxDLLoDK1nj7SSftNfMSbxacmkeX5etBsVks28X2PRDM2QuKOflxWsUWBZn1xT5NVu
j+PwmSc/RZsAQQSRhC7Em1m2qALapi9pG0QcC4jE1RxXxACul0JvCrP3ZM59H2HUNeu3F9NiPsc6
FiGKqc561ffl9eVW1znvZRS4IajwLL3231Qs47lowUup7b7QttY413QfnBNNxOv69Up7ePRMm0/L
yV0j8ILBodevOHHPC38hH/bVNx9sowrhDEy6Z089yaxz4+aWcuTYRzBXlgNhwYBkYlpofaZS6U94
nsUlVn6bZ73XXSKQwrLEkhbxMB2KvHuDKTiQfZ//5RP+Y9v9hJPNFXpFa+048PS2FOiIxO3xMaws
/w/x7uWNEuNH+VOVx6f5FZk30IaMQ65b1ODa6+J+4df7fQbX89NimVuGk/sZHVzqhlMhle3zw5zI
lq3dcCZ6iurnmFV8oJuH1K6TANrnqpmJPyAKsDlY5Y8IbbW5iyo6C2MnKSsy5rjCa/E6RM9gaHDM
jJTrojTZNUQJFV9KfA0Zln5TkCsbzvTnnGvaLeqpyDGZ6eIxxvPyArh7J36ak2YlVxIhN0d/QfUP
/FITW9fHqtNUAFiVoSrFM/fEDdMqGivj2fHdX28WkroNJ3Denj/g0H1YuO1Q2f68MjLSVVBiH+gA
tLVhsh9ZZxKYvgb2LAWqXkhCfhI1/Q//UaWd0HQDbFFCznG8ad7aqQLrPhcBv2KinkpM1QpF1quB
c5ugsIfGgp71kINKsFcErstvHjtQOX3KPd06GNmnmLjaQavYtOeFMP31Bz4VG29E2XJlEIvvyxeG
1RD2euJnF0D03aTb8rD7f6m5qCo16wkFpCaDVQE7eB8aVpZk/RDFxyJoGe74kM8LTG0TIgzl+fUJ
m95nSMAG4N0/uIfRjOkyKkDe3gYcpc7kUjmeKlzt1T5XHeLXZRc8jfFquLvRkVIWh/RBKegLRKod
JYQlSlfGwunVhUM/C9wHDDspGVYLjDr2mWdsQ/KKrPuxvxmp9PV3bL0PNbDvVGF64pOYv9gKgOFr
czcz/90GIdriqo3fySCNEF7FpWSTf+YucmIddb/L5nQD88ymuSceZSAe4USK/gnahj9dZUG8/BEF
qnX1/bshdpalRNCsUDRVcd/+ePi0TKqrJxU0Lq1I5vv7d04EdARn41w1pAD44dvmHGC8NmgoPzaW
nVLLXJiSVn6FeO/k7O8okKxCiDc8nvUabYCNbdmUXDBXDOaBX4RZ1i/RIvzVuqCdRjnThViwpWDW
mlJqU65H/O97N813z2bpxBWsoLWwqD4FUwZqh4BsIb7rAHNBJk2eFjcRtJUx/qMpv1ywiCt2lAX+
V+oVA9TWMoMGfjAYb3FHpQycNMbbUYm9ni62Syxbph+98TV1bE4ZumQ7TLy+MVIZ9xLsJBIzRn9g
cfVxY482w8jTeH87ZsiZ9a96kv6N7jMiC3Ydzf9qzR06N2gu1PL9OuKCQAr/RSYzMFgYgWqrIyW3
mzqpv1vAmezeWZbpne7z4RjXwm2Nxd7/SdkScY9n6pv1yAB/ejEuFzN9Jowk8NxPLBmyASolhvD7
IurOrc0p3ICfaXPgWaGcjkfiL/QFBFnp5rTJB475gVTLsrE1g/tZ3vu9Lnra41bTI9wrrlqO+zRw
ywba25M+NUoisl7v8ccx6qjI79k+lzhx6Q9d16R0ei2nMKOU7axUkh6dTSLZFwK9Od5noqG1AJbo
5RWBozCP3m1Mcz+pJ8eo+3LvOWY2BMm0SKfenNb5CkuvTXUqWfH89Jv3pzIISYw978RW5XhsgmhQ
MMQ9y1qrmffjksJYxwlvA6g86o6cKIe4VD+EOXYYZ2Cu2XHRWOYe1ZqYM19vH0hS7KOd1SnN25qX
ITwMqamv9oSC7fOMh+y5BvqYGV5h+m0DTO0eZopUSux4h/0ZW2iSePCebFTDPRAF8GnehzbMlNH/
9BtKhuRG5RYusXjkfq2Ge4OzVdnQgbUmvPvgQOUZmWeBnpce+Q3yGQQcI+Cx8tcE6E6uxuyCIz1U
G9wa68xjjolbYqgjfsb2orm+P0MUrHncU78r7f5RbDYMHL8TxY1Azh74mCRFigxUZl6JEJ/Jqglv
UksL+HulpE7W/QV2VyDD3k8qREUOjD2rS5Ka5TM5+t/0aLWMfU8NtUaQh+HND17aN8q5Rkg+II8f
GHuQINCvOSbdSiq9B1uMrlzTjyCcJVflI6Xa+qm/YANLiU8OHEwbe8efl3kxztDJp4CFLKryoFDb
24r0E+WMDgzdZbE/K37uZMDupOUFl3ghM7L8SjJuaGQ4ZRWahRs6F8upPnEYdK8LlyhlQecq0m4t
tCCZ6u2puZ7ICVu+LOFnagsUs6mFHgCAskIu7KEZSKdzxUnU6/mqvGgo6q8LcanLz77eV90+kyc+
6kl9yI/zstbhS6HlXoR2pJVegMpZadIZx5rX6HvS+/nShLT2Wc0AGtG1NPsqqXQHCT60NPu6kKDY
4HNOeIGijwmEsnlg7PJBqxvn4aWk2WaoRXSSYFtCX7E4QtVQbj3MuCHg9daxWhPDcq4jQ+srWVo2
QOiTStD1H1EjV5BlnVeGUiCASoAY1wVttFGPKMWzEVdcMxMBWKYQX7qlXx8ONtjFRAOXMuk7y1ZD
gLvKDh1eki7U41KcWicvtGFE2cOv7PeNk7A60ha8xEPAH9Zq9dDlMSBLZlKVi16ho1odKxPXx/Z8
66i1ND7/bUWpsWQW2p1EgoGwjt77eGgE+J35lt6OyG5uoEoOqggPue2aqY1xXk1198yXfk6DgvKf
ki55lRXL8AEvL00l1np1sEcW94It18TyMVSM/u2XQY/qDvk1/GVrXjQeZUycua9pda3FtkokRG2i
NxygV638s1dt87dkALacDMGUmu870xBW1tnCZjbqI2+iYFvlRsJAkRnbglzBFCxfz0R6SYemOClS
2wmxfzx/x9FrjCgoL4DbJhi9KlwB0zgfSfeseeUbWu6s2+T45Yx2L1sTillVGAqZL5pGGgdh6rb7
+i1hX7wc2myAwkfWL9DlYfvxe4i9taGjUthVLtkE4kIhspLzlrjroMdkpXjV9MANxu3/pMB9mEEV
czrQvZhezvQdimixGXzJ0wLaHOFZC/loxDVnEaxxFJd/XlruG+MgK38YiiD3TPdFNIyuA+bs38b/
mgmVqXH6ZYJuP378yazCd8tClcTVOC1YFW+opTpaMXar+++6uUCINaUdffLHCVH3N1XQJD6bbTwO
UiQlDyWKd9x06WsCRQz+s75kGxkHiYP/adadnZVJd+6UgmJ491yCUWzVuLpV4JZmiY85rE1mUxTJ
jDk0drYNH4CmWhJz+4tKpVzpYfRrlKTTH+PlVZ3zEvxfyGBtMW9kC4Hgv4RMUZoWdePYeIw2oOta
9TE4veZ4qxfJzEBG7JU7UY+TJbb8Jub1Wx4kKXbZKbSlWYDaMSMSgg1Od4TZiwSkFTIQqLDUB6x/
TMyPOBkoUkp2u7+1r3DQBeRuF4EFbJOk//8mQOQXcCq+pHU8q93h95Crgd0csO8RIRs3FDuToSxf
ahahUS01BMcHzBSMJrV8+zTQwjZn8Z8Lgo/F92Z5G8lEiJm4OypCrNXcC+q2HQKvoAYmvbEqZbxE
Tzm8wLUZHemCPZ3To+03oNAHB6rvHoMhDlVpJMNbgD6s/39k6/yM2xRD1EY+x9XGqNgYvcwcfHUj
DF93SGAf6rg7Ftg1OrdhyW69XWstIXJ5bSzdI0GbYhASvlfl6mi0CeaUQI+zvSQnFLrck4yIXlQk
chLR2zf8l4DOodit+AeBl93dKzXSvXGDGBlyL7r73+hggYFmSqRpa6o+/OjvJjZl6qoKxQbaQNPY
Drq4En6ZsHB9XS4z+nT8/N+dd0XS8M5LDlMQ4pd1LLBbWu3LRQFedom41SRQZsfa2grt76JjLUf4
tLjO1egPc7vzfs247IOOvRondP89InnsdNfQb46/IUn4nCjllltWuQ4vmBr9ijrIlQjfK5tJvNmb
fBRN4TORlzAkKPBJP1NPgIkbgEYp2PNdU9kalJZ61xv6LIWUMxMnpIXL+JiuAK0bPVJvEM+HgCEw
ke8i9nD8oKYfuj9/Iu9jaBbZERQpPDPZvFndmKgCLU3sOzxpq3Q8G2XGYHPLJUmLdQMTWf8Lw2vD
UFswXbnEYONDHnGiFpoFfwMAu8rtk23dooiEn+eRzKM1i9dG6ibAlngMMAuJXR+bj7oRDYlhsgUJ
ny/UXPwmYQAIsbESPwCjl+5q2yEE8BAsf3Ha1qEP7s1VhEdwQtKFrsa6L/6hTe+jX79cg50Z4z5r
9a2ZwW0fOL9qbIJW4NTTXr9efyWV2Lw6bNUWq9YTiwRqj1IGFHEdHlDokN9kTb6mHNShT5oqFRu2
vMACpEOYiIZ8ZMpT2CbO6BSuR1/D0t9VXTEbIGX7N61/QsgmBK7OW2oQFNc06LKAYpy8/p6Jtgl4
RhxJ25rV9El7S8DI7xPfhPgG8g+wByccVH6qqcbgr2Je0eJCkmj6/7ELjHZrPwQMAYfEx82Epf/0
znBayEkhJG4lprvt8C8arLrjRb0gptn6l2eax/8cScySc1hjkRUeCEtC0uVAsqCpusPSb6x5DND2
hcGdyaPFAL/kJgcCdsaVZAQDWA9bC6OZPYhQMxcw1aHlpjBUNdKu7OLpGSHxCQz2IhzjgusK2ZmG
tfVcxUqQhesAHA406MoP5C6SlGpnNQ3gwBVGTnEivTVnkCe1WT3EKcOSLVZUzlH1AfUR026yG1mg
upbgoPa11eCx80P0gg3ix82VPbXdeM7dtYavjqsTAIuUksdtNBDzDYdVZDnyZE1znNbccF5vwsHD
YBaQkqT/z5yYBGXAEnESrHMp0mGlyYpOQqvQWg4XDeqUHlm/bhOk/cnkJ8wMV5pw+V7v9QT/Ztcu
Em1dzYzxbdz6f7aGOyKKvncQky80MfM5GLuS3ONS1dwmH54C66YqzfJEVtfx+sg6rhktOX0dXdNw
8eCaVxZH48G+xeCjTPDs5BWOO2lraLALYofNNS0VOCM9z8Zdk0m/phLluax4m95Cuj/4Qa8rm2J9
Gh71OyWlDb/bWz7lI8CI6jvpJBwt2+YCNkVFwwsMDsXul5qiAAd1jmCY3eMiV4QpuMkb/dVKJkzw
eaSk9/GZlsMLUGGLdc+XiZllmIPRwvrw9koufI0Q/xc17SaBc9F0g0tV8P9vhaUJGylIHhnAWdS8
f8HTO9fh1g+ihsKpotYBuJtYLmpgs8RWho5Uw3Orriu9RI3vbEc1hnlKr2hPhz07NVcY5RGSunUN
KcAsp+NQHV38jPTcngLdAYpWX5MWacwKVvJ+JxJHHgtqbtaFssxegtMW5wxkftp9uVXSqAAfirLV
lFzgGKkKjr9TMNpjB6DZMDIK+60AE77c1hRX3o6feOYITflogkr8bMNK7s2NDElYk7AnDja5A9W8
+v8EwWbSb1VOJ5/wHB2lNbN/uchrOVdMK2Y5JPsifumEw0Jn5dNqACarUZoiEQQtVABmXvJCm2ri
sz8uG2RNrfKxlaTvmbNKVMHLt9IwE+ukAlMUrPggpDuVWaNG+4i5lPsInNap/mM+EPY6P++bf1GC
dhwb3Boru/2UygHx+Ke/5qI9j3oMlAINgpssUa+7XcLUAm0rkWtF6ldF3f7fccFyeDyU5YFD+uvj
DQ5d3B0czRzA51Yc/JbsGzILkg0n7fKylid+7xj5ba00hPmBF7Grqd54/Y59eTN6uYfyl7CRNeDo
dQGCbhCVt2eWjqINmGfZf6p6EJqjAGQIOdIninb9zaznzP1eRpZIeqSGTikfmNqI2nWYKBQFbxUu
e0ex5PGBSdfujXFG/7WVVDUPzUwTzwEziaU9DJIvUENvYqKxChO7CpwtV5VoQ0dTreV3CdTM5L2D
t+pKsuw/IOg7qDDNIpcR+MekLnMH1r54i4MC7EK0PUbzg7bhmTclRiyT9Ds3v8aNsTQz07wALseR
eAOdnGesIBGxujPVACZMHRkFxmzALIETLV1HOML0SKRhPNnQeRGTdU0b4rVQ/CfTQG+LohGl9ifT
6eSi5oujBnMEQ35xr21HmglWyPwd+XOVvAs1W0/G8Rv4z4rFROa3F4hMCNNFotfLcU63rO8TY+Xn
FE+8P0dvi8nn7ysyZUL4UZUpcUHQLX4CM6SKctuZJe+Md0ZN3RDCfjb+mrB6T28tjb3TXUpKzSK9
nIEA2gUSC1kos5C34iDVCZjzmJ/XMSblOLXDgrUO9SNaV1VFl9l1ckAkyfHE5z0FZ4kAG9bLNE2E
MqJHwSn+U5R0jqhHLmcCnrB3HPbD6aIecjhTM73AcsjruAKUwyrzpPjbckDsVZL8E/zNjqC/aRRZ
hLKoQACHpLRlaNX1ZZjzMB9+zr7D0FRsH9vAvsE5on1WVUw3eyzQ1vWZCKrBwnQMa75HnU2B/u+T
rsOsoaR5M9Oxvcp4vgdJjy11CWNAp7yX7K24hR//q+7omcRFolAPWOMzfSXBTtBbTNbUVPe9A9QK
6bIaRHqJLXRpkgBmNrfJBlvj+T8JHUeI9pFUS/V6vluKRi79Glhh1Qe1UE00JfcRr+Zf5Pp3WeCd
GEp7LyzWWGaXd26UysV4401AaOdHQj/pq2OOcyIpGixE2rSNtOKma7eO17CdeAefcI5IAVgHn917
fRKUkbHwvC1LniAl0QwO+/bS5vy3GxAS45ICnCINFSiJ5YDMpYniAI0n6uknS70Chf9we26JFLew
8y/mEUXZ3Od0VDHYfNwS+ENp3qkwDF9BTmeOvvgOHtltHPhtvicM+rgkCwA/1BFXn1PbJ0/Vqrmx
x7LNY8M19utO0ADbY4Cw2Kzx1QQDI2USNm46NxVShXVtbKi3XGRCYcuxLm1TzFn9ed3K09QOZMsD
evdVuSHrwDpqmYmtBD/NLrkHiWeJf6ZnPrt3abK0hgXgYu7y/dHIaw96AdwejC809fGQEv9s9I7+
VshTIQK9REkQThJwuSBDSw0E4AlKz4+6++RGN5wOZzAJrK4xFoux3WfbzKwUJ2YjkuFKviLmhxy3
HZlt4TsW3sL3047FaQJB1OIXNOL13plT1Itxz5y3jXBacmo8OfFE/f2RwWXS2AUvioApvd6S2Sfw
QqlrPxtdr5ui7R6VMeTqcCi7/CKUCOtIjFKMV/yaEKOeBPPzSPgRSzsZk+pZ7sv7KaE8rAGROgnf
vDNntZt+z8kdzZCHxINNlIYJcYKvDul4jAwFG8RqqqSHGlqGJvVcoem6nO1ecA+rnE6/MG2oxhzB
POTxnM3t2bm39oz9T/Q3YOMOUKzv8pJl4frx49YEkZKTsQV971UFxIYKVcqyfa7ZvAyCkgB9olyH
SSruOVq1wIljMpyL8M4KDZ/riKtoiLDQoBZOqPaGuiDrndTIwPF/7f7mlhgASpBcUxq6kO98wNqa
E5GPcZLUZU+o6iZtd98p1Zg3OvdKDMvlDEvywhxqaa3I/w2JKz+cPvDQ5nODsUJPIs65SLlqZ52W
dk9tY1jKM4/g51IZ9YDF0ZMUIw+NcDn1Ubif2WF9U4REu2egLxXkojsZ9dFHABvRGpUnBHB3+kHg
MuwlKdG4toKpApwzzyWWWbN4DcDJL1/XArI1c78oXUpffXh9+Eg6b7CNQ/PsBYQCyHjkXnwh242x
it6McvNXd/v/iHJMg6JVVuocWm3nI9nJcVsWhDvOjRjxx6g+etceqbEnF/ujKsO6NvoSeJNXPWSz
ow2VSmzap79nxo3QmgU1Skcn3BmFTPAeESWx3J/pW4073bNvyqcNbbyNtEjx/vku4A+LMLDWFTun
k4CGclA0/4ZN8sj1658htiB/qyXwKhQDiIXS7I/SH/eEbOFdo2/1f6f9C0KEJ9+EccDnDv0XUdR6
UMhDMxH7w3A1J0Ra9wADC/JuDc3gSBuOkXFV3vJacIU27qRojE74/ksugDTmegt+tE2/bAvIhMO6
/MmHX1urmA5pi3CqwqhlCGTuVS5BX8E33a4FcQg5SnwTIRq09KDRtW5Xip0tyLOs/9N3+lBLiU65
sCgVSZtWc0gaWG6deSY6tPgglPrvcw5QdIMc2pfzg1BcwwliJseHbsyk8tjEWjQsqqUViyxomZiS
uxGBTPL+wdfasTf3YgaA+1/nWKwbKz3+J4L7nTIcA039clp6XRiz5JxyVaKUaPdwuuokcJ9cxeS+
1LWKipU8K17b1O9s5WgMIzu5/VmDz+4mWYql/uF4YFueqVH89NcaKen+ZF9DNce8BWXf8HU22hGF
dIbSBhtuVQPd77UZMFBltU/PdkKZ6yLJFEZSiXJGWTfkOKROraBoNxNYc0vbyQHNgtdX3BDYba6t
iN4lgqe3HfoRlC0MRpj5q2DHQZKdISgjpMCsrz3h1yeU/CbMUiQq/SZJif+SmHSLdl2Nwp8geNbA
+mnzKxQlVA76lJXU/L7mXkMpuLxRCFOqUGhiAXOR8QlQ79Sdmal+5UPyi/0ZPd9sBHOY8E6tAiEY
x4CRBc45rRoQ5oMbXfjeXP2UEMAYqDacjvIWPJuOyGVAF9Hq2Uo3RQLHj0myeerwuwNIIpdnqN2X
4fGMcAqtVVHBXQ0Jjb2LbIPghaY5WGD2eh3S+i6pVbU4hJuA+NKS6KEwu6VyfDPqLcUfhqvjtqOU
jKrlAH0omMcmhRDnrzu1u6VjBZxz5zm5wvkwHgfQnFTGaMbPCRFFOODcLXuajgOiPPK9eR+7GKA7
M7JyQJ6FU8ujYHFXkYRZV45B7NI1wUYuiivR920W6HKPIlPnZg8AaOqJZxwqte3uLkFYX1dbPiWn
qH1p5ZJbynwrq6iNf4hs8NEB8jXNmvCvmtoyk74uMymK4KEQWF4zCxzHsZWFATpHRI/Jtr/+kBtm
pYkyzmdLmpG/cn68EWmOxSQClSoJZnDy/hWFWI+4mHNQdHGfA2TYC/QpjhmQgqzQJLAxV7HIMu3z
+UTKzf0oCrB3+zkNHXe7rwOPTWuo4IqaqpA2QZp2YWpZoZ2RpYpESjKyxQeMG4wtV9kjfQO1o8al
VvsQ+Ec+WUxwnutIT3Y9rmMLeADHe5QNX1Zrfuh+Us+sSOJBLXSTd8phd9KDFiN/STrOdx23Gllg
RvcV6QAcG6f5nOGkU9cETf45KAxD/paLcb2h38mx6qBLmjc+6IskW4BGw4f84XrEcz5w/xvdYDpv
k4d3fLi3Gny4qjar52Tqc1MEWRRA+y864DNKK6HVxVs0vqSLgZ74ic8UTdxCrIAepjRvRiLTKXps
FMyEjkurFNZFzhAdJdm2czWfES+0pPbLHpkJ+TC05bemct6mhXWR3jt4OXLEyGP9E7wwQTxrrbiQ
hPn6Y24i9c54cnXdnx9pdGN3m9AOT7t6W/09Al/mtZfOtwcM6CqSAbSFnQO1ZWodd5nXlJ9hneLH
aP4Btw5Q929DFquJzSO2WlMnj9QVNXZzMCuWGQaOr4QqvcXJtWVNvREnQs+TdgRZa3zmdei0CqOb
QM3bYZ+a+x5sAVt8iQcCGqjSOcwwJRUjJBMDXWhCYOXIFVRltzr1bYLrG8U1WTV6sXD2Mz6JXsnE
aIwZpuVDR3LDirEaPsodXhLXZkBuyAggVq3y0eDxZ6l20GgXrHg08x6diPDqcqK7n6GfQtu9u2qj
1UunzvznvuAzedHz6PS5r8JDwz+eB23J7f5yXUQDy2jcUrs19GjnSrffwJxJL9NAdvCIZvrMj8RW
1xaNrAy+0a/i/OYxwYWdX9FC6wTXaKsO8lJ+yECDU2Kof8pVDVZmxB2colcHOYCrzVUi7cOlN2UD
Q2VdcuVe/YBXPtI+DMTBWUTo6yAWVXZPBJc1XTvfcD64bnhpWY3xZTz0a0yRev+MwhcBBNjhu50j
Iya0zSzlHZjh1xk47DluIAxxU9V/IhwXyM0EbP4qM8JrdHZb74mqYgn90VDVO2gPRiWgvvg83nt/
gZB1McKwdo+Vzv88ovOyHmhB0RI4sphxKPo72qOGyLLWD7GepVeobC27w1zklNZsQA7R+Ex1Enzs
eqs+JiQ8hcVUtvaRSwsPBd00wvYyPwKsv33aYl/1g4TFQloxhJMg8Ceq8ini9yELxl8WYQqz3/E2
LvArZjpHR1XKKAeXMbLhoPTbkJcvHYZOLsCUuvJche+dRL1oolSagLl2VozTZrOkq1UifOO35XJu
b/xZOJv47X7eyFSi2Ggc4ASHVau+P7cONcYEKOU8EXbL8YXIE+imvyl/bgRnIZ++8YDxDZD52Eke
9ZyHpRBrmoiw+Smx5wOg/sHUERATu9yXLg0xm10UKBocY+wcwk/OrYFr4fnYxs3oOn3g3XHYvwgm
exVqrXn+kC3qN5BKJHPwmi+3E0hCsCm/TxiwgWo2az0qxqSD42ADRfdRLNqMaI49Lu5i03M7exdZ
WegDkKSHGjVFxE09nCarhI/T2VxlKUquuY3RBHbLhrYMKWYPUdx1IUtNRK9Knn1OJOgDmIjciHaP
6Nhzdw9oJMUcTGMI1lfYmy/psIHxJ3zTkJStfkx3o4+SgjpurCwqACu7aaouRBsrHVehxW6IYBpp
ypZEvn/tqjGL8plJoFQYNu1wAxzN9+DylZooXqQkSTbEezrRymYWTC0+eIzgEjkPtSOtD/Z+q0ZD
d/+UodQIdTaHRQfq+YNMJ5nn8fGAGmnimCcvUNaaTt+6VwO7smvRVE224Eke5wKE/Oshg8X+zQ7M
RKpWNXY/78NNZa8dvSVzgEZLRURx0Cdtw0RFIUS1n0h9nq0q6Mnc4mmVzVxphm1oAklPJM7ShGCp
5iVrV7bQ1BwzHsVBoXLUiVeiGFF+4mMjDF0IWmEsICjcYKAEFtwb5RSopnazpiX4Nl0k/1MQe1kV
LQzYROx6qcfDIxewNUuhh1e4M4hwyl5sfVMB8wHTO2n2nWg5GwOJty+mFP35ratmEqDsvZAore2I
xjHI0dRoKiMGP275s+LnqXea748QJGL6bE5FusfyYd67wFX+xjhR2ocQwo26e5x+qbtkj/OUSK1q
gwR06h+b9qJmVK3hkJPpEQvMH3FbWUj2aK3SRhPrS1QzXeYaD5oEzqhMe5YUZHRAlDQIAKAYulzQ
yZagWd0X3xy9D9uWCNs1RH+xrVy+XZtKypibS1E+UU8Lttuiqdj2TtgK8oVH7P/fi98V/Ec5c/ok
9xmlI7mD5OCjhMbZiAtIfVPgBraThjpg3n9RIR0WAeRSnOeKFBB09yyAPeXSOELF/5SBEsgJBz0E
JqiUtPpQAPHAZu1nZTGqE0UCeTWmG80rQ60aou/CpNRIFLEd946PTwTaqTcrQcfvw5PDOnc9t0G4
qx7Ggar1TLSZlfg814+5FmRI2ISt+2k+2cwCYOjjahut1x31BDyT3KmEGDCh22o4E0ykhsAf3tGX
T7dXkc7RMpuHZ11AOK9uPxgEYZ3LSIgzKHvw3Tsla86Hemb5W8jeFA35JkjjDXKb8i0PkDpT5iry
Ls2VZ12bzXqKEwkumtE/9boy3+subsYSRZIRQ+Bux66MFl4WbXDXl/yiFUAdsNBbgOfAgBAtulLL
U060zowU6cs7nj+8ZHdyn6QR0uYPVW6IdR5Nca6faFI5GalBERHCM6me7aQxBFrv5o8Rk4dpVhWa
GhZrivJivrzNy/ozXbQKjhcnRO4P5HNGT5C8iyq/umKELbMoKkr8S7tq8U77nbyYuQgSKAr79cCR
ogAdJ3TCW7W4dQeE72havDlJwK/9TYoi3ftZloHSWUaXuYHiPCn/dgzT+v+mQXMjpBUo8N8FRjl0
KE0Gm351ewI3V1m3SIrCzjOwcz/A0+Iu1PA7kvHFmAzo1Xh2DGYcF9LkSG6rOo8cRh7rgAzGL0s3
VarNv+nhUFnfw/COwT5jC6t+AwqKA9d4JK078BmAoV0qQXUeiZrNTOYtrTZfKwnxZUAB8cjkjAbX
+uwWZUWB2McUvI/qJrtFfHcK55IALoUeNKB3Bl/PQJThvYOpzD2c6hStZNe4wMpQU5eaNl9+yEpB
BCICoeJwFHEr5HiXiTKS0AhdEisauDiFqR4UIlhGNxXOgLL6QzKVAJNeEX47rGwopyl15Hrga9pE
aAC2TbaT9JO4rv0NmLUTOpzODPPF+Psac6V1/3ORwpUSob89IvcpDOm/eWXLotUs6L8CU+xCMVUL
XrQD1bDnxRVgi9+zs7ZMFC48WibxO10vAOfAjzANGmdhS7Tdxg17FpF3n8ZNkPfPiaDFOhsYqtJS
N9VC/e7dXVHXiKZEHCTPOwC2FnK2KT8iiyqgNrDDFnIvIVPKsmEaEMIaja3lA4nJYKbB2B4Kjr4K
qw3S6h5YuZmqUdehuOdTVethj4ug3O2IOgnnIbhmAueKeSQSFP9mgI7QqMy3WifqCke4NoNvoWnE
sPjjAXdFMjKmeLMOoQi/RcZfp67tOv8PIq0ZxQ1CB4ktml0qIfd9QVoZNbZjFN+903J0EReP1UUa
frnwJ+XkmHk4kgVAGeIwMCVRFFgFynCciI/lg07K1aqgHIZncrNktjnSRzSYjInAhHOTyyTKZ+wI
EusooMQ9rCE8a50KPg7/Tk7YqjIwDgp8+0sDalQvmISLq7zyiKQy4hasv1p/zX//iYNyjChnFJpk
eGzXFLpT2ZiHLEMapVZT9uW+AjAPWjZFeQduywqQM9QLgkasy0d0jGmr+NDjjyAK0u5QXkNyHtMq
KDJta+zuuUHHuAa8WtTu81R5emoT91ku7lZ8QcSsM617pUe7e8gDgu/sPxJVHsRe1cdTHGvTT0x/
ADySLYFwUfYWTOC7CTD/K/T4h5GEwcyv1Z9CIByBGR3Epll84cyGothZRLjPvCKbb6CHScE+mI16
O+XcVkPJtv/HKNF4EmbeZonQerHS1RxiZzEDNOdOFjZFnctIiIFv5/VA0NP5C2SXxc+gfSa5K9ue
U7WN+xo4sWQvrNWDo5qTltTR55tFqPaiAZ9Wr0uf8Qouf2DRyb131nwth2TlADwtajRmhP7GJ8v1
keAD2z/kanASRwiJAAkua+KvjkeLaEUcoOaj7jz1UzQj/2V4f26BebWkiyTuiWgEby0LG+CKBfSN
mRTSh9czkz8cagwXqKtMp5dwc8tc5C5gGNv07WLrA6PkPdjGmF8ymlZ7c/czXakmxmNkH+LLgOxi
Xj0R9N+9+NcLNZyq0m0d9MBeb98JDosDN+yKufIrlfiqG5YDnB3tjhrZvxAmva+H4xLRCBWpgY5I
VZXzgd50AfDLobZtXQtFbVu/9DHV/ZUZM6PZmyIjdUcmsvw9BgYPk8GVLmaP9wRS3pj5LTOvylYz
rPt55eVkA5ecXdhsqMm6oik12UdbKRfoWAQY8+uDzSei1QrtcAt654oZyWmG0cuV+JPDJj+QaTXx
BbKyaef7s90fouyONzvEF1yn8lkwd+Ob8MLrBK3YTncxU+lcIY1BMUF8rxzHpD+1HeVp53hvlnlh
a99luY2LTxOwrX02lbEzM8k3ucpoz03KITdLHGIYqDL5H7ZP4BU2EANcGK77/tmOFGrbBNjZ0zi/
qFsoWO0R+ihpAkVnHt4yvCViS/NnkCo5qY9UoJ0A09yot9IVJZlXs7BtI+oXuALC0Z9Bo7sTh3YR
KK5GZp5aHyd6k/2SXT+/po4PCwlPQNW6XZ/gDXnwG3sSMKXU4l3RSzasdlluM3pEfisTsPMi/2N3
VAHDztc7X54d+fXuJUz/NAn0GbNYV1tUVhyxrg/8zzkmWJqYWGM2witk7NKi196VrO/bLy79fq1I
qnANg90R845iR2BnTNTuCRPeUzGDrtyUtHwKCgQY2rqaVjrfGSmt3ptwvdYBZ/dUdXyTN/E2rOqR
AMdP57Wu+4nPZkhunoO2MhqyNpCoeBokkN5NrZI37RSvpqsWL5pK0zckTIbWM0ejvcvihZeiNGJ5
p1ApaS9+Jloah4hY+u4JUf6jyzo5JUyBOZJ85NP1E0UaxEtSLlioe4BV5MN17arGc6GuUU4KsSG9
KMM4n+IStOOmFhLzTlReqPhuM+eUmO9Kak4nTSzw+lVCqaPTIP0JRkt2mOWOd0+ldGGNk7a2Y6b7
lgtNYvu1rISIFU6dgaApJZ6bncqAMwY3Xdmq7yGCRBsrd6v6JblHWMaJOJugV/8niIefaQKESwRl
NTng+s67b3C6Wb/YpQf1pJwUUiNtHf6uK9HKQhtQv3ele61DPOF1CEcCzZOphr0hYtK6JBPyEHKK
xUfh0Pu28yBF40vWXQMRcBA0X4P84YJpWsLfb6zx/D2RfAmHF8QCVJOksnrzyf/oC1SfrCQikpW4
k69C/gzEkFTLq6aXA9pmxYds7wX8eiOdrTp/kieLZeEyog1tzTOdMPTuSzGyAvvvAo5t1pW5sfS2
P1MB9q8EvqBqtxX/Nu3JCw1uFGd4TT2p07Inr9KXLjX7i1KqEAex+oebPAgQy2XIpWER+Q+8pZ5i
Ug78GEyuZvFSlCws5qzLGIf70r1m4RfqI1KZGtoSbgzSXe1l6EJimBt4Bc6YH6YSySX093W8l79j
aZdMveanI0o3JPXU3Tq6jtm+71w/55fGkBqNFTY4kJKuX4h1+6AN7M4173aToknGOcSAKPx5k+Q9
uX8uO5WuCb+ICIXauOb5Hinr8Ycw5VNT6AaHGmDPVw0ZNJucB4YD8X06OfSvS26ot1lVeuQEaus+
uTMwDCEwsxc2jsai39P1XQfMqvrbqB4HqmBU9+dscRY0kfc59zZvwFVvrnnFyFXNhaZJ5oFviIjj
v02qsbN5ebLY/LaB5d34EguGMDfWg8jYETDxc81F1jOT4rzwc9p6l6TxzCnikjAqT2oCp5pbcGIg
DqRzrMi7R3g5LfWR+HfHWbMhLR3mEkRVJUrgHeWOZxwVpIvH2zqYL/ZJBviNelWxqACvAWQGucL7
256UdjTCGUSusX7+6yHiD8minv6Uh2KLDFaeSQg/5RjaRiAUeZSJTBC5ch99h0Ym9pe5gykB+xHy
rQRAd8J40hss+WKK13PUtiG+rkWzKqh3JEVFcdChtDS6QJ5OJ55tuAfJRvoWKzRoeRg80nuU1gVE
SSWfVaDaokERugL3pskOXlbv7IBzrN+oZMlRo1OuEaVe89AXoDBsLmhBZFkPpyT1yN29eO2K7G+U
vm4ODXtx8uzbVOSicv9SG6EL8yXR8W7kD3v7qRZXUa0cyLXqpZU7KSRlWucmMkJUP4XO1AdovvRE
Ow2mMLg8tMIZh7TDs5uBZ4Ae/n5njnuJkejVCWSsLEV9cO+MRf+cb4HU+PXyVVsoTue6/TTqItvs
puDPy0jLIH2MFGjiffp9bLk5k468p4WR0Ui2J5DmeNK/nF5oarM/Tul3ZJfN8ijuBsZ+sDuoRprH
UnqD7RDvwHi9sCqSQO9WuqGS2Pk9fRM6lh6CXQZq95sGAfqh2LmXPp6u7gF1ZekMO+bQw1Uf039N
IcCxoORElADlqol4CpCeli/4nu8mJ1hqYPGk6wzRSEDdT6/GooTD7sF5YY9nSi1Vhx37QwlLH5Pv
4mIdXs4UmgeEpEIPnk+T+sYzDZPVPRFuR+HUOsSTKLNDiGEULGgggkDws37lGium5+wJIYCYIxQY
mU8a9tmESGbehmL1XeiPVHnK0xMme5MjRi2wvVJAbzm9LS8l9+5Vvg6Jrs0xjlfjUtjTzFg51cb0
jkA7VHK2Jnp1a29uXBblvwPeJMKRx9UE+zRD0JRlNwr3/i0KZJ8vkNTduoyQyhI17ZBdzqQ4VP/G
JRWgXA9n73lpPOAkvJE+y0x1oMPBguB7ZNmaNxQu+fdUjpx8u3LAQkN4QUDZGijgv38ijDsg+eQW
I1060P3PacXTZZJT3ScCwP3E114n0UIPdP3AT+LD0QTN4vb2jiF1VxhI7SnhBDXjvSI189Slf5RA
yi24DBilyq8lmUfG7PsnYYSuPKnSQWbRxAEi9eJqqIPHZkX1EBIwNI8J2WdMuEjZ1CUTSVvkFHzu
sxb5NuiEku5R4tbtcDR5A4SKXkq6XGnBYL0VIT6TgSJ7AGZ3A+VFD6/7vr8Q5jduieBNsq44qQKH
HjR09ydAM5m5zod9Um8HBwJE4yKwqwJKmWUJg1JWJ+VTlq2Tb9qKgAIfqRw9R2DmWWwloRk7Ppd7
bxYCMMlAt/nIyilsvZ5I115BXgB4CGMTQ+wJ280MryUXc9UcTB9QArFCyAOTBrB9CKTGE8YfiYDN
m4lWD2wyffyiNhdkN//kNa870lqzAh+5mb9xtgh33qiSvjN8yKnUMISlwmWiBCFsGcOc/69JwjJM
OFYbDFssimFT8wzihYBdC4ilFgzkHjpLyNjsWHbjrcF1u565yfnw7Hi/we21q1hX859pQNPqKesh
kFCa+LvCOpLfSnbqAlqIjTX84zFPBYK8crs2RKgv4YlqaLLqQrn8lqvPxeSUP2z6bLSAKJIeANMA
Iii1QYf1A9BSkTrgJipEwF4VTEdcywVBSTnjoVwlPv/wtMmQcBYhpr9BAaUZ9Eij+Hxsol2bZRCa
QD4p1E32SguFw1hIVEJQIuedBr1v46ezMbWd01gyb6Ieu2QdpGuqIiIZG20uNMm1YAf4CrGH+q3d
zF6aQOA4IjwitvCvJVUKGYxusPGS6n27xMH8FQ7VKRXygXqufSjw755ghlxTQlNcxP9G00LfZP+j
qtBB7XVF6Jk2+DFkUwZdMk5/Ywf4Qgp9oI2zFPjhj7pbdsontzzELQVCLT8kok57jZWnHtyCk/9n
a916a9rRtlfB0p5CHQcQq71V1wZhzlSj3rd9hSjeuL22noStDZniMY0z6wOMUJG5wcX8bfFZy8Wk
SCbyFhsjLBFaQj8iRfSfVbMjjXWigsySNcGfR6RBBjAt7A/NBGAUaEYGsQ+U+FFGknej4FmYSQNB
LAgh758ohn3OxOROlCa+GKdda/urkFnJOtpBw0/FQO+r0A7iCR+XgX+y8VqU9+it0yKIOpu+bFN1
vHmHSf1R6Doff1Nc7OPuIv4PegKzsuxA/BT4C62LIOSdnVKGXqfvvnTaX6WMUWKzsp8NvBTHFBbJ
CwWBHpqY9togtSza/iJH+kuHMx9Or7R4CtMpBPuZxEgJHGXwKYGlhjqPxHtY3kMd5nK3y0DksU4r
p+7MvhXKelGKKZAgrygubGB0NF2Wb+ranfAcJe/KF8KUoZBMdULRWyAC5u1KGJL0v78gtHz5/EU4
4tzX1IioZyDmD56T/gJ39joc4a1/fIJGVTjik0SJCLYE2nap4j3Y/Mna2qXBhQu+lFHJ677i4XbR
4d+EBjXSeT4sj9vaB4wnqX/s6y7+1az1g5u2yTydPyL0JkIjyQoWjGPVcPGVB/Y34nMc+msQ0w+f
gsdgIB8UVRMoqz4GUNJioIe9bC3hy7H28gajlyOMJkG4DnWHD7bQKMyZ4f1URY8ahRBXxx93pny2
493wB1ErSmnQ3QhR91il8svG44axoyNDtoz/McD6bhlECkojop0RpPG+mThmxSIQIMpsHDURKo6A
jn+rhj30C6XoSLxAgF2S/nWCnYY9MLPmi1FThxJCWD/uvJ2KrBrQqTMxleM+9+Y/KmmNXqlFiwCP
sBIQp5ZHQfVVJaZ7n1I5gky2skaDeqYEG57H1gUWZtfCjGMqFYQi/tGp4NF3WO+WOE9ULLR380s6
19T2KeP+XKYCQitJiAvsMYCUV80vGCaz/1EL+YbVBj8+WuKpUrI3xx9PzTZrjjYzVzPAV1GlihhF
hDCZfR0Tdw51HJjtGPYN4BjP2l9ko5S7tv+44ZKNEHZOGacf4kSwQZnvJo9+KKI59FNxBvL9lhw1
hf74sZbarcwXLrYRUARvKy+eKhl9idY1m7AQE2E8uOSvjnZdAMNhKqXKfu+SUYcnEvYhadkqSh5F
snOdE8kNXFMDBwv+5hjM2ysAYYyoDvjdFEz63OMAP3bZ/MvhS3f/oKiPCFfOtlKEpDs10Ich3XOM
4ucaJ4J17fkOO/7K0N4Mmv7HtulOpFi7DDK5iVrDgsVf+72PKwVa1polYf3cZnzINbwYEW0j4MKn
b3is31i1bWmIa7OK5oSB0tBaGFw6dLFNH8KpuqsUnVgPQfszgD5ahMnB1YM9JrMyCfgC/go3rzt7
2rB4clGhKfR7DvLApyVGN5JJf8v67nQv5w1Ofz/YCMJk0Pla8U8bYUmfxyE7Fy5AkvfYxZKAtcee
ACifaJ+8sdeVraVUA2WCYemAOcu51j0PlErwrsrvZuEzP3azwcfmgSjHxLS6wVccmO/EDLRaU00m
+i9NfsmMdvoFMEKywnQ8R6pwFjyf0ySgCAOsyM0nKgI62cnMVzs0ork44wb2ste3JvmMmpg1g6XQ
jxqjg/31FNjzEfwsRJmSVz5mpERBh8s21lFKhVwgkfUZh4RZ75cBaGlrxopN/PB8vzcILg2/mC04
LsSm0kGOPQ8J2EKSKl9A3mmpaJ6Zrewhse7j3PUTNd8aZGblyjtd1KzAx1gfNsERwXvpDEE9j7B7
ldsGlZ+wIh81/bqaClzeRL+CtbVGHCUSX7l4OWvBf8oAKs1cLgngbEYOX8QmQ/FRmJ6BA8q4Cm/v
ifjdbn898a2foeJNgedGXpKG9uEgT8pf6GbmIL5hNUYia+43G6HD7m2PdQoSoU903jCVwMo7zt+x
f3Hx8ZOAf1qKKQVx3zr/EDYylgx8z8aZlejo5zABVimqL1uNudhz/NNu/B9sbgMb8XZ6Ia8XSnyZ
OZ5Jnd83czGhwLb2top59azjDH1sGhcl3KJph++LQAQn3UZ4t4oF9WIP5Ol8Tq6DBzxGymLv8XU8
B1UtyY3fWEPb5b4ls1E/5Hg0KQAsQZUrptQCYLjdGRJj11gva3p0SuSdVVaqbw9UiFZT19PFkqUp
rQwfSykjnt9kiyRvBQxfGQGNNfSYncZ3gymnj1LhcOFs8mj9dO57bobcfd7uzi1FVStj4OaE7bKP
3IqdzcA9ffnKhXOWAHrxsUFngzERUFpSLOM0Zp5MmT1XWK70Xep/ZplDpgGDf26zCHgt04i5LJ5h
P0fHkOOC8gMQirYBOUSxKqJUDErL0YGPQ8jAi6PXiDDk8Y3RCa+kyxQX/1w25CR9jEQ/w0gqsd23
PeFxLLYqEw9MJxst7GycNOXtAdy8ZdqVNf2JINRygeiWHc+XmGdghw5E4arRd7LYfDYbuySRi5sa
W3PHVXoi4+ln1OiFV7R+c0egKsHWinHt+iZvT6cyxECxn2w8mKxcfIapiQCFeTbuVPvPo8o286Lf
JmCEyyiICyALnNIRWFxJdQ/ZejqDqR2isIgL+fJmJlwkey/+Fs59+MYcRifKRNkTogg0bHL7uNTu
mXQRGZfaVLK65otMKXz2YN9SCmp3V75hNBzJAS2zF0pk9SRGrQwtlYJJ9vuflj2ZV8tBnG5LCEv/
O4yyR38OyAK/4p/Agffj1/wDDXqJlgzqoa0wJgXXsEJjUQRgDhO5DjgP3lC7VGuG3pcJ8jVULc3b
YoS6HRJVmkL6Z+L95x0OJnVEsTCxSHk9TzNzuO0LOFgql3iIporxks4cOK1gM5ZCiRBs6Qf7ZTYi
jwfcsyXz8BN+eK4VkedGubnVVRpj2od0nCDfJyhhURnSjaiGfSFLTgUx1CBypCl9mkhTGIS6NnOb
cqwrMmB8P0LohD7nFSAKiQznAEymT/0I+hnA1nzPg1ybvsqg1GfrDGd2F0myJd8WVF4pT90RTRib
OkENJs+LfiQEO+eLsXU/u303FyVRZ5Hjy6b2XMU/jfeMX5Y8sDGeBn+iFkttezzpuK6/c+n5B7+M
lmOEQ/73ddq+YBOvDZFPlBLuogJ1y6q+xVSUi1IfvAdVZF4NqXIJ+MK29qAhA8qiqUfRrc3NWyPO
5+IxEwVUFO6WJBrtwmFDt5y2qtxEyHHnY3Z4fKvazFpin+sdQelugYNGk76ZQRjgSPBoIWh02sYC
mk/KIBxnm/SnJMPkaUyhqo3hHPWqEALg31HK+7ZIap0FyWk1lgBPjUluKfh7g0dS2ymy1eQGhCOi
YYwPHmSfroiyXNKkoqqndDNUT0dfJmvYJP6V7zeFc0g0H22sUiy8WQKsXfJUElL9MKJIY9hjOpxq
iO3jxkUJXIJrf5gHI56HuWwd/BgJ66tzj3j6Oicm01j1hvgzQRPclQkLK2WM5SkFaP11+gc8kyTF
BSiHMfA/RLlVUgX4+7pB4Cj0ELf2Vc6S4y4izNOCfdAsQ4zXUsUudKZaR+fN2+IrYig8739wj6ob
dkHV1eGTKPaoXpUsuraNFs3cvap2VOHFh8Zr5CIMq61AEF7mZApmPzbLPAA+tkkLOgWfbd23UJfu
QMYYr1ESSAAOQuAxBGvyHkDLtTYEFmOH87ekaT0dZzexf9f/+pjvBkcD0ajyDNyTyjF48kbd0xxd
vO4bGkI5KvFg4Pmge9T0pjb9hbSu2+XVug4P52x5C9LaoFdryoixosfe7/BzOzYnRr4fOHNofgDk
qKZqZMCMgUzt5oWMb+Mpc4XM0FXjR9EXCS5jONCBHCgNfAJ5JUGp4LMaUCfsXtv4zMXGk2/MffdE
C8Ju0tGasw7MFH4V8AnfBh9Gt0Zw76ZlKFRkqhe2kcAzVqYcAE7rJUHjQ9AyvMy06BpxObWTyZoN
8zC3tO4cYLJkI8ap0t9YvftmJTspvPk4WahT1eEfhbJLnctqU3I8uzsdzTefJt3gbtWid9KtHkMJ
+RECEAky+yLnVcYLB9cdG08hsrAiHo0ed/1arDTYlHbBvgJ+Rynm8dTp/CYr1nHaa8IgQhGk0Bo1
9l5rKjbRL6FVr8yFt+GJD9NEfMdRoglN13RItNuc/ub2ZVLuU2RrdX2d5lkDu3qXf1HrGH45pjdq
RGa7x3fYogR3N/JCkTaWlRMq9E7GLNXwZ9Toob/ajxDSOeuzs+/+0Q3g/CGHdMInWEyCfjyi5Mek
5ZnhDqoRpCZPuVBca9AHQb+2LZyYdFc0FAAR4WyFKQ1k+Qb8DjweuZ4gCMizxRQ4sdj90OG5fLQh
rCzX3kCY1A9Uy0LfFBA94SPL7kACfYN/LRIGifq+quJ7DfoSwvzuQy2N+VJRcc6TGcsjjzfENiT+
UaYHuwD51jb6rBqKtBY9gTQSHWY464BVijp5CH2Wg859a5AdEowz4w4zLjDaQgQxzAUx3KxgE+SK
8l5Njs8uTstlovUDAfuPJQGuC+ZH54hDrkmG+MVFfhyBqqpnfqdctUY4poZjwwQwXPqPNyJVyFYE
nrVSXOkp8xo0Hu9kqlm4B8YhDkVSDEuimPJ9l90BN4nwMbFZwgSDWV9CdK1Kd3aeRg60XUygneNI
Zeof4JPi/8cs0wLYlHeRcd2NxsNFvnefdcW8b4Twp79ZoPWeaf3127NVVnvt81qAVD1puxHwWxu7
+FDf8/T4MQgh6kW/MVdAI5C3yVQYkX+JiDhMBFS6Chx7JYCHD6q6zN8p9TMDkWqo+QcvjUsSABDn
QPdu9YG5zTtGqRO0sBLb6N8Xfx6JbwXNJD4MO4kMWC6H/NUgDj/WYqe8kKXnF2bEAcylQP6bNOpS
5ryIUgLcPCkW6xlwpX9Uwfkh1Xkf2jAGg6jOIwU8OpHU+kR8m1rGEU5l2pW/p1bvim2ensxGEoW3
ebuCQ++iE5cZFJJgii2OymQC4Vxo7eK35o0WKB++nfIOzA09Ji2PYY0R0fcXLEOPsfhY+8elbxR/
XeGI8Fqj7vLkZOQDjYqSRCSI2Z00PqnNyFhdn2Psgv2+tEZgCKAKMftppw18Gl4a40SFKbFVFlXJ
UOJdUu94GKtGZgIIFVhtmkbRc05pwciVqJEzpep4BZltZyL6YuvpdV12U747UBXp8HLdxsicuYFE
aexGKSyVKhrM0ASEjhlWWvledyvlnWlOz8to1QL5lF3wVf4u/d7gMtq8P5Em61iixNQTf3lFknZn
hMAEasJNc3txYPRmZAUoK8jHTqDheQzFuPo+BQmGTw194dhDNf+8nbk0OOvT+cdujiIss65gE4o9
dl7GiG4gNKnMjGFBXv+oImauIOU3dVOb3NbLojXF/0vQ55nJro66x0UeRL3uwBv/gfldEaW2SRK8
Qq1d1TEsy6cBWfDy4IncSFhp2UIet+x5dr6Iwk01LJq+txiEVEOX+YNoFScrObZbDXrzLydQY5PN
ocS+mVnNhiXUNfU8wIQJIBpM3waKA7+jqRsesUfxlz9AbktgQkAJSuqDIfHtm5F/g9e5wV1xfmmo
hscCCQ0DLjcEehvIRN2N4xgL1a4iBdi4FkOS0CKPBVsvCsnyAIWIXB3SDhtMFxfm21QNV6AU2IPh
W9qELrbQ86j8q4pUFGQWXbSbsbFv+7KuDE0RwTrGrvgoHkaGruuDVCCG6MyI9TI/Pfw7i1yaUXHY
/BLj59xeti6IsxQYBpBYbYYSTs/SNEoK2XJ3cDeSLsNPARvz96C9aS6sIKW2UzU8eYU4Ua8j7npf
EEc9gzsQmYhZ1V1SxVcCquPDVzhN9w8NPB6ifjr7L5m51KNo3X4QgU9BFfTi5/oQQZ4UBLmN4PhU
H5/9OPO8L7YFtxI7WgV91m64/tCxacjYGLF7RkcTvWPBFhzU4ndReXIqV3WpXhGHZMZYyhI9PmZo
oehQIKvu23vNmBf1SgIMXdaWsZr386gA5r2GnZix0u+Or7yuX/XcKIGvPHQqd6F5KhotY0d2kHvE
iHm5WiUUQaIrA+VFmdfTXIy9ey3/OA2u4vfoaiOYhS7rPjjQEmK071yiNIm1M79skTK87SpwM4mF
9S1yk30OQGcdURpbINz2f6ZpH6fJYI8IBs6CYAaDI66g8BCVEnSW/bEH0NhxRXMlqS9aMVjUWZ3N
fvrLjui5oqcNFpcFGmzaEoN6eTZLkS93c6UaxZAW1NvUdXeOA5q3iJgCwR9zp2/i+J8U8snx3AdT
P/M/jH5M/L5FTEK9CwahfsMo4jnodFjOZ06uGFH75NwsfebLLq1aot6CeJFBlc/4vNRqw3MrtHZs
jSkxfjt+1R+AdsWgPczzXO3RaKuOJAxCGxmEyqSvRhd+VFIeEshmdvgKiL+WcjLsIjNfsd45UMdP
NMl4i/4e5D5VQEOWX9ttgAjmbwQRTeekjLbkLvVXSuszr7Ic9lK7lK3sOCqOc6XbuHx9bQutvBV/
uKsokyt/+Nf/AOMj2KeR3SYQWQpc4Cj5zmArU0QGM5Pp4hpcfwL0y7yTLzYfKzTBtwstpb9jRpyc
G7Wuez6hgSPNozizJFg70dIbXFDp69mEsx36s6VD19imNCke02GwRHaU+MVRbjPjRQ4CD0HVivqk
TjRI/AZ4jFPoAujPMhR8p89HeoKbjPHwBSh652XtirchU3OgG7obIV01QdrnyApMxyB8Agn/WyxT
cdheaK1Qu5jJiu3puMkesb8yrL7A3nUpvHs6gEhsBce/jx2J4S67SDW027DMat0u8YH898conIDi
tPC7o0THYWJ3DrZaEUgGl0xV0B8y48Djj68+TC7Ac0MssnZ5heTPmi2z47QqpyDSOTYIvhgp9Irg
kvZWOvf81mmvPYAy8BPTJcMZT/goK8nfB92N1kkB5p1hXHb7dGKv+UFBakCyRLm7XbwlHe3dgpC1
JLeuZnWVafwzQM4/PmfL+DEUCeA8uWyFVjojblUGS7GaJSc7r48cdBmUcomfbVyxdwIXyDjR+4pK
XcPwkntFygS5g0UtuQ7rIm3L6p4+DkHBcegJfuQAm/1nw3Nn2Wjlq3RCg8LJDdmEiKM6vAwWR01a
TYyf1JtZNBBLl4XPhFDLav1ko0LQ9s8y8JkxAKxiSIl3Zi5WjtyOjXjXaRSfymQBxx51L5ZC6Nln
2Hg94FcJY6kBuvklijO+pyEZZnLhsJ0/EZR+Zb6msyxZwPhArESoOlDIv5TBvpOI6w0ER+nKCNci
A5+fytrPzQYz06lVqZ7QhhdnXJYALNWg/gY8BDM4chyBa5cSHYQp5XHUKvmLN6gjxshhqaY2S09H
knTwGtsPQmmFQosMV4vZV5DF2iuKPTeOdjbt6wBIiFRZt7DeQy8eJfwLN/jdWsoeidvgLG6uBebc
N2VJFXnw7ZR4dbxQa+w0o85CYCUxmZ1w6vHB0xyR5HbA/QLKom+M3iQjnjhwj/8ApPD1dodBuu+F
JylLliad4f5yel/oSHfvgD6yvVl7VJPaZuYeMog/0j2mE4iTkUEZhIOgaiD5zptJiBLQ5wqwaFBS
WfGxBgYwl36+6LsED62GQj39c3RYtr81QjrTRzJp/EX5BpJ+pPCK/J0tA66fXUY7kahzzGG6R6GY
JzrN9wHxQ637LXwly9GY2SzsbuX0mPo53OafQTzPBWXP74iP1t6+qChAS3Y1GZpzvR2Oo5kys1Aq
3iPZBbbganUNpGrt94JaVTO9VZg8UR4XGRyd8jqku79W5uutBoh4+l3FTIjeZyzZZs546PdXe2J4
xjsRXyyN0of8r6TbQ7PIit3jBmuTviFrb7EGiAIRQOYcywHFF5TGpL0+gsT1ozTgNxChm34ps6M5
qTjcgYDEIOJv76VaunEIiydI/IUD4GUUR4zo5MAZJqQoH5c9C3lgKtShNnDa4KdMLODpsmdGspro
/zU8lQBDLtBXRL47BxXfrkGnPUiQk8XeMyFYMHjDqbdizE2F0haN3jsSO2XBnbZK8yz6LhZ25Laf
FX4C+BLFDU+RQuezIrZ0PaxhdnIFQmQsXtAigGDISjBPWIOsQN/etrQxXLZ3NuVRr526tW+yJ+C5
UPTLsl7jYBV/HafeNDdA1OPzTJCPQhlnhxsW9fG5wxnbjJ95C3/EchxD+1E5GiZXTtKqCd8K8ozc
JBu6AZkRQUlbFV06A619/9l1SLWtqObXjgsXnrpavEMjvU/P8PMYNp1DUdZduvn9w7aTDyMJUEKs
1L11UIsNAzhUGyiCH12B+NEgDxyf5Qb2hVFVQvvquj4J7hnTSjXNXDtOTaVNbi8vA+5nysArhFDe
c/FGHFYSppuQoy2uxXo1LSsyLRgZwBpFW7tue8S5wokVAwsx8rNEwJ/MDUFFAtOPGAsla/f1WcxA
uqOeaJmm+rk1qMITorqUpR2Rl2W9VJozvmMEdCdjznBiPTU+HjxERvpG5SWdQocB9zVbt+UZVlyw
jSCcBRIS8GdcgN7FWEFhppEhBqchmA6YOESQHEXGP5RNzyaN7z/44tuEai7M58qyYMIKpIg/u87H
yw6jq92H0LhVrX8OeJPm7OSIh2l21zM+9ZCaiBootMPxXOJt5rhd9jmdzfKhmyvrxKE7/H8auIQ6
dqyxie+58Qp0fGRbM2poxCQDQ5de1mxs6rZIFlbCox3RuQxdZmZSFD/AfHCtfVBwAtJoqK9YeVBh
KllD8mLd0s+uV3kHyd3+MxjaV0U6xRfnTqZGbf04zdeVSYAWzosxjCnESIArU/QLPiynR2Oq3Uy4
bgoz3RYl4V2fCvS3eS6HIZ0DlOXv01eXsytkHtj5O4jw5F+Kf1OquYzFvFAdSU2NW9QWBrWohvU0
fsXM2XEjsRKXVXCEh2FHlP/XFtJDZ8CGI6XmALW8txBvbOWlnIWRNxVnL0dpcXk8KALjoXvuk8AI
VwKWGL2Or34N/E2UxG9b4tO6xALIzD6kTcNKiyxeb3FeuPkkM+rx8scw5nfyqIzB+t7yQU7X7kNF
NAYamoIXLOcewALjdihb2EH/sXISLfHFYul1l/GAdWsl5NoCF/p8mEYcJaaAZO2ykBH3+CYlQRGM
q7WclnwTKGF0G5LB7hGMj7usMBH0drrEK+1CoyD02DaxJWtE0kvB1HMYEsZrJpvOQznHclNATDnI
aGLe1E6boR9OeAazyRESHfGR5x9pjxTO6N75VeN2uOPV1of/bjehLl2wGwEcin8s6fm6CplMmo90
dBFQlsGuCUO1tWB4a6YVS9DJpWILBA5aMfHJpqHZwYyOX0S1O9lZfGnoCAxHiJT7Kta8PU/gQI25
57jxWgHoyZM2zC08GBPgocanNL25Uuo6FghrJ86uuvRwnmD5FdFBlijCdjW/Zlpod9mlzLmawZDU
z/Yzqp3V+Z6jU5eXRdW9uYc1Ql3McWFZTZjhNxAbiNdsL+Zq9fS1T1Jw5j6y2kjhjwmAAxzW1lOz
4e8q6HIUTislJ9zReNMAZJFFUaBdcxzjgj0Lfd9gA/BkVJLK+LBzujYegblMKZ+PgoGE5xYJ8puO
LLqv5PwaUPJ/9q+ujzfwMk1uLgZ3rDvVqr+vudLbHHn0F7p61oDwWTf1Eu9gVGhPSXF+5EXKFnq7
L7HglqBlrxdaM3Hs2nTUslVZ5dzAQkDWQDzBgdEei2vVbrqnU3Re/IUTxg0OmUvOOtnH+g3D2T+j
rohXnuhZu8Q0rahp9sCr2AiDOLES9LCRRU8ssDOJCo7tpguyGVU7HLSQ4/FgVH1ssENckPOk5EJs
OMmwKkkBf63IjGET5WqTzNNyzq/bcWKlrgB4rV2YuJrSexbY3X4OZ9qYpJ4QHF8+bYM5SRTU3X3P
uoIi27h65BDSPKPFBOHLtRyK+z0Vs+qoqDqAF7X40aMpY2n6RGFHaEERe1bQ7VZSWLow2TShhqsY
Ilod7BPyo2209h6WCViCzFkl+FrBybHpnBkHIQ3vj8hNSAUPqECl5GjYahl4JVyftWWeLf5gY69/
iaTDnmUicLnBB8caIuEvU3XiDnLKvF5F8SIucDw/+zYXgjWRbdULrCCvmC5f9bG1rUFJ/1PJmatC
AY0106S0TWucswZTwccIWg1HlwqfGrPLK4i/Aer7gOcqUpY9wCN7QtR00LYRM54ekc4ge4p6ELlq
h4GOirrMXc/eZFkQXzrfiYjTTZuiBNRbI89X9cImorwRZ8roTVHjymZUNNIycWTnab/gReP/3IEl
dz9XdMSxTF62ozA1kJpNKZUP4G/ZhtnXoICoKSxJt7C1Ba09toLKZ5hA6kWzZFuxX01NVtTUMJd2
493X1V0fBZK+qn7dL27Sf7t+vu9AYoh423kCz4NuxsVJYE4a3OPiBz+m9UFG5YKHkfFKhQg8wihR
bGonZ+km5ZuRs65XQEst6mZe6zdMNtotbIVY7i4isZAdPb75a4P2guESueGKqBw9io9hP/nDZhhJ
gO4+0Kk9Obq/oG8s7jnbSoULGtU3/gpUvOpttxkzb7e7wGMcYqPPt+o9BiDZAByfC8zVlj9hDxBF
DbM4wu8Aez85EQnvj1t7Qn/xiOHHRwX6r6xYB2ASOok1S+8TSFn0xLT+E57PcnakEDtpcXgLFVIM
chb7CfhL7wIxPCWpTpk6icdwxTN2HEGuOvy0Ym/fNVDWdsGfNNga1oPWgMfkYWCU+kOreMVHBOaa
jVaLbCRhuG4YwL5P8h5giCByhiPcoz2I1nGkwKKLU2F+eM8FqpZF9Q9AtmDQRALbomhgMcdRhPpd
1hZr7rJHuFZC9t1axW60uQSaP5ns9vhnwH3hJ3BgfXKqnCyEOpH+qbxh2jTg7EpwQJlYtM2wwHyk
uH7dhuJfqxECQWTIvo1EOqB8dA1drFH8sBt6aJ/bu6pAF7Z67GbOoLADnWcQqRfFy/NOOpDLvIfa
bZM5dFO8cs+28eP4sc57/aUeVJR/RmhY42jJe7RYGgo0Kg4dfJv9L3cWaS5hr0jKGqqrO9mlgkS4
dJaCPC7BZJ04Uy2s3wMQACRHUYVj9xsMHpeTu4n+Fujt+n1+Nci9o9eefoIehos+qrqlFzH5dZbc
EdylKubKK2S7BhFzIgiK+kRdeC+gMwkDlLZiQ1MGEAzVmzGMGzWaqgugoCzHjYWI2djeDn2KjTQ6
OcoYyWytFcEi8g6DByRkWwLrSE0qFVPMdDl6bv0JRCUBTRzTeQjAcziQPoCAZmPl6GAavPLVAf0L
FX1OXIjwotNNWbxiKcmgx/371egWv9ffgpe4MNAKFkbe+envUBtqeR/DLQoSk+wpecGLZNjSKFTs
lAJsetx6sn83NBT+OoYa89dpp0JGGgxMdo0KwFLXXHM1KAI0h5P7xRdLyvaUtPyLN62d1CtgERDa
A9fLvsF2XgwZteRvsOxRfCNAk0chYW7H3Vbiijgzd2cgprU3oTKPQq6M2nW90w2nPtCmxRvS87wf
F4R+qsGC28dLSpkBdd2FONey5Kevylkx9DTzhsJof1wBW+Q6uY2n1N6VxiFkSjFdWGyxQv6Cd55V
sQCVqT772Ux2F3oIT8tW7XXuHjSfQ+IP5GaicsUSuxGhlqFO6gpqnXD7QTEz/4ICBARBTum/EuLZ
gOpxCDXGOOkt198UCXN6SoX/mErofSfL06/1NYk1NhslrzgsGIKJVoBzdQHh0zRQdVG4s5f+iPbI
H3IE4c0UjROhsa+HUQUPTuf7ObC6AMPBa7iIZk2tikAcrsR0l6BkDHBjIOXV9cwLOl0/E5msvcDG
EVUaHWFdqkZeBk6P4lkiRoSiiSAfZf1qDBGXO6HGjVg19nqUyYOAwyZ6/6/rdsb64n+b17TryPhH
l2UNn3tkH/cGrsUD9D35fXmUspEh1ibZUooPD8WgLxqZzm2COEPYIb0usttHCtXdScjkS3Txx/UD
jjUTJ55Lo1IYsQVWBstOJmukQg5qRpL35dkde52oy2Czu3N9gDx1dpPCRKA+ii8rTEtJYqxgYESc
W/lNRtGaIoRKIAga63oINSSIXcohP7DcqpntmxE6nHcnphy9IPEunJngquF2tOmBm0216f11EF4a
zqrs/DLbw6LnJu47mFSqu513q56g6oXjUpMa8yYPf0aeUvFiV/TSMbmt6uy2i4oYZvzEWN5g+qB7
FrWwwX++kHHAfzHeDZFDZ9U308MLLkUBwv7l6W+J/zQnvUPdyukgYtNxYiWJHIB5pcI69ktQRAp4
wWdnD0VN5+bT2xg+vkQoKvBrzU2hy5K/Woy2mR0JEUaxTOgAWvTgCcGlXHE83sq6IOUn74t3xZKX
PLGRA3D5bq5OYHPtIgF8rl8UHR+eBj718BbixQ6q7IhARGJb5BiploeD9VzD9KMlH7aYjSLWwFNG
/coaqjKtpTuIsw9o+hKgztWLq3LOWDy/n0KuiiH5QlXsZnFoQ3aVqlFsfLuCWz+5+hNySjOD6+Bt
QUZsfrJL6f5CchM7zaeGmkTCtIUnCNO4E5oNs74Ra74JOozQ8g5e6SNvTb/Zsfi6kR5SyB5fQRfv
I9znuWjyvbjIAKAslmBYLvnelW2d0P/rAOPxgckibN6LulVqLUWY6ijRLYXa1RfZLSeo6JJpU30C
DQT8pdVZT34R37qIvs0o3b+a+Q9xeMbOV3WgQAKLxvKvctMjBqbP73rq/od0TAP4NIaRhZIDcsh0
96tlPxYlf+akzkqTTj5jbGnpHwKx07JyMUVGMt/z1mtnh3x6JLAxcQpC75tiap2cr6xIrQaGeY2A
OWV/GnHzHbtRIav6r4FujVZQSgZf5D0Z0HWZDOw9X8w29uaN9LHMA+0m2G0IKax1x57knEk7oW7J
AA4lXMpABK2Eqj/J9jsSogHwMvajfJHL6wLnJZtIqA+WsFfGQWDajxJ+ufvEKZGGRoIqNGU9Urpe
THWOLPTLsqbwqL6D5V5MdIHKtdvlHuPQ/mRpC0FBvTlqlZUq5rLMDxtbTsm6a0gFqpGXBh7Mgmg1
YVotWlayE0MRP+UIvuO8oF0WsXGdt04nAjnuaWgvnXd1/tQYRbZyvmHAEZ1HQjaQTKsr63nZ7xBl
FoLq6mKwxYcSY9FQpyhr/Qoyi6MG0eX3a7W8Tu9xZBcwNkl54gVb2aiwrCl+5c9xooj9SSixco7w
O4mUoOFZxzpKhhZgRlaZO2Gnd5417cQ9cBb5qQRHCceyLGz3a/i3/L1joIVgyCvNU7JR8jmuFaui
Kpkr+A6a4FWgvWc8eX4fXWTEthJGhLIZlhLGZHBYKpZLBv5owSbalTY26Jn4KoEAQkjD2rVM7LP8
7N5PTIyfikHQV/vgrzf+M8KwPwpV72U5/JqBdFKHpar9TWOeJ7ffKqvGWezwlPj57VHjXTd0E4j9
7/OuPJfGJsP971DVDbARFtuR7W7x8rxksth/KOEb9QA8xVjlKbVzUeD8JOlS8wsIcULbxwCUpwaD
o4d49YLUqvHqckY4kKRweMHIb0AxsBcICVCSgWUzLbxSQNW5yj/jfbe6vP6gXhjYML+VGt03DVyb
etAQeDTqC11FNiJSBLVF+umylKJeFh0Tpp5uiFCKWnc22V9zE7Z7T5k8orRROMoBYkmjD4U8WKjT
U6DxQhRmGyiIy5v7YOX+Y1nn0DEAg0f+A9pM1S8qz1HCtocTV6fAiGm41Kec3bevfLABy3eGnVZH
Z76lCKl/wTKLvMNPRwZRJp9yzrAc9At0yYUM8aGyMveSfMvpckJvvyKet83yxfIEUXav2XxkyF0P
t15c64TFKCa2jn56t6/JQ4tGSCoflQ1umTgrhnGmGUlheVwITwgMig6Yw7cdFxu39ExhepZ8EBv6
a/a9FI6NHVEVDPNn35qYHfY503vjuBHPyUfh7yZGRzOD9QsSoVTPEcV4SBAXWVdLWSuk3KzdAmG8
ArzSh72ZlAGdXTRAknshtBj4apqSI0Xs4t2G37JCoVzXT3kBT16PnG7KHBxvfGAz45li9fdn1UWY
98nwlybP/gvVAu7IeAZnfZLCbJKDDx9/dKajdxf07liB9mrc6W7KVQ+o7Hlv59HIL1QyZT5HZTQK
SBK4ZN+yCKe1ucdNUretpIPbZUSj4FGwPRhrMvZwj6K0EAZXdUzmrgcqHahUMUVTC7i7nroX8pdH
DYtV5Q+kyC3ZYmhAOPMvC3KV3t339zUTmBTRUxU4Ew/deRwlnghe3WQ3g/3vemq1FDrVRsxhXOCV
q0VFkfkOqRnyMSTEDL08E/o3SAZMgjDS8wniyNN50H1t9Qie1B2PDxTPg8lCYRlWYkOEuZ9wWvI0
BRGO7h6fEXIacnAOz0gN6OBwjCzI9jbVfKHbFsUd/nJQASmaWGfzjI4HDeFBrqaRmyf/xvhFlCen
5XUGThtHQQvk2VMskHNoFdVcU+hbLgzYeERTh44EO8V7Gmv9OJJsSqyypEkV3j/aW0XDJ9Ss933D
X9CJwyvS3YZtyhr5aQZ+vVIujhjKx17S/N1Uuj8T9aZPEmy0JFXr4P+mM+fRz3bQl2TPbQc+utSb
qVofdMe/HnUW37ZThpj/YXEyFSnJaxaLXSyxatEOjWNic8gY92ioUK041mOepvzeowKQdwo4Wkkm
hk1Rj1d3UcYt6B/nSHSITPHoOKrhQtIMUFLgr1FdBcKooDefFBrK9hou+p3/hF+c2lZYqM+9ZQvd
8jpgY+k0vymCTu2QgmxR4o7DCgBTBeRWp2qyEcfeSghvt/r6tMnj0qjqoI9tsxxKHYytJ5GbI1GH
NQ7B59TaqDnLd4UHil6YsFspw5IJ4gRMqAy3cvtX0XcEptuKCcrDFfBGymdqnNtd30reWtuyPJQD
aBDWHEyLbsy+vt5fcY5mLaOwRSRe42kBtFit1wxsWal7/Thn/nG/j+0H448QO2m2padqZSusq7B8
Pslz/+JVok0pyiAzzN4q/P1srhMiUWtrPsuwr05UcdQiVqTT239ls7y/S+8SBr2UGwR6H00WJJ54
xcKyDcQazb31236JCpAX0oXkBSubJXuJRxcBLrmuLS91zh7jGLWcqDh1w+8xi1KxX8D8HrVbwwdo
h+bsG6CFLCE7Sm7UxBz0X9jx7S58eU9btHPdsOds+0Qr7CZ3jxzlD1iTUdwlCR4fN4SGDh91EP8k
gGqUNGQFQaM8v/Gm5zikHLscIBg6MVVxZCJn0qvAisBiU+yiw9uuugfBstfIANwrBzkigqz5iO+p
OeOfIk55TNFUXP8Q4OPTF3tZzQKUrEzFJv6y4uobWJna+gEk7kOllBdh9u9Zoz6foGKB9d9HvtJX
J4VtrfAWTXfcSVRhK/Lk62FkZ6dOHX21TCYdXrGJWylf0JTy9MPTS91wAepfpJKeRMxqK+RHD5iW
0RI1sEbVrbpGZNiZVzj9MCb1OmvehGcT6AemQQQkhGwmWl7efC/HR53UeE7WwLjiBTFKhWj/+GUj
vBW5c7AoxgNCIKtvha7gAPgqbJu7XpUdqbYajYAwI5bwlc0S01EZ6efdlBSM78uGyWcPxXUqPnNv
QvYXtu+6aN4J4ag+aY7XtVk0PhjxzlVCbYJ/cmTo9F3KLJ2ydCEea/x79xH59tJNkvxL1jWfmSqx
mOdw8DAKoKxao7z+W5tBAX3+FfhcU6Ye3qjwBxpjeUL4uHHFGkVJbEdDEE8BS+9Q4yKatmkrDFi5
/qANcaY+qvcu6GtbGJLU3nz6jCst6LnayRhGscnKHgwMEloH8m/qM7EzL4sPnlei31Fxk0rbNR57
MCoTX79nc7Hqx5AEFfB50BkSVDqZ0aB9FIIs+S1xg8oiktjTQiYXet+H5SbGQXu6JEqqA4iT8lv7
g3YmP05n3qJ2csWCA6MqMmaawZ7Be4ZosJVpocF+OAvjxrWhjsIv1SX5N8BWmQyQOXVhscnWYzNi
ZA5FoblxcvJg65ssru9jMKe8Mms6CVR01FjeS4QhcngIbj7DkZ8oW9Ag89KKtLJuSSH3C5u/oCqi
RmoTIHMdNcCdHgSFWrH6XhgikAaDhkOdlqd0lm2cJQzmLZuF9vFZTQhZT6NYt59bTPoilj3zse29
PTQoNKmeVl+pWZddUn7ZJ8leOlfRxgdBLfD+QgldCNzQwnVgSo2bsW8ubdiEKAmQLyb/Rn0vwOVE
u/97OP+PuDdhMH19mbaTFDI9dl/k79eqrvsad9ixV0tq52wzub0rKjSJY0uEclxXAzI36bTnQvE0
m1v7ZpmAh3USo1D5FoS4ywsTsxEcypM1nnhFL83BiHhO53quwsujJDizu4pIgm0Ls1ErrKkzsVRr
C+g6YGlv6yCUEbmQXghQS3S9iVC/mqb8SSlQiZECuWhe/dGFbLxQ9WFDuYacYtjfPsuY9yhyqXGl
AtliLKjRXv/fxW4DaVPKDshfioGavn9LldtihHOY3sUumOzXzdHeYRNbVkrekmdJCgAXddXRS3JN
MbSUL3hF4NtdfFYhAsz4Pgy2kCyXkMhl4z0Zd/DPaqXNnSsQ1a0o6NmRQeHoZBWhnbEuLd7b6QGK
k4Rpf3g34JR49Ggkqyj+FSvk+RAGm5yRafcKkiLIdgLm96a98kThQvqq0JBcx8zBzjT5s2W8OqlO
FQRQxyeozQrUrRIw8bwqokKmqMR13kgwqCAndc8RGoSzdiRHGqFl5ZiHuDNtFvi1tYWxSSiZEQkr
1kDlRlLBr37jZtVSghu2sUNs/ZDCHcdlmBCAzqNCZGGR5XSiTCHLO6FMqiHJ0ae4JWMKXVXqXNxU
PjASsjL7bjrhm6Jyg/5spaUF3cu9wURLSPc+pMwVDykgi5ZIOlvNp+E3pAYYAUQSRLHOopDwKkKJ
5cEbLu/Q+86NTUJ6SixSv3dKT1nq3Q4WLbrgcx6FUmfj9ZCBBIsy5YSLT4zY/pazuPk50NZ8PCFo
xD0u0UzXSPAnhaBdBOXGzWJTk1IYk7FZdTX7URN5vSjBOVYfzcj+g9Ne3PipVBjWyrnspTCkPhz5
8weZRTb/dumDyIXs+BzXRVECUAu2KrfAE0V86O05T+aqSDKozOMNWuz6EM03YoehmeDNAhOVLJZo
bH9YwiiuPjcfkWvKrXweHcSnAhBDco/PBR3Y+RAsI05h8sKgylpdjMMHHW6FRWqVfMn9bB5x3Te+
HkYhwG7OF3re/huaQwnd9qD1lWvt8Tr40ooasJuNNKnEYCO/XxAFcB5R+XQCX7P4wQIlGP6/xswe
kI8LblULyhWyEEgPBXiSe/qwWAvs66QoD15AWHKSZnldx906GnYa/PZlW42CizIX+RRPHNimWAKC
PxgjYKlcyysjP43IBj0tTBNyAE4jh35OxqVYXcGWZzuFiiLk+3kAJco5cGB51E5aIgNm0+BU1VnR
vhPlxD5CCVTk9N7O0wZ2Yrrpa/Qy1RaZWCd3mD47l+EUchi+TBlINbYxm2GsX6U4eXHpoeOg+Srk
FJd6qLD/fSX8aS3GHgdAbD0HjNPqZ89+qmegFum+Ec52/bAw/7iYNjBx9HzATdBICT3kycgWVR9g
lCkpZ/oP447L7ORJUNz0xmA1+g9OKaYnSyzQ7cuUHdvgRstOCvoNoOTeRla77ckSYgAgifhP40Qv
KmKUYe0eOAU7uyYpqHgoYE23b5V05SdfU8T5vki23nXx6wT/3HrtsVnhsSb61BUbUjwBljxuIIY1
iAbzkqiyrIprwzEQAVi+PRhFbwRlW574aPumeuQCouCjNAdRYkDchgLZ7apZwa8CxfAskJD1fuuF
CiSIVc+gk+sVB9Ss44uFh5yTfVshNGiT9zuf5kFGM4IqG3rtbAgEOY676ZIkPJbNFbbwUBdKMsCT
ONgc6R2WS6a3Mhp/wAyT6SQZWEVj960Aj6xVLnOhFWvpykIde47ZhrI0ndvhaysvoTuidq0VRJZF
rgC12Lmq1KBdp6rTaCQoaAjTOHmBUBIY1uzhAcvCNTAHPOqtWVZDJldQCxSPd6wRWebR8cC+CWEA
45HUVPPW5RFxbAc0hZLOVuAVPu/9TOKVDT/vi6q+lpJY6AqCXtSHnFXwGru23cXP6vYKdh0hQwdi
MG9MqypAM451YEe5L9JY9H6Bp+6qvqXxN+tJQbn8lQ5/t/5mElEr1FU/cXJ+ANxveBMrA/2/OkAq
CLFY0WiUD0jjlCN7CpcGD7DWRX04s8nVmM3WhQu3I7ZWuNvNEcb258iuY1ZcPdV6xdMwSQShfDWn
r6LikLz0xEOKxMac8y1IaG56mg496FJay1XeABYJX4LL4K86uUdiD4GxGQEFCBIPxxvXv+canp+q
wbyTAbsXFCwQiNLfWev/aEaySm0dmEnKkGChT7RH+HJODRuNqrjg8fcgb8GI79xAL+TaQkCqj1Dh
KkDFIEO93QQwLCmXPDZgpEssUzbQa1QZV3fobD1ylCqts5xI4VbGj+oRh+oivvIjobqtRjMIObUc
XzUCRe/qxEdtW2H4HT52IYBnAEr3ildU+4xdN84/YtH/4F4aDdbWdkyA+l1iXTA9qWXekvfJqZcW
74kRgjTfXLKINJcPNJYdDjFexM7IV99vT5ER2lUzluAK3X3oQnBm+re4dUJ2QpZ9dL2roLaFgWJM
iLJ3TkaxSQaa8ODj2CVYnM33Szc2ZwTL076C0XF3T6ZuBVynkGBKoGz03dJ4gwIHHPeu+0271kAO
RfCRKIorud3v5VHEZd7Wm+5CX1WPwGpSzeLK5loDeNnIP4lFiWoJXbJL+Vs+hLR2NsTFRPJstD46
4BZgCDHG6nu5NUD78ktCaR/FDbmlg8haazo8xxVZyYBbTBtIEEYJGdC4r9bniqzP+Z4L2fGY+HWl
kW1ilxwwgklLaHTy48aNN8Si2ze2SA5TkqHxoEdpS0uqxurxhYP2ltl0KrqYeNu16DzJ8Oi/sCQZ
VLnnNqEte1o/YlvmbCBeSfxHlqSNc8ew0ThMUiEKCla1kPT37kJHaPI9+iCQuFaqc7XT9CBqz693
6+i//H0GN4/7FDic3JdugftmE3gkmFBaeXat0WR2Iazm9rGGtD+REpHVwBJXRcngUNxG5n8vC9iV
X1J0uUpcwmHU0jH/fYUK8q/ooVKeEO1WKm/k3JekFrBwoL9bK3nfIfjgOwAq64SrJDvxQ3ikiuaS
OnnobnifUyazp/WhvBfKu3OqVTi8A9EAxmCU9F1Cw2nj1qmnokRGoJU5kgRo8DO8UmT2c8EpzJBk
lrp1WhZ9Fo8Hum5RwuuvsMh0y/s+y+U4+O1ddC37CoWBdoowtWFPq4unbvJo0x7xEVXep0qo8kE5
+nMcpds81CxxPtNayJJ/eU0FaPbQh3mcRWx8qyiidfWXCvcPLXAQVUEPUJf/6P6znqgexu0DZ9Zk
qSQXxXm0He43wycY+xHFjONncss16TClv3Im4Xo2Mb5LXbjKGXwC4dOPnXQ6PB9PIX6rK4AQKjHN
FjyMxYAgXAuvHid8fYZ1tjGuEcLXJyJm9GHNeJ0+UXo9zhiZmfMp4yHwQG9eno+WKF0l9TzzLA/c
V5Zuhnl7JtQACZerDtyYlmb/AAa/u/AvFzrPNxMoK5Xgn6N/UjWrNHQzDuRWXtvZxEnlQDwpD3gL
UdO9cEddUb8F+HEBJrCiaqvqKkgiLMc9QfvycckPkJtgg/aKiwghpgrLboIC/iL4kM31WjK7rRIb
WIXt2YArv35WRf5jyaV3Au5ctnxnniCjJX4napGikSsRDPLMllEAUIEWSgNnVinR+8cwTrA/5lx1
UdY/WtusxvpPaOiv/bztBM6/Sr9nkhxxJOBS6+jzaRlBXmtPF+Pwx/vj7gH8AJMtsGAh8U09uU24
s8pCmmn7DM9JmegHlFTyoOyl2VBM2jBAH0vd8gKkzvTZp+PTqmql/CCBqi8nHUJbnN08jm6Rl4Go
Qb8g7UO+OQZmvVmk4e9aTeKipYFB8KffJIwzO3RHB2it0P2Chh8CCGGTmWSbmgZ6W1mIObkYtv+O
OXwYy5+nh5/hxPxDbdvWKorm/WFG5o3RNww/yMn/F2osicmwtXCfCel7zVT5gtvaIjW36j4R8D2v
tHAz/XeAF02zSy5wolgxNqXZFI00eLmelRhpigfgmOs6bzMJbHfaBGPe+tuI8zfpd8eJNZegV5qq
tUGM+9AzplL0E/078CDzB760ENBazMe3loycsAJmLj8sTMcL3Oo4WuAzJIio/hYTC1oHlNiskzYt
KjccV+MoCcACRZgoHF7qIQ3rr+BeNb0auWmFZNi9n5YOii39wlzOBuUqzE9qV4hDU9lKQ14jzD5h
kzC0/y8/Xe9k60rmHmx+GUmUIbgBkg85cmXG4umUL/hcXHXZzXk/v9I4Oi0p2B3HiJ2a+WaNxk1U
d1MUHsFY+clfjY9UC6eIMJab0aVS4LSYtAALSicRUDDDws3mUOyyOHG2qNSUsLoMyrSUArBO2yfV
Mn1H0abipnhy/kWcFbAYlV51eq85Cpv7f30yaxDb9MFtNYwAGH80SMsMdnAr/U9nD5JYzZ8oLewc
3FPZzvGH/nAP7PMOA34SxpBj87CQnb5hqRADW7TtC2R7cZ4g5pf+e3MvjfCQ97z9yfn2SArX2xs0
j/7me8ATE6UjlncPdYvRr3CuT7mN28JP9123wuN3OVAz/WRGEbjBWVDnx3QVpCqrnD67nMv5wI7V
SqoRL1FRdfLny1Xz0zmnDe0n4Zwtnr/QsBH91v6Kaebci+yQbBzR2cGyR+2eGkg5AM4cimiV8bU9
rov/ihVyllsAANuZGTrpoZ5k/kl0pJsuuY6Go0vnYMhBexim35sHuc+PYYEAec9NO6ARlir8kxhi
yE9mSmqfhF9w4/x20Iq77fZF8Jpa56DqLnOmcr4MTFh5qBy/eyYzuNEziBq7WOD0p4WOoYuQpPbW
74U+ctANqcNnj/0OBwAX+crxObkN3HxKNEVOoyrHUQoSJLDIQCk6s+V1vJjM9SbDQs72iSpJC8r4
/ra45TZZT0j/MfAP12td273KLhLoNI+QxUJAJxG/ZAaFdqKx9gYYZxNVNfN+krdRRz2R6f0WupY1
QCs3e4lhQ8JZLvBOV3YMoi/ixaQyENqLYPwEDzTXz5LS6CKKMbphF0rHkxsmeJ3S9DrCpQqjWK8x
cuUXlXhZhSPc4noGwO510DzaQrPTvR3ESdWm846mR2FPskLbvbwzi7E9leQwDfEjHIiZLsmqyUV0
24osuG5Gc85spVNipOBG0JJDTQVjYf/6t+JdKp9aOPlGkNuQpQtl4PHZXtknVqL/x6x73Vn2buPV
lNa1qFZEwBBtk4iA9OlPTE28K1lxh1/ManOoWzLJqEeEXrOlHUah3lBiH9QMhgPuuHegFhv+Vsax
hm0kQPJoEOKoYPeIWGwjj/GEztJ2DJwiviniAy+W2DXrkPjIJlSPQ3Jvm0mkpy1lISlZwS0yfMSs
DF1vl1rLlNCzpDYqioEb1a/+qOf3z8NPIg2edKC87++X7ZJGaFWSFzhzJx6OBAftYyKnQKrF2D6l
Sl1/1ifgtWuMlS3JfJPSC2zHuPLXolR8OzEUTzaNGIa95o+M2GdMFpemZsymBoovjo+3xzXXCHvs
3CB58LsXQvp5fpwCYFjERygbNYVeaIZyajUGhPdZx3va+O5R1w/BMq4Gf5b87wcH2BqJDLEnnHaj
0LpKGiIxX52EAcQqUdbjgaQ7m68DNKqIOUDdDLSJAGtTpRJNrSp/ggH3wtLHZLvdIIFRTCvWDtdE
10YUlkcAAQLLCoVDW5JPbf9W0v6F+3JFi6YgG3bA7Ura6rkxBcbC4nLtAxM64JYQubbqZ38p4vwe
N2uBrADrqIb13UO3SVUxvPMXu8yOlAOy/w2OokzcJk3Q8hZ7irdJ00AV8rqBV/Q8lm8EOGkQibrn
M7g7aPz7wKy8/N5PHFaslFSkT09PYKeeYHO+6efxSb+OlgZUsNwGaPmQhZBYEXdGye83xbAaziz5
tKrbkEgJ76+5mzMHGZFIRzmEE5gKuXXmFmarsJGnV5VfvBNglI7bGL/6rTk/jGF2CVyYGt1B+vOe
Xh8MThKCDqKi61p41FHevUdmOyTT3Yohxn8uEamwk/jA+I/5XCBFts5RH+XLND85zwOFwkho07PM
zyRXSQgNar+KaAmkxgrZWoxcLf52c09spMknSxYuNxspn0p4JjH4mUf0u6dGTep287Hc+uH7Rj3q
X7sccp9nuT43LimjIzUbPUM6EGKgc8mhTQDoJWT7g1y4zo6ClS3r/GcJ3+1/jONHROlukxEKTQH7
UQjfKckrHjZJSqJZ8se9swmS5uf3fm0GIJaW/FYuhrm2gG6ryPco8tPNz9m3cwoBdviGTNBol0mz
dkHG7ZuSQWKzLKcKLERaPi+vv2UwMN76ECxQC2d2pJEd7Nii3r/IOIPTwd2WgWuKxtNA4ASed4DT
3lBIqdzg5UlBG+2CtizSaAFkrcjMwS66S0mAQn1Nrvg9d+ytlgZKkb+U98dS1kaEjnAPI2TnaMiS
liE7QZeI6rALhMPkOdUrOdI8LTDT30/7mQJ20OZL1bHceSzSwWmAVl9eS6Bdsh3HHozhGSS0amRU
ovPulfexwpWf8YV3LW+oej/JS1yDXpq6ytDRgxl/7Fc5i5kAKA1+GyvcXjKRn7I3fcQ/C0Cy8wBV
qsLz1eYBaBJPaOhDX1GF0CPqCq05OHhuiBln4MhQJMWQ0tD31ipOcnHM4daZt4sVTTgJ7UMm1yZU
X5UfO5tOoa/H/xJDNP8orjvz9qCPDZ0Jwwb9WzAZ7FvGCYgRZC42n4dgXKw59DDFvIxzSyh5h+0T
bGYBqsW938+fF7gx/9P7srmQj6KiLLCcgsrtXiC/9bYDuEGAdeCAyf263pKzUHkgM4MM1bo0fZme
6pCbUa7ZxQ5TUkWhH2F8/HDbsKm8ISxAkTUOuZVCFibVE2KvDLpCCjUaDae13/Be871EOzu2nTnB
h8WfKq8at6sqXEvPAqjmE9ZBmKLSLVzrAkUhr1h5OAA3093IXsTU64PscbUD87A3tGfExf+bYvVp
1NNmD8xJ2LmRYoJVzx89kMGsaXn9suMe9RsvUQb/QVDn6bQ6skh28/9Y8Ch15iBrfiL/UspYbrP9
rCT5owOfqa6IevcWldC4WBYobG4xIc/WTpwVZwMhJAIrHcCKVq5ulcTKdgDHrhiWRy/4yliODOk6
LkvcNw2Ui8iI00UjCxdnXPe1zBTtzx5r7yYDGaoNV8dI2X87m2GyD+iFgrO2zDgIZyD37XT21MKk
tiIl5qmIswvfGV57qLpfswleH0Ng4JTvNuQ1VaHIq7+GN3HXm5y6ltO9BRrp/NHTqLd8/BewEMTD
1u8uvjbQr+iH1d4OSQDQCQ/rSvn/pKhdE4ef+Rd/5hsLcZMb3ckIBMYypABCElCo4R6zlksPoOjO
kB9gcHtgLEAcJTjFlr8zKubf6j32EDKzZgXzbh5eWX9Byv8DaCfDc4YowM5QYyW5j9/Q4zNG6KVs
6CLEwq0zXpy8OTFXZgyNzZlN4/yJi8RfyDiO+bzhEPi7iSp8bTPMvPxU8OOjjO9pHGgRwYhHnZLX
DCevh44b5+BBOlRgaQG4atJ67kQyhERsYW2X2KzaPKbGpIRBMFZtRyi4F9xLVF95L+QChyjT9mUt
0Fgwghl8X0QDnJ/FNhd/e7KKpT//E1foKUXyz1A6Cw7237G/OT79WTdbKTwOLkbdVnmVrnqNtVuo
lRYYiclwRrADJ0FgiEKMgwAM/pqaDT14pYVGfewx00Hi0IRoCk0t36+7CVO9QuDtZXKY1t2oddUl
M8QQTU2GZ7G1wgJFrHRj0hflBp9LH2C5wMmOTrRpRrNSAkuEph1DPWREpjR0MjShKwGPhPRNsYvp
96VVEDg7s8TavMsYXtPjNl5YLk2oVMzqd+HC2r9UespDCc80fwiarlopqVGHJxAIiHkSTHdNspTw
YG/65WUhTkbr5YyQ9Qu0+k49dv4U5ySPErvOdVWJ8aEszcq+gF3R6oI9gCRLm49yPg9aN5aI5rNS
+enSMoj+aZ2s8CqceC3czKlV8IH9vHI71TBsPryEnu2yXBVZDRQuz7ad3P+zwwTxU7GAQqlyA1ip
2vG5MiP4v5hy9EJ85iUijGSneXW84EAGHpOR0bs3lid8+JQi4D9iouiBCT7xK4WoJZYCfaoG7NGL
sJMNhfMrAxjk4zU06DvZbby7kQTEMK3raCN6MID6bI9/v2r5vYgNjucR8FZSQy04IdX+OWFBPRg+
Dg9RoI2bMsLmboayuLOW8GqS2vHjALc6BvtzPjNxpM8/sMNw+2nwM0BWS7eqNcFT+Pqxs38jRLaL
337T0TNFMlPN7UkbcdbsH7miQny6E8XJOM5dhA4xBZCrDDwVkOtsDIoZUSxxLg+zWaiFU/9o6JDQ
drjMk/VZq1sOCqR1OA+EaW3hZgEtJOdACxV8Qy0cROGaZXSNywyVIQo2r5fM9QbDwKBRqfk8jrsL
KEqObr3I3TTbH9/x7FIpFKQ1xFzoBGhnzKAYn3ou0IOC566PUQX2OfY05TGhj6YdmYzCr5yexcqD
cyFeuxuDRi7OpgIt7Tm0KG3mMWUnY1gT52cLNv3CrfRLGcoIhpIuAxQ5mm6QAHX71aU5OxleXbif
M47fogkAG72PXrq5oL+8rFfVpnGFG4TUARnQFcjl751BtfNXonUIssTSfKQnrq+wdbfy5CToMapl
ToZ0KqblHusi1S5WFhWvb3k6yth1IP3uluh6eqFwTuRh0g1YvpSwt20dQwLMBWRNh6EtvF2OuCij
bwYYHed3oVUPs2Cp/d3crx9XwJ4z2izmN5OSmzqaVglE2blmWPXNAgHdtCMyQ3TIas/uIDRmCoMS
sDvfPHneRDE7UWdr6UhwhZ5ha7Sozqznm5FqeZ796LiFEzxCb3Sbf9GjLYaVKWMhJ6vpJFkI8FXu
uwjMQ0WYj9B8DnqMfZLq0LgSn3Ax8RV/Ns/9wXJdsoVoX2zX/OUl2pCkIFwhRv5Izh58Ybwa+yqh
naOHhkDe55Ys1oZMKEu1h925XotRki/k/YexL5aZ/oAcSl19FCEY8wlzHs0nHF2USqWHY2Ow8OxV
hgsgQJABEeNUNw/k9srM2mPwAhv0Tb/D1PKwEPeddX5Y1bzlrsNaHZRpjpzqvCuLquGZMNSIRN68
+clPmjPB3blq1/WbElUfg7n7BTJOk+Ivry3tVOqPOfPUxTKDayrzkOvDQFvViVhuHBhnULb2WxZ5
2JyGd1KLsYlb4ilfPW5gX5mLWyX8P5EH826CKoVq16+9h90BSZszZ+2do4oiMHoM/1dzsbd5zwK7
glS24vPtBmlODiGIhks8MhfA8mEJDiLBt5po/5F7hUun0hXkur/eQK58PdTULZcfz3fzYSoRZ4Q3
eniokHgcTkb+5XrV4PmOpYjpqtd9RKIbkUjoui9FmpX/+lnJQvUgW7fopyucbFqhxVTU4EHZBVMF
9mt3+SlHVsIek1xPW67pPIL9V1B9EKYbWZGSPUXtbDwNT/t+aXBfDIY9aftOtGauIkPAaICkJpXF
YYJ4AzcSFkbUihvPtUSo2nCdT+nfY1tUfEm4RqUW6DANwYiyAa3NALuHdokYtf93iwPDpjMxhj9d
lhZ+m9ws5J+5IHMLLg9qGzbl4drrdAxavl8jISxMSevrz7Mj7mLKiqUM9qgy0e1dSfxcxYpOIVBx
ouhg8V37QSa6YZR5a6s6ykmbK4l1toJ4gM5C9WSpcul5VjpFABqUizZmo2MAXnNH2No5lP4htykb
3q97Gkuma2NqLUo4gCdbWtVyuwpeUU59aurwTgTZ8jDq+7DunBC0rnJp2/I3OUKWdqHtbsAH4LZy
6PLvuXEG0VBiDJEvsv4rYK45iF6LQw70U3snBW/FbllSVBNfJxW+caYY5nIu70+VJM0SNAj+xr+y
ImKyXEMBG7WwPT6SjvhF0Fgl9nwrYS0iAp8IUJP7JWSIT+W5u86Tmjjv9odEaH96638jPc4/p4hJ
pYpOIeOHhiT9lIj7Kx6sXXdbvO2IJe6C9Nu6KlMy1e1pk6ZyDDjRiWNZZa+S124SsX9CWCodnUbb
89MX1FfW9ihdicJBwTHDlS5mPK1yspZ7rsnA0Hdv09kjNMliI8yjrjjhPSG5i+Ab9OtAy2jBWaUo
u1rRm8pM+nOezfqM2ND6Th3ZXulM+IQnCxNkJAtSlq4GSiMe1dUFWAjVv5zZzJtHEAfTj9CQc5j7
Y5xL7SigPDg0/klQVm+n94tO3fGAZ6ke7zcYTQpyzBlNrC2hIeANrmeXUAAx0EcAxBcDxjnypklJ
yv+3Hzp7RKHHcLyXH2uYsJBsPdQtR8NcT1XwcnhiqyEFAtkMZy5nvYmY9aG2e+NM9NfaeBqGyETb
FqCNzk8lrVkASamvURjjvFun0SfsLoa6AHCKOPm+BQl0GXPVflzvrQMyo2Is4wpSv5ZC3MiWppy6
F1W817h4VHydMsqaRZeI8FC47xhlLHPwUY4MdfSmcFRVNpc9lHbsySA2KnDn+9blfKSd8RFqdGmM
FGIUFLqnKEFOy+FzLLqEQWQbZcx5iDLZknpqA2hdXLlYcI72Yof53BUUhCob4LODhtkDv2SEDTzY
xt4KAKdgOwOi7UEWU9ncY4lRpOms/LGegjLbXWjufWDm/znNd9Em8QIp5AuoxPc7wv31gl35QDRA
tIBMrdjpRVOVcb7PZUZrWJxHJYLCl8uZSjPJNVDEf9MhcO32k6bWMj/OYOaxWHwixjMUCaNemwLM
Z2ImPJoLZHV1Lfr0IdQ6PbzVhL02npON92GDk94qeFnH3FPBA3zLimc4cYGp2Dh7px9w6xJfjJ4G
Fx2Ybrgih6b7yJHAhj2+TeIpChB4I0u19tF0/8R/bdm4UAXw4yHya1lbX8hAMRb7APJjo66GE1Cf
IewaF1aDL9pLBvkzN706kkDJBLLI5vomO//awLYonBJ2jWfo7IADBgba0zrpYym0vj6tRpO+zVzQ
9IX5OjZsgs26ek4MxP9RDOkCxlL+8d9gm7tBA57DCmDOjcCrugSJzJbd/NEPegnrzo0OjKvZDnb4
+gEXMPv3vntFAeWzKpruGe8xyT+s7gxXqnZkcK0+jXkO7F/KLRZcKASWVwOyHUTs9Jt4rbdCKh9H
owlKN2QKaZ9AsqfVPK5LElwzuzgDvkAyhOnUnxbS2zuELA5Q/RdTD/yziziS6IvrFbVPyznFMgTF
8hLFQvewXTnMBnYhUZlC0qDZyVIwUm774yKgs5JSuneqaKG9YBbDx5sgpqs06HXBUo3UmDwVANZn
cso28lwhpBZr4R+LH2ctC2OZDL1EybcbMfcKx71wInu+5iG/gP+/nyyvmRFSGAIJQ2fuJEs9gkyG
Ph2aO7NBdvaBetUNuCivepyPy3bDbkq8Ma/Lr+RBc+f9i38KNYAa5a5s2eBdxYIGfJ37RxNnLJjh
SbhVV7qX2X5DHNAxlNdPfQqWTeyYDBqwzYmpmx8AN+o63e/RxTHHPWI1nhhd8ie44VDgeYclQ+V5
B8aKMf2UYkqk6+I2mjez9WIyb+id6UPvRMIggAOnzhpC1qR4s0NnzIyUiMt4Go2g7venhQFXPU3W
BI0278G5RmzS0TOhgKMKxuocHLIUI4M8HriwmBQxYI4HnfrfBms2qfnkT1WnCN/sdHfP2Gkwt+6M
ECMmekbz77tCVvRLGw/NwXCFVnsu4M/UIf5FR+hvJJiTdlWcqyz8m3OVoRzo7wfPqyIGnVVzFb0K
/FZn/Hr4TcoHCgXwOTIMP9ykmKJXxtvP6Y54M/oNDKFuXnnYJvVnHLj2NRF+FK55F0KEx647HU3a
YtEwQmPHASZ0afKwnpqB+NQhIacrlCKMcQU524BDMD/b8XeS07nA2itVLzFjsjFMocsw5zxPhWZ6
jxXjBom//icsSuHRHzTePoEFb+gQrTHAMSXRr/CExCdKPcNBMZ0Ch6qlQZbMd043Cxn5+EawgOWT
OSSMiul+ADtvL4FBr2kAv9VjLsZdMDsbf37Bou8k2clPrUoc7LR2oL9tVvIM0uqzXjujcJ7jZyO1
/tfrOQwGT6Zzfs7yM+R7ciBzSxQ3DE7fm5SYtCOrBy+XzuRudkP/FKUPOd+skKNcY6Wo14SBeHsP
rBxh5z1J38rwaCwv/kiWl+g7JziiMb7c+nXi/NOWxpcOjTcSL73CunYhZOoCmZpIu8cAprdPKnsB
VqpupS7dv01wE37veATZYG5dg/DxQJkL4rPG7V4UEgxu38m4qEhJAqboa24O+uYIZVJIz0bw5EHW
ECjroH2zPpIkI66vZsBID/UzzgQsMlc86Gcbdl3ULCMKlGPBk4/423mOvz/uJvQJTe62YePT1MUQ
oQLio2HlCFd6yoW8Bmu6u33OlJhD3ldTMcAw0evOPTqbbgWygjvJteR7IPy+1Nn1YEh6GfsrzgrP
Ipd+zP1Mgl6XaU8MICd8j6bKQxyHrqWBd6B7gVePH29+ysh/Vju6ajCPZ5x7UqBNm/A7dgPe+eoM
WkJgmoNVZRQSl8bN5KONYCoRsQdsUFk7SEwYcSyWhRbOkhXd6zKvnPVcZZVXHosOivDS4McTQ1r0
+oq5PLeQpnSUPbWqVaDRujdaPq0w5XYFVftxKe6tgdCG7742yNhpqO/WPrwnSH9uEospQstGXuyI
CwQ35eao+eNJiDgKENj5KabpEgvCk0C3W2zxzLVFm485IJmulDir7N6IVzIFunQAQb+xc30xVKf2
3FIz8VEXtnIr943p09t6Wh0cyr7Bv/9/Z5DDCjnzR//eBmsS+plKVjG9jjoNK5y4GHUZcTVg90SI
JC3bER0oZFs5chzIzoYWpm1g/EN8BEmwB4Cyls0FN2Mjwfnxsj4vBqPF66QBoDTylAdk+MC12Fdr
eA0RA1ocCHz0k1T+5+jJt2uLfZi3tvLAy0rwGuN27epaCoClNKb6wF50KCQUkzEo1Wyu0eW/cAXu
p0GVQ22e2lSFFtELGB7K+8GTmoaz5uRnVE1gqiK5Wry+xN+eytyGBzjUkKr0asJ7uB2eVk6qIVX2
+/x/kzHDhO2NrWU0HeGJFPjeIw7QoMwMldKBzyutLVyMne1HQb/VosI0by46CSs/H3ImzsJq6NC5
tLccdE7jR26Bi+LUSIcRX+kh4sQ8Fzh/hJeG0jnLAZFHuXh5U6v/+fkXHEfbaSoraFhwHc38pzSH
mviRJBLC0kExUisQKj8XeF5UtVz6Iij00U3y6CbO/UdW4/4Rd863gl48iHyewO+h6nWiM1t1Wt0o
vyMWP1ol0+5KTG9PxpNNR2nDo6t9wwEHDLrYF02YrJ5bg/qLcOZdB620/FV7Dkr35Ay3OeVaQTeX
qMQ0CeYIZXq6Sx0yqqj9am8pf9b0fYWezsuKEO1b4lYyH7dEC0FCxC9qqcOEAaL9jQcCnBoI4uRF
tunV9JmOBmcEsIzp57kpCaavWxC4+vKjLzN7nnQrtIbXY6JberehEc+sxbwphCBE7xkv51Ch2Tvz
KooAIG634rz3St9Gt8LxHlz3VIUQSjaDpfWDoSZ6ozWNWkU9hi8BRfnCDN/HwHkxrK0FQR8A0/rr
BPfk/bbhZvrx6Fpnd1XilC5IYnRNWHcL8eABWBqsGorwDsYEskRjRXU3eNa6l6bQWDMGGobOVl2H
KnobOwEXa7kmmU2swsh/2HffMhnQnsYeWD0xGTy9x9N5OB6rB98/ZTjL9GVDRej5AwzEcZ6O9otA
FtOSiJAxEABgcYAzqUAkJfw3aVLX1Wsm2wFDXxrLERY7NaqI7DqvkE6WTK/ISJm6lqExTclQUlLU
70BwtmNQ1k8FluVnA1Ua7DjHerI1IsKYFHHdR/IWp3zsC0J1eGvRLypsE2Kntfrw9ZvsMQduc9+T
W5LOXMzxp/QacBosxPVw7gXE3Ketv4v9Z5nwzj+1cER3/upoNeHtq2/5AAHz2mSL31s5u9/x79rg
l9RIiY5NaKwJm6rNzz8mENgtbTK3hFcPdNriV39aVQMOSg/rWquUqDNPF9+dbdOxjzkyZOaSfWli
SG2H2r26uSKMQGnQb8sOcCQOdlGuB1rde956rckyBb5748RUtPIofA0tNM8MLVOtlJd6RfbpTGOj
TwM5D/VxjabZmGYjEhCXiKrIPDcuU6dPSJy270G62Em5IqptcJMw5qwFjlHfus70YwynxZVkxEPJ
f5+PF3nkE9yvRUX/TocOk0t+qG+Oi6STRDpINeP39h5Wr7PsR669xpplejj8kAMEurSOLNwQyTOp
huRkREadObiFNrvcVqcW0HqkQuEcUyELXViNQmu5zVBRhDsPi/Fu+Ml8C+XvHj7kMkk3d6JaQLiu
lj1HRByHrBp+nmHJw0XJE1gdlZqaXbfTz/8i7htYNzzpHNxlEndRYGU77a7XYAImWZ/QPSbuAtOd
P2Tl44xThpOUpfSv+5Bja5ePyGf1r8ScHANINr4n8D+RgWYGBQwX4dqQrQ+RXEy40Wf6Pf9MIQU1
YGJElI6ZWueeNff530+atgtnGIMTzDelBA84QLN7jJT/wFw/vwwveJx6EyBbHVnVX/07o0bSwXPO
0ThAPhVIWw4IYn9IgE+/JyJZzj4FZwQU6EEJnHVo3qpcqjWNy6Vn2vESOUHs24AAq6/28zcGuSjg
4JdbJCMHsjjnIbiO3tjfSb5Y2pn4PpDnjz27QTuEasOijcDg9xShVmyIBLsTI8DwBF7iQ4yUvaYM
1QzrSeoBbYEKqw0FpEsuoUAjDNir3rsVtGoMnkW2n04R1ZqB4xbAf6F4+uMqXGkDDNFFB/gK6ZET
37O201Kfds0B4ZzkG13WtIcFvixi9mZuY1UMwl36x4iQPBghVIpAFOd+JHf6TirH8cww3PhUmbam
f2y8daMXtBhbKMSE4ZqUXXwW3TjnQKQMWdTuc/NpTP1rbwIbq3HC9T+N5rkp9MyLJHVD6eAPf+Q/
v4LS6e4ASbYZw40+EudA4bG8KqLjSxlT73rckFn2esZLWyHDj3S2Fr/mdrOKdpLUUplCTf3Y9SD9
CAblAak5TUj4NUaBsqOtlu4p2kH2trgq4txwVnfkYEVMhXnCvnfXGfwYYBnANNb6D7+uudSOjUDg
iykdOiLnLJTBztZ1j8m2vVz1I2WVJvmj6S1eKfpjiH//6apnDQGqgKu84/KVB22JVZOzjZzoLoBK
tECsj5bQHr0xxYMJ/dGKnojeH+dKxyf+3RyFk6QeZO5PPxVR5rsFoxCZFLHvy0kI4xmwKx1LNchT
d15QuCDuK3C5fTw9eh/9EGeOUdrT5Y0nzwBKJ56Rq00zkzwyx0b7ADuUQw/MyallarCojqUmS63W
dRa8a1kPHaIxV8QbF8sJQ7ybFTpBvHg4QXAyCgmNDZlPWsKXn9yv4MjRyEgF+kDyuvSui8hriZgF
QwidDRdUnMbhGev7pcvmfV334V0vimSJV0bfGbKCXi6V5UkEcKrKPux4AXy1v12NSzZpYAwz3Hp6
T0VZmVRaiNkXqKDDWfxcd+zXRnvgZuhAKf5YZLy9hz9aWYcLDEuT9R6g11syk8BC2gL1tEo41wSy
iovI7iCZsiZA1thSiAif3gFa58FKAgaIjs17HGz5JyQqmuvzEb3AJlniwjgxwuRzQ1P6eww4gZvW
t7QkEh2SnOhA8HQuByRg1rH6AQRTODS2KIzCQ4aQlrNrSaWckARocMB+JZXqpLHOr1KQMlJDQ3KF
dEhem+JZvfwdihUr6P4zVsAVSBZS7qSmMSLOlpzyQ2ampE5tB7GJCJQoFfDfsjs0gPlFw6HKDmfK
wr4fH8soPzECkakRdUVRv9huyxLq+72nXjKDuEp9SwuMWdufB1/e87PzNmAwpYspnMLo+64Gpkpy
kxogb0jd3WFVtsFTYW+YdZLX5SIFYtlFq/OYjXM4CedK8tymoyi5Mj3QvYc5nO4P2xeZz6aISNZD
ZuVuHenibWr6cfME1mycf5Swg4wz7yTpXbLc2NvWRfSDZpbZjJuqL6nS6OChMSThYsS1zxl2608j
/3VDUT9iZsAhFasyARDZAFfqD8CVS0wZw/xCeYBMUq2i8KdVp2T0PftJgUa6EdFNcR7TooxWCNAM
DnolSCjgRAIChDpK4fbjD0E5VfcC83s8WSpd6yar6XXhblEQSUtPVS2dFERlxbjCHYKybf75idQ7
CnOnO+RLh9WrUA6d3oLOcpajEudGaF4r3e344+K/0dHSLqmqlDN1jdy4eY8WA+3TufZz5ugp9ah3
ynjXFhLTnSsCPLEGkrAHtCqIEhmddK+8HZ5kzBTaEIIk4D1gPwlI14lPBaDqhATLsdypmLUVrlfO
1pmc5xhqoOkOgyAE+UWOz47zCvA08ZF4UWMYyCnFvArc3KZJUiWkD///V13BZp0U/E6LEO1mdb4B
4PdcvIGFxDupIiJjTGdc2rAIhENGvMUIonROjeW94dO4vRYZks37SLkghLG8hB9k3nQbOcJ48258
zaxmWA5jLg7tQbqx0sBBbDrecRtzeXSFcbEw6485LMICoHSaYp1aEMJQkLZlcTweFjVjf1yO9B/0
s9YqPJZdyflsZBDDwBU+DD6/dBjJTri0L4NdrWw1fvSPpS/kz8tFewyLOmjxRq6BJVb2LHJZC27j
RXl9qeSbuBfGSwN9aNAGXRfnhSkuODmLBV5Xgi/jKcXo/72UhbCd/UF/cFw9foZ5rCdU5CwK3VU8
o7qSt5SgfANPG87E7n/leLBnXhObsWLn9EzhKFECfAjilymy0a44sHtGQQas8EZeq29rDLcc6vXg
BQTe6+mXEWiDGpz0as7OFEzwW45np53QS+vUuum95wY2ardIVSdUMG+a2BQpMiiXdIbPn32tFpWm
My+HIBZgGMn3c5XR+rIZqjkqZZZe+/N/xOGu1BATVoevZ2ljI2L5xVC4PMzONS7Yrjca+WCCp/oe
qq4JHWN6LehhBqGf6QgjouefzQw8NaBW4x3lynbadFOcPV6ioy+BqGXo+ZM0Py5Bo/IN/dc3mzv3
HkU5LCn7dVaiCSZiY8CP00ejgfrJFwMtdmIjwR3ZPne7uWbxYK47yuffN00vQc1miUVPQYrapZNk
akW1wmeLXsLZTvqBWKiVK9zXQJpR8SGap61A1Sj8uriVMZaICteS4cULU9Yuu/aO70Pa1EwdUDEz
K0Y3MCrbVQc1aW9aN5H84e9o7SeADt02NO+NfHjy2peHg9d4e798FCf5snFXfX6oKOo1qCQXaTPt
pt2ayUfgCTh6FwijB4jPGMbOos8W1s9dKnyg2W8ZdRfr35r3xwvg9086Pot8BbYeuCB5n84jx4Vm
nq1FvHluBJNSeIJlLoDgibaQhp4nh/hZUG8c9MlMpni7RieDclH295cxYwnp+uTtx8LCyXJvUizQ
/0tBltCgecF6t9kadwY7P0vrHf9vWMej45wPlCUUaUPGnIYUqCHd3a88kSTdp1ixLyXVkSBrimlZ
Ivc6MjTZHUz1VuuAUhh4wbdFBI474i8BaiflpK42AdBN7TFB6pNHy9gcZbbqmh51FaIlkx66/t9d
xrlDUJgpGoV1IxTxwryuUxwYpW1iMRfL1bMaM3Vhj2tLCKl3ztoEG6SFmActHmVuPXVW6AoEgKfW
rTU40wf1z4AGZfPNw3kyl46Fg4HdeG0cm+qF5cjPtWi4Mo1rRQQ0+WafBCf2wOkJbGit+lE1KDnE
6lYSS/KJAb+3xrH7BPm4QWGnX82bBnqyfAqO1FAKB76IXicpPZdCfUl/ERSmKN/CnZEhp+FYLbRT
4sgghKSRZVExie0rMlZXIrPghiD7zR2WB103+LkqMZl9EY6UWUFUMzaghmcU+Ljbv96no8lrfE8G
gTt00yF0IKtc/ZdRnamDUQjMvjXgI7sFLn1QKYoGF4fXC40TfmMKA6nGozlKRpFJT01TFmYNVrTY
avefgrY40oliAHSg6igFSy6Jg/69ZJeiOSa3KuWIQ0hbNEbX6ASfR0eo766LYd1iIDsmLlJVltWX
T+sgOtmuIRVe6hEbTNDP2OMmCApEcu28NMOni05G0bOJoPS3TrXK3xR0LTD/O9riYdiZ5VCYO0if
Hf3RgrslUDsWlzWdqVoX3FRVWBW0qbfvGecZnjHWMc2NcLKkcVLjkNTJiF+q99aRDIIldMUxi3Gl
SFAnevTf1aOnUt0ousK/N/c6BoNtor7ioP6fszb3R8c+y5jPsL/S/97S/VIAAtf5QttG7DMHluit
iUEFg9RykpPUlKZWXZ5IrPAwJZJSsxp9WhFBnOk+fL2XK8Jretz7oZKFBtbhA3GwqoW9WDLIhnDT
ZFscRx7NCt7vpGLLYZJO4VXmw9LJKEwIqhW09BXwd0YJCe699lF/cNTMgh1mcq67TvtKLKneg8RV
8xk1kazSoqdLRya9370lCV3bCbw326w0/FLtYz871pTY3BjyW/7QHlKOatGKOqCfpI6MdDcRxw6y
U/hTFEkStplyx+Jjd4Rwsj0jvdU/fMJ9sCBnwZVIkTQe6PFbE2kfnDUjpRWJjKurpmZyNTLvFGn8
sABw9jHrN+8Nr1Y5evSJ16bG4ZVnlRVeBIKCK8Qx0e75iqBqIagg6PD35CFAr2zfgc7eEcZXPbT8
sywSufVWGgOpsyxP7phDW+4Oz3p5rzO3JWYIThByNXPUtTfKeiKMFqz+k7MmXx0CsI9/Z/8INERm
ODrE7Wvu4lU3lqn0BSaC0/EF0UFPy4q6dEO7oc/TGw4wBFj4ktXgjGV/yr27zEBor8PPWXe8WyNQ
87l/0pXope+vZnsawCI7lXMfaLuG6QNDzMY9l9eXb/wQ2US4rJqdsshGqotdl3I48qzBQf95Jksb
yG1yFtDexjjP3RS0W655PxDGArdgSK5oRrCQO4EJsELlIpI8om4QfVC6mq+g6R2fTAFB6yXQyJpZ
TkSyKeJVMKow2n8nP9TjQpBX68J7hzofW214yKr6+V2Sar/fklxLiuTqc4gKjJx2x7xa2L38B4Xh
HH15HwB+IleSU0HmNj3lRl4Nhh9yim9zUE9t2W14Dnsk+ir8CLnfYJ1qO9+lvalj4D7h10hS/qTv
hcCZZC6rMR6SI5Ily9zVjTvmJzbKVnE1hjZKr/IVDTGLaenwL/w/5JKFTK/Ka4nUEW/onj8fma51
M29cL7XajAB9MU8Zzsz9NnN1rhIiBdYVHck3ANFM5vMtSLKmqAUYeik8gQMQwmy+1P1AR6Gz/D34
TSaC7CBpaWKSy9pTzPNw3O+SEEG78jyOCnX+tIcX+iq1zRwkIMtFno1wLAObBZknyLV8tZXhdVIm
HhYUwOoYRm8Nw9KTScxAVzCxu57T9q181P5LotU+twjfI8V/Lh4uC3cw+sEn880fftbvYCBcE5Mq
9DVG8SNp0b2fWcAihaae/wBQJHbBM1W1tPM7KgBR93QwP/RcKnu9cnbyZP78SuQkjxealrCdNIMB
ee5oprIW9CKenKTE8LMWLljTyE9mMjXBaeEVwREGv7p5mfk3cu+b6KqaV2RxQvcyVpYVLRe9Krqw
+xqEuZ8rwDNT4GWXCEXgcU7Nv3jgqePKLItV6qGV1kmjTlbEwFnoTRg4UTs/J+2jAFJAKl5RZc6i
PRo2IOqGR9jlQRLKSuJfJNzSt6PDgoEi8WJZ5majBns2+JUGUywHX1+sufzFKyzGxDdRRc+VEd+W
IMRQs1FhybVFWxk5WvE8N63Yvmiz6umFKo8W2BrB2Ux1w81HO+w9b1ZOStzRaX847/1Y7TcVx+KI
1DwqjT6Jp7syJi6cqX6NN/E6VK2BPXsZ5rZ5c/zrp/aaMksG28OjHDS2QG1kJeu7gxCc6low6+1u
aVl+YOU/vmCyxIBAp8WZMsoVN8AYeKTPLw+VXSZYEJCROvefxvS4tx9S72D1wDAMBPXmgNEmrnrD
yNg/L0dNCviyEKC8S8vK2mA5BJm4+IiB8c+pgp6d7Ra1/MZ7NefteCaa+xiBcloM2wzJrX/awZ4W
/Uy5zwXteh//mV2BJD7R+SswpS6eY0BvIyV1uQidUSdBDOzzCXkccqVHoxrgCIBZDRXDNf9AEZyY
P26JyOCb069BB8ZXJ2WDm03hGEohggREUkkqimOuOyUDKyAWgRDPnribiJoK5hwqKRZJ/d3vFxBb
pzbYr+7IZD0UAmnU0d6isxjsohxI/bg38tE+ErDEBbKxfUWHN3NssW/9gGbiDeQ6zniQfgUwgQRA
L1uN1kCwteakE6+nPQaGrZPye9e7lLVPNMNwNQ/WIctDZdAD+BDSrZSDWgoNYJCqPee1OiAf3CG6
aEyqWC7y0RwO5dmrAloiOpP28O2xlU5mTWm58V5Bz7ptK3gLStV2iAV+b95DsJlfd4MOmWs7XSTm
AAA3L1yVJV3F/tXoStq56mTG+JrS6fSBLBxLrlknTYXtYYLQm7uNOCew3p0khK9BjdLRuDyMQMQF
ld2V7S0JUHB38iHmmCXnJQRa/OmKQCBzHy2dpBgF4bPOjiAjRxQnRj7eWHa5BDW8AZBd8hvsGwuW
NINxCcgiaGj5B4YrNhMyeTXmqMZHRP/rsWfyiwVIUNbfCb33l6ukYZh7wA5D0lqsM78yYKc2fKUK
A5JwloQzK/sZVvhx1macY3K3Y9zkkjXPVDQm7RzP0Ry0Tn+9vJ2boNtGUYhx8oCCbaUj5x+UqMt2
W5G6Vf7k5j+6b7siQbdHSrbteZXo2UxQbELij4zTAV0My0jCKihJyQ8Xt65kRDcpXpWkTZQSF7CY
ha3Dc8M6Cy3D+G6KoKpxItwmTgP8ipxx+tiC8C6ozQUOLVfAojAuhPB+Ud94FluNck7XdYnkPufW
FRtxz+2Ez6ypUV12ixU4V7BVYn7eJYbfXkzhGQoWfuhJgeeGeyMm9x2YSaLWIIjOIGTOUSMD+mr/
7etjeDssqxVFA+zVupfwA7O5u21oqVyaUW4cZMAmF+EuMUOhA5BCTnfakxwLCYUIXuu5V00VKDxt
+J7uiDkPA8sHSTh11E30r82jgvIDe0bnCFPHb3cKuFHa77avbnE3wGWDwJP2E0LPIlC45NcOYlry
Oah+mrKbgwJouePDAWzRkkiyoS9cxCCr/S5/05t03DSbbs3DugpcjL3It9IxoqLRfjTBarn7MobY
6qbEyuMvuaL4n9nnkrTbAUeJPIYoNv0+l9yYXF0ABis6z0IwZHz3AfAwr8cM+nAkUG8G8YJVmK9o
TTEGY9l0aSx6fTw8tsoUh2XZ85caLNwO+c1Y/JzM6NoH3SiuZaQqcK6fgQWqRtSMWyZLBwcztDQn
j9Diu0DvkkZqFAm1XEqSIavmnNEtVxCVP72Or0CPPliaf8usLOc4b22Ye0cuDOxKKJ7edjvHMo49
TUwyTKksK3gumfh11MAE8a1LIV5j1Kkhl0wRAD9qXOsp95ibRptKxAOaPT4/K5GQ8iWwpLTVD/nK
pwDvm70rZXBYLeukAEyzayM/yUlIbIieAZ+5VOOLqHOmsdIcmdxsfRZEtIWSkqLwE1fdcRClMiqv
fAmmoiuloRQl60L7g/4QHT0b7fjGeNN6XWlFmUd9QDjwZ4VexO4xEDKwp57BRxcTgobExoEnizZI
S0kZW+PcjcaB2GTS/wJhyEEOu9N0BpMes7ekXwBD2ABZvN5WsbXulb9Nco7lqr8fi7uotIVKj0ls
cQ/irSf9EQO08nuGXKkjxFfaGpICW5tmFwW+0m8LhX1nGQl3GMxQxoxiqfTYxBNRvQsMkkJHd/B3
V1y5qujUYPd3vDawShawg2UZE11oOt4hqE9LimZneZ9E9jDiONS83gYH/fLnBP/8YvFFCNTMQsL2
ROYZq0D8iPIEay1mrn+zVcHxxrRwjFjoJRpRyjEXMn0GrIe4ObkO4rcpTyaAE4SG0Xf582Kyu0/Q
yW8wERVc2WNaZDWMVfGKMPFLrJEG3YdnLXZmE6oJB6k+CgUYp2v8P1NxrYP7e6pJxxat7F8N1/Pt
Ck/UxIENMDfv+PQajFIIS12ZyiMPGu6qyIllhhLz8wHRS6hG1sbWkABH648nedP5ETOY/JDoGQet
ZSoNeJzW5ibVFZ4CqFwFunJvRswcfsLqJTPKcLUi+rZgKTt5p3WZemzNu3KSqV+IvP14Fwo/mXiQ
eJJ/Vd2hv+avSlRGDbTDY4DflAXKVfz6LB8hTgEIElEc4f47JBU7SYlzX31S213dC1fQzWGqUysZ
A7KGYSe4RxnVsoVqIaOzrHPjMZ+/X0Psz4LxK+dfDAf2W+THVfbULERh4dH0wH7RSW/BJwAbG+8Y
yzx9Kw6JnP0aTN4pYwUSMgrPPpa5fQwTSOWBwBT82HMHUE/w+6xSShwnheVi9WTmnY0RpaiAY3NE
FyAjW+QEOtWCpz0On1P8tHnz2//w3a1KBhFOy2xX514DM+ZU8N05ac5dSdv7sUJhkwziUFw484Pf
5bl2gcrsfe9N/UzCBNLy8StBaKQjklROxGiodAxdluokdrrN5C2jVxC0pa56O+yoPGwTSXWlGBdW
XizD0kfMsRrwj5jBxde2saSso8TI6O/cjCvbnLS8Mpt1BKTznxZ5HR92N2u6v28vo/OeyGkGxSqE
Ds5z+n2ow0+wvb+MX3fOfefkZFAXZKlYyjJ5HY/fE3ZnuJIddpAM+pUC/6PpIvfCctkliodA3ijQ
Yr7qIjEc99UGn+9e1OzrglA9qgl0s1Mx85QJiRt6fK4MErqC3Cg0uJlcuC40UAxkNkjYKg+5/AVD
zkietMxVsnIWscY1SiGRM5cBCVGY5gJg5peyofne7CB/t8gHYuHaVKr8XuY8UhqZIrUYhepBSYum
/SvPR3nrOtPIhGPfu5Sq/wj1nYrwkiq4Bpth1gbW40hkO5XEy2vYL6rXDf9aFtnnjiLH0Yi1edXX
JeouGhFYf4j9F88I5JXpRgF8vws1feAX0Y9AyECwL29H+swmxIxg2Pw+xjJoDdU/A0n8nimQuZKg
V+vVq2XMW2VAXqgw6qnZoEHUbPMCYcDPlqqTXLD3GJTgWpfUJgRuK9pSua4Q1BmnccG4koFqBqVJ
FgEvnJBgSUWS+XB21FeI7v+aLGoeXl4PedUoQnPvyFo26MgrdDlQpVt8TuNv7mu7yGjd1IhS+oWa
FUQxyCJ34FRy5xGFR0DmTbOqJ4hZ2XWxTy041CkKkms6g3P4dbUy6rPnHzx7O13x0FC67//DCuXO
4/Mp0p1sOIotuPT71ntDHSzQoSkoUl2DU5JRqqcKUBfv6mR40CGGP2fuyn8Kj2iQmuJrY5/EdBm+
vyzDRyVt4Cz+lEyY29CK4L3WSnDQJYHVZjOdUIt1mHudqu8hnx4ancyl/K2tK3zwPUnFmJsjqFoC
aa5+4tH3GvXwYWgCrDNQlQ4L4xXIklEIDAV2FS9jZGwYVi1fuUeqMn+eKUlLMKSbQKk+9oH9UYHX
UEH1z3Btne5aMNg9hleQYP1/jRrBP371paDJNzDuBwiY0DhJRNpTDNtHKv1SUrKKCPXIZ+Y6ji6X
taVlUIIcLvzZyzhLBKuSiZ3hv8PEh4k1Msyyz/uTKgvSauvrkMYfTFDPmBdWdtO6VWXBKVid5b0W
kyZAJbQkzP9xne0ms80aY2BOzZ15McJaj481fj6HT/gjQNm63LHfThTXDokeCpaYWxJZOb2kl2Uh
E2opC3z2fhJlITEY33sqdiFkDD10yPs8TO0W0m+r+Rh4m2nKx7ujalaz9ga9wNJ3A9MehK6PTSmK
cdEJt51+cH3WbiQ2f6tyWFiRXJUyYE1CVwtLBy4A3jHu2uKXSVkEJ2GQn1mxex0vXE9qy/pH2KoF
3n9MAcquypjZoXPyNWS3SLkYJIVaMR+/QQeLC3+eGcQTcTBjPaSgv/jUkDX6l96MDq9mjTedK12F
CTWXTpOyp8L8kJ1vG5BrENBj3iy1XBnU7KX39sOlszhYYy2oHI+br6mU03QdUjM0MyRSjcuseEoz
GvONgODY0QuGlC9x6LJDzEKf8bCBAPO2xdSvF972F90HBhey+sQWUB2lL2DWa6KkeWe7hYwvLxv1
S1+T0yG5bzLypyR9bgHJNQ0ysrpF52LqpT0P0SchE2I21nYYXhnDdkxxdaas3ANbwH6ACSamltrE
Paao0izWpqceic49ETn7+NzP2+QosHtRsfEUjcWecKtyaVMFpBIHFtjkHg2jHz8YVIOho2l2MSKj
yGq24Kr0+rvjsX7UtBBN1UPkv8JcUx8r3TcXwgOBs23phe1hJ1ch6q77ZqwoIeP8i7vcxrVRKTaX
8PK04CO7Kx+iFees7RfXzb590nKuYIRGPN8UMOAXWwHFBDR7swHHbZ5gs2q3c/oj2YDX2gbKdfuC
TbtD97lpchdb7nWoOlSu02fld5jpTj5AIghznnyy158trsQHUj9OhwC9a2R7I8xAiFSbiyimKG2F
zjwgjzLG4iSgjYhyjds20kYv3GjM9ATw91YgN+ImzUN1PZH/UO8YOoDXgpCSprAxoe3wsfyk9RbI
c336V2TUMxDrFG0imuSV8ENceAE9ExIPlZ5HfFnogjMEQIR0OXBrPlaYe6RUCBlvxAwZpfYk1crX
Tg8YaXTgkmTtoqMLns/pAKX3qYYOZKD0llOiBOW+AxoomX4rcj2O7C1uFeKixJ6Wisf+L+wwNUuy
5zHLSd0E5qSCdGtjjVZ0uArBiRJEsK8RwHdvuyNaMOx3JFZsco19TT4aGde4xWxMBnIjO6mQJNoh
5BZFyk6XdYN+YiWCh9L7jVrdMpejMQ8GsI54q725Jyzv4rF2OpHs6cIYTd7gECnBroA7tgmyfeDh
D5vE1S2SJuBb28+SthzucMH2onjpJb+KMapA6nz7S7q8d+bbL1T/Pu1HZ9Ndc6q/yfLvPUdj1fBW
mCmVA/KgeU4hVj5MCilrGvmpe9Wn4S0UDk1dRZ/2VcaavYy8kpoB/AlmXy7o/Ls6qo6AZeTY2BMj
oc58wzBlw+qXtNFkYPZSdeJwvQBiOQyRMDmGVRYASNxqGfBScrOPcnSzyUmiPRFbkko5kcZHmuFT
38mFL+5WKsw+4a+NB6XZRDBDzNhqT8uglAoYl7v0CgFinUhoL/Se6+a7ZreCmtHa/yiukM2gZIl9
2pvWqkq6fVAatUFkebg6wbDssq0XfQaXL3jHJXt+HMRpQEJ4C7uyUtyjljqVooiBw5ba5Wprz90C
7i0VLj9i33kkO/bTTMde3osjNv2GzUBo/5jTzXw9xSnq5AtKu8KTS2s4Csm5bZiXXuk5dcCMvdeJ
Ve3Go5S6SrPyt7E0oJ053A6B30UMbVgI2+XXCCS0wybY6aTa8cERNl7UbqA7Jpzsv5jPRSiJTBOa
fEnZVIw5xVwL83jQ59pI9Wi4ImdPmQb9nIu3aa4H6Vrbhq5pTXITtH/zz46Fg7RIOnyefHwvCSC4
n1ska5iYY8Bcf6vh+5q9Ec20Id6cnUEU9P7DZIPw4IYcf7HkH9xO1JmLb83HegnZyPDzl6hKTPZG
9DtG4UN9oFHgSbP9FdF3rtQu9d+ehtXUsVr/D1ygJBhTJFno13ViFMjjeStpbFm+gvsa1LsEYMx8
apRsAFNPrQsnSnYvEo9eV076IbuRjoNEpyLbV8RWTPR1KPYFmrv/QZ/yYcCy7O0YGdYgptiL95oC
RwIZBTD5HrehiQGvEBTSjmSfhgT+ZqR1g/JMi4l1pvB8wdJyxaDUrDFsfpodfK+CN8cvxihaGVWm
nEKX54B6stxm+EbLywAWn8g3S8lbhXLSETZeOlYZmYAL0saTSzOrzNlhfvMEu149q6zb5/zg9UJK
86jpEqVGEHOP8O0A13oQzGluNCCo2GAFqMCV07DdiI5IbvZByzmgfEvOl78R5X+IDPcxwy5DX2dw
MZgutjxpTQbSdI/+wGauIgRVRohgndYZQst9xST/rfl+Zr1dsadmBOXPMqVQfhgL25xUbrlsy5kp
x+8x/kT4zpZ7qzIdnIYZpaLcVTi3ANGeZBwmr6RWnhvTtp3lN3YlFf0OQfvyFSHHPu2ukoZnRd/5
kWmnAQy9YK2pWELEy1D1GHpAsxuEb3f70PJK4ntPHNslHinY0PlwkOrTnKVjuUzVv+Wd7g9KSPoz
EdfW9psinM/xMJiB3Gon6OrLMsA9UtInm9kBiHEJ2BI87pJM5l6Z4L7Qzy1x73S6hHrvBDgD+ivH
GYe5x6pPFRbpGfZZUECIbdTpoxVYe3tJe6phY8JJN2/bk9cmvAs1eXXSGF0/J3U8g8qospaB+RsH
ivRbL+0T3/kIxNska1bfnurttvk8alz5uKVD92PpPJ2PYNKyN+kkNqhFiWlTvSSrhkM0FcU3QsDR
9FsL25XvO3mDaLOdLhe0SXcC256PkdWRtaXK6sg3WPhvqRGinQWWQl79woD4aoBVQmFPSr5LbPRN
l+So5K1aEoJsgduiMs8JRGAs8F1QvbuYP92QBWtr8xW6PQp4HJnAU+MARzo6k2OkG+IFAVLFxXV9
2O8DhpMvCiYFPEnMHvXUXq2j/fM9dD8L/2gAKK9TuKpQvaD3qzJcA/jP28yuO+dwlPTWN7+bwY5r
0HLjs/ZaN0xbL5MJgRdSPLK5k2YnUuPy9bR4cwJHYWu1WXToqdWO6XntAY9GbaUmNrL/n4Ni34x/
M9ZMbm/vFsf4ePv5roki8Tpds9NMhYRBIjDnX3z1JZNtkZWkQzu8sTfHezjkHZg5aOzrmnueUi3B
XnAKk8g0nuGjUxk8lXSJhI4BtwDWk+kGYM4D5MOH0BE8tYMGtEs5nuZt9nGdqrVIZ2LCEYMEBaCF
thwfd2yO1lOJ9kHcteuxYsJlGz6BmDEvvMgoaJcrDMT2wiGeHj5Xjq0Z3DTi7/MOoZ1IYJeH2kTQ
UdeiM1L+M2lCnyW/KpDX4LKRsASYLHtFvwOLoxFFH7WY4ogaqTRRmVKEhFbgx8LwVRIWSP09bIJv
WjXRz6pKxOkUBZvuU1RQj+eM9M6klk+0NtTsQf9P71a+BdEBB8Sn/GTDgMK1cok1XMi2C1swjLIS
EAj71Y3+qOvIoqwxuiAlowKh2rbJB8mGoBU0Qy7K+84jA5Lngkzqlyc/jQKZ+hhkMeIoS6uqHEll
ERE0FwgfDcDiMbhUTPC3xEKOoDoiXFLXJcBM1pIQv8Dsp9RfJ49V1LxpBr6YLZ2tdN8vHqyjawTy
y0HGOxcH0KvHufySgh23n512y12digzNoOSGHa7Zz0tS9qvO4iIofzoI5HGpQ5eIn5pNCZWBlBRj
vedv6aGE2k4KaNQpeEdQXe+yoW5mVzdN2cnfV+J5DLdPk/6AhlNRHcDQRTMb05MyfOwRElIPWTf4
Gf2V/w4eD7mcv6Vj8pVSKhX/e/+MsMYIqr2K0Ym05pB7f6DQDTdKQ2kUfu29eKQXuEsHGU7E2KNR
AX/X+gF+G3hLMH68hHtYFB3D/x+HrwJ7er8dKtbeERRh7+gTu4cdHIv4HNZ0MiO4RRti+A3MpYia
hJNd4KfgvIigbM9sGc6No0JxRgxKhFXfaTcvO1szlYV6CIXAVGJEqjpvZZiaIetWzULFMqDTYiiF
cRAPwkzsQWQpQXfhJJInCZ66W/qqPri3VzR8N9hDp/KD2+hY+jLGKMflSZGAIfn7C1i0c349NFCQ
szca6E7cWseIkYTl+Rv52fMFH4ok58ZMe7WbTYFGe/lP99GXmohWucjoirUvaF9lTmUC5vO3ftl6
MHYOlIWMopm91DUyCDU57c2js722w1lP97ZAgc4EGJvTQjBmJ7ahoSQ2FnUf/rl1FzRbWnrZ1wW/
Hwl8KftEqiHGOBn9PYyBJgPjI48Xsa6eypURWp8vU85uOUhulpXqMtwgE2989Bf+mRy2ZELWgX3e
nKKCtSD4GG5kP/9WpLHuj7ODqOqa5e80WOxh1KvRpFxUYpwuLbL5d+SQGTaDJTz5YLOxhZoIWKQH
Mwyi/Tn1Ed+dyLFzSkJUHd2hfxHTd6ltkDMZ2Vp8gcNrMq5galaN+borLuwn7ej8fbaMTO/ax4gn
SNAGjRkb5+8ryAnSUnM/a3jgUBZOtNGwlXBBTIcXxZCHHFmIUNnisUo82fOp5+IkOgNgSrVktFQm
c7cRyJWUwvTGBq958X1DYno0tehiYnD754TBwy3bP3PnJR1k92fh0Lgje2fiEFC0uVFq3Rcin484
xksCA7moLCEERpJkG0DrlyRsvDUOB7s20xkWo7cO1YkOI7FnsbIIG00VtvQ2HMoO8Y1uD0DrY+Pt
B6ILH40iYWR+DAGcp/HTuBA5OVh2fOQP2I5DNeMghc0TADFAqvqCdCMyC2/9vTH78w2Ir3vQiffg
b44kz17BGsA2Y1RSN0PQkM6r4Hwi5e+YeUutEbxNM4FAsrJtwafUd0MaxbgFXAYEVCwNaNl7SuK9
r7+kKjLGTmwNCPQoyzOa65+lEO7Fq9aeObvnmV29STCzcASQ1XW4AkWUpqB4r5fkDsEH+1z8SOt2
Gd1mK44kscbmZEkJbOS1FRXqYXcUxEJc4aPE8+zNy6OtjD7vLqTQDC3k0Ti5bO6bumLZk1MF4e5S
n6TBSGL8/pbxIUK1TA2Usfo7woNUppUVIX6kQ669DAhCMaCDyJH++3Y1fWBIJuGSjerKu5bzd1wX
dqwx8K8eKhgf9j0+vF5sJRFieR8YldBJczlCIb6Iw6v0M3MntNhzqOOgTIU4SyFbhJWlyUZSyRZS
1xfOCjgynJvyFP4e/y2MaNbeoL6D5Dpfzwj4HacB6oNgqzVKD3MJjQp1lJ0hYTe3J65hLpxuIr7n
H1fAWgNxq7xwyzvlj1FN7cA7KhmMIdXblewu0lTgSZJHyT8FLUEjkjgMLDIfhhtYUj4cEYELMygo
kYZ2oD78M7n8sqdO3MNcA7HCYuog9kRQ7Asn/Rv/4H6rZQ7vLaOB7cOnkiHrRvSrwVZMsnavDnNP
yo6DmUTz5jTdJ5RbyTx3mwDx3LlmMKU5mXCHeYabONtYbcodBNMuQPUOlSaFKUxifIpR10opLoVi
z7PaqmfrQTZWn+RrTOJGHl8DqJdQXK1yQDPXR06JXm6HSGMTeUWfw+QSgmpaHGwzAH74myGH3rcv
n2LMDkVS4hMb2vcKkYuzm0XO4cFcM1ZKf5J91oAUatl+aeZeX09kRUkCjnlHg2fGDkQzheqt8XNq
WllOllhyJRqIYFPOQgufaypVD3oZo42o1DPG45SinFnqO8xidOVxoLDt1CuDJF9Crll2rqWTbG2o
YTEugjxXulTHa3YCo0YTktbw/NzNmwicKCX4F6fg9u5bKo04AmbXvz6tI8fkDLCizXepqtZ1f45h
hNHXbpFGEjD6ncJlAGVVcrA6ERezdQjf+hPZNmfffmvyqGHaq7oy4vjDfR2VraXT8lOoCYb4Qa/c
0Osbm7rp8a2l6Gtzw8Z8l0vnmQgaCYRbjIBaglK8iHSnGjnjTOPC4xhWIMzyr4/XCJJ8EzG1tW6N
fUKkQffuOYpnfM8w0fzRdjmCJZQCeI3MA3Nt6633yrL6PC3AQYJKj/zCFhaWpGH4brHrZlIHkska
+ARLlMBKfoJNyVnBndqBL9uV5QIiYrcNq4NUiexqWccddFOZdayyrbYZEhk1KD0SxQn6EB6dSVH+
Ha674/f6sGeGW223GXi70xO2ZTmZ4KlP4zLeHUSL9mODkYxxBBpz1wiwOPCsi3IymB4Dh+At/uQr
B5dKSxrriBhKYnfmZm3/Yq9X3gLjalGKvQWwTt/ov1VMb/WxG0RJuZgurjkk6h28Q2+WDJQpYZv2
AXxVUZ0/YRHwYlOp2OXMEpFi+8piJsFHk0CvZ5cIkT2SoBWUJ3QzhI5Tncv1pphrIJQaLQjqlq4d
ldM4mLQxgZtv3pw1dD1Nk7wGHgXKXh3Wr+mcNsT2LzSj2IXSXv3H8DL5dJaIyBDwvi+8/NP4n3/8
2t9Nv8jfypbCMoVl6pI8VwNvyZHXYGFF7WEJGX0QC7jK1Qr4bhNodWeWELqUrlwVfoCntY6E+3qX
0vIkFBJQQ+D/gMQNyjw43Tb4pIH8SKATt4wkVN+YHIBl4ZJni6lm/bS0JYvq5yd6M7YKquId3boI
PWZpQwlv3uKh0i7Sr4szTnPytH0zU38njSlwA3ANFV92HlOHfNykmToxlH6KMjVH/RTE69+sPZsr
2kMMl8PFlBaYGvs4zN3/umywHBvy37zQvmbCx7ZFg/2+Pfv+qH909VSoTuANT7Ei9OEZyLqYMhvr
wJ5jiosiJ9fXOgaxCo4VKpir4RcgF6D8+ZaflmJ8lEkMTOHhRukeAEQEzljLSn6OckBPlrCvJr9Y
+jb4osbVQqr6BXDRUGP9PcvMxCPu6tIxOaiyr6+bc/asE3kNkNWdp0dlPVJmKjpoofwDJ7HOysfw
O6/XCCMjTq2/bxU4qtNnNBBzgXad/uBITBoJljrmxPs4+KJMycWB8Ac+L6ReSr19HOER2smT2Uru
Nia02baYGpI4KFH4yKuHhSEFp+itKujE90B/L9iAiuMpHdbACAtAu4iaBUPoPu9tsjW7S+hM3Tle
znNpyNzFK2S6VsTqWOXBFeB4u/sHhsy/rLQYfIEqDG24r67ldZolqH5mRGpe49W2+am9j6xkWLBP
qDWaKQcOU+CB2JAPGpFcZx/j1yskbLJ1TUZ1AUG3xf/q+AWGm0xm3sv9VRV0K08nDVZqyjQ665eF
nJgzzVWX9PHBxfCGlfa2va8Y1yjXvAmFpTCD00KMg7q61dIMag6Rc8xQjQ1FFAw0ziPa5CkjkwB7
gcXSw4uGAOEEYRqKow+FCvBPh7h/6wB4ZBjtqMQ69o038MzqmdJUpr1SpPQ28sMS7FZAfAqBITOW
0+IAbsnmcoFa/gsJIp+SZaz7pVdap9nDAdO7xlIO9PSHabAV77dg7S0MNiBvFCoppTpw6zWZlUoP
22wP+h5bP3Xpj8+sU5e7J9sp8aJQ/7/YCFbAm9Eau9B2CWTqJn/ApBqME1S0TEcNmhwmwxoaey3a
Nsjoa6BKgSCcLUa7dCr8wSlahPXAfeiA7FUJ4Pp71aYTXLbfx21u5ZFKQ49JSqSSYucq8G/aMdwT
Bk6+ctAGPtnfwlfU92ftPHQTwOccMzZm27oqeF7suFi0g8eau1rLvY1AK235Sciks7Q8wEQepOre
yUw94d8tBHrc/MNVIYybgci+tevLNs6YXb9Jb/gEID74Fc9lqPw/iaeEyp5C99GN1V1t33ZvXZRR
jzFALpFxGig1P4VLWtCGu3eqWX6A7V/2AressFf6nUsks+UHNGDnPtLze9U+wXbT2nzjKVAmRPkd
ldeDFBXuRMERp6D+hqY+UmFMSm6Uk/8b8qVLhyUFauuE3MmHaMIjEkyG0h0HWV4eaaxRnsVTUDQS
uHZ4JPdes51M7j/BmkQ6y3zrjORim+3aaUxGyLbXmWd/INrZiRpSahbpZL1uFz3b499K6R6hTLSM
NBPVm5Jpt+5SJD47wQUTCaFsQZAZBDUp+65iEvQHggpfuPn9jUL8kbSaua23jYUlcTRBQkcYZN+G
4m+DFht033EoiGwCo1R/Vfe531T1+JiMr/YY6d1ZfWy7PMemrgM+cdnP33OpATtGWF03n0m2KkvL
9DF+TEGc9mh42tST6uCtIQfR1d6NykTXucPlY+gNKV7IznuzUSe2naU8zFPzIPF1ATccLkHoL4Uy
HAyayZppyTAE6sZcjNy5OrexbEsJ2Z+UyYlwjNImUKFEysIh5rC0ZJZdYN3SY4CSxv7LX+Wygyfm
ruc0538ayusHZSVpjzK0lspBMend/xjrymKGHxJbnxPZXV2K07Muk85DLA6BgtaAKkKneAkooLUE
4xcLC0ZBc7Fl20H71WIoMaunPTArDvPMvkSIT6Oo7BRkp7HwAOahRw9Odgd+OJzALkngJnW02Gh+
9X94bmZICHXABClJv7/K1+gFziEaO8Vlg7Cl3Rx8UbfUjsB/14g3dZQkaeHT6nKxXpNuC4sHJLY0
ETXX98hTDZhaQ/oMIPrVC+u4hE8xLX17sKgvPVZAWGHmT15SDZC3STYxoTjFdFwnB6cSYOdbOBSf
Oh701D5cvJppbvTcsI4tAEiUtzTdfZdT3LzXWX8OkIKVgspnj08Q6wLn8DgsCWrOh2ops+MocPTK
h+mPRA2kDrcBJOUbgB/SL0sy+BeHvRVad2pKj6x7967F6TBTVt+rEsiskDhMH8QBMfuXK0tkNSxp
VtIl2lW2MMMJjaG2iX/OD4nmQcPPqiIj4jFwolozp2IDWXhAfX2FB3ZONCN8MxOR/he9fXUt0tk1
J6JqHjzUeWRbNiLB45XeUVCNjq5kP8Im/Ud9jy/MR4nbP7yaYFnNX1fX7L+uqXnJyIZ0wfG7bd2k
3vDMmnJEdQF8/DmPL1R9XRx3zQGAx0bUeGDkUovAMQzbGIgrw0qfGiyqG1B/JmQoZzH5QE2QS8h9
1e/sOcbxoN+aeiEu6toLZ5sFrWsmDS858tcMdDN4b1pouQqh4xt4R0PwWwpqkirG+ceuKihEW8ez
2Fh9by4FF230lDFLszV7Hi2OkVBzJyBDPN8TZ//2JQStDKsnyC8ber0cCHbvRvsSjj9WrlLWNwUN
QNa2nozyH+ziSEx06h3VrEgGo6I0A1npqqL7Qb/ft86482oVvsfsKkiAmnr2tZSZiLeTQTyGZCCw
Y3y6B2bzDm9fON4HPowIMyObeA24ZX//Ui22zPfg7LwCfbnYywO6nRMZmh/4ij7h+ceYqwnyDV4b
Z7idCBxctOlnnF0Nmnn01Iiykk9V7JSk9uSBEQC3eMEZN0jO7DYFDATdb0xCywE9+Yzve8NQ8HhG
l4a9BMREpbcPgXTib7TzH1HnedT+TN2zcUSY9nxqCNEwrQaQWhm/+LBfs32xlWCHwtPlWyshRHXE
5FZcXM2JQyHDrRJ81QcGNdwwC4cm2VY7BAftGvhzpt2xpCAGvkbPAuVD0U+fUlc9schtPsH/oK82
+enuc54ESYwkc3kN6G4AqCsZuDLfYVtKV0uymmAIh6Tg//ppXBYi8y1OdaWkr0Sp12Q0QAoMlEf/
lN+nvUEXONPb3lkG0frBDIEzDcJa7hTZkKkzV5Nta0yKMITeok/nACDyWZCbUC13q2un6/HRD1SQ
P8y0mO3WSjQCBtoIg+yWXKEJIwj4mk5hkl/PDfVlaYTCvOR84noONleWyurVukNTKe4aY4iCg0tt
TvoydVYZqBOey37w6uJe99ZAwpfuFV/L3U3ZlSZdHizbhRhhSmGtc/l80W0QjXle/AQWf1NLOk4U
1kbUaCXJU87iEIGKtBVcdDYcEJJ86OX9nM0Inm/TGry7dR4AfLBskkS8xN1793nHERENk/2/qj3D
AyO0fI1lTi0hrtmbOFpGKrBPw2aF+Vjow5ejbo6GOh10FRt7XBjzMCztk9iO6iNjwjZiYRfWkFF2
m1dv9qmR5RyjMzkzXSkSUowb48ozHvBjPGhOn5gu+nrYKnHaN1rNM4qBsJKyTFsyiUKwFn+ezLdy
QHLJVxrHtblI2hKEIRSD93U5uAPnmJwkYDQNsP40bzE/6VPrDhYuqFxQB64q+SNYg4I4CA3xo2HH
x5J3xo5k9aZPeOZBOj+iVyTrQWYw5GhiG4g8OdgIQ9RufLB8HwkP4CNpr0aPgx9pDe7L277PR817
3D+zdh8CAzN/lPduPCo/VjCu6oL7SFhm0yvYnpxIoO7IlJTLs6YN1m3kag5VkMFoXjVEOVN/YZbw
RNaPfFcjyX1iALkVKmaq/pKddh7bJp3970E48W4dBH3PhTNG66lXO2XZQ5ITnCDaHk2KvM5pcwh6
HNdRP5mRs1E+csoM5W1IsiLeNKh+uivwdPEcMmtvx0Va64esK77d4a8SLo9t4XUAj4VurVpXmd77
JskzbrpdgIt+NEfLpRNB5KrnJQ/tFq7BrvoZvs+Yj/C5TJfuywZnfcoLFpJFFefjQIpCQCBnUmau
dKovdFtQHvxd+hgqAVt5tZwofdV2FW6aQ58gliHcUkUBZFZCLvp0ymkw7W648bf/UmSZh1tPWrmU
iNqqdf6yM/HNLWi4mWDCPzGCcCcLULa19tTveac8VKnIZF10I5Cv6JusnW2patizP9ASS/Xi8u+0
n2kipTPive6iNsL5J8c+a8Tfp7hdTYf9o+rYhAuTBLFE3vDbBL4c+7eM4dfNdpP4GgI9Ptg2uk1r
u3MrxVxfaNHmt0ldINMQq/o0WQ8eZ/vLKI9jropFsCs3bGfluqN1iAf0qYCtfY+TnedBy3SmFTSw
SxhCubQOevyQmUllTZ0UII9yTmVA4cuwqZcRxoha8OMzfK4Hc3UOmWtIH7YBCs8NLZi4s+cR4jIv
bfIKnlUwQkP8UvctuYMuqXW2ZxxBNR5Do37fGSqX02MnEWsv6pSyz4EYEPtvj1FReZpmsMHj3hin
eg6SwhnqTfZw/4uZ3JWyzHsE40GIE0N879Bgr4U+QXMOJeN06DTmEwJvdyeEHwLeAfHK48iEquE+
xA5bVMCQXqdxek1Td/TyFL1kLpGHGpAO6BzOq5nxwkMC5tbDA0shzFbv6HriFRT+W/Ie9CjTNtpv
rY66mP+bS1kHx4mjiS0ervJscvWVcNm1tb8hiavOuNvEXODwPkx2WanvwKiGs/M5UszyzFxMiv1k
9BLi8WXBvGlqeX4RDh46fzS/irP/t2D73pRZpr6wugA1cALQqJav0+DJwyfZ721S/tkkDnt+Z/Cn
gYQlsbgkwmxEcmf7MH/NGR8AjOHan4oqKPbl36qV2ILFbeolHJWvnpYJY1VVhvMKh34lUna9LZwI
7nPBRtlPZMKhVTf2GdSaVPUIOwTtmIwsA3+FNeS9kYnJsT9BGNjkH6q+hCzqh7XvzaoV8YXSqM0k
tjQiTV+5vvJAnpLYIQ09VAfIkjnxxf7YNgXTCEZGVpUVuwQ5p88nEk9b0bStDmFIGpmQPvaxutso
kiF7I36Ky29T8TY0EqYltyY51pDay1TtaeZK4KfDnq5VzHvLdUq9dGyd/hz939Ra/akGH29V3l+F
cGub09JwsHrfuFmnS0JF2BA1KzZmMnAaaZF5+gd1OUswOr3XrUSsLEknPVbMnenQBqihtgvH/2lV
bmkNZqLQ9rcHQXnBcyrmLBeZctXIOeQfzkYq/mFA8Gr6zngwR94LTkp5VodNb+ZXFpNoJ7WRruyr
BAldw6GYaPQ3UujqNaiIa7TiVIrZRceTtcUXj8FcBhnQiCg3/g+9iLgACR0Gbn0XWLHaB3V+xMPX
tUlc6HQeNo5gkGq1RLNST9ZwuiobxanQKBNninrdB3E3Wrbi4iQrmaHT4E2RCJmBurNqHIarNY3d
txLljt0N9IWOXpD6ngVkuoUoThT0EyBmL4QyVxJ166Db1OZHx4+zni/SJq53l4TvSwZvZ7ZJPCPy
uhsWuxClrrQbQFAEwu9Sfb/fr62JX8SPPEGWIeI6aguFzxdtyT7ijtk5VMtcYqthPJWauGdL7bac
dIdwQJGih8UTq8hbpY/T6xGA/sw2tzbubSFSzypZ/O9Ywer+W7K/BPhGlTSaYgYg4n3+DmkAm1JI
6f6AXBBMPx3agqxjRl7qlRnyONsimowrDRoNcAdgH8KUzDV4gdDoOpk9I6m2XHTRMLLHpmUKkhxh
BS6QP1pv8xeVGUr/Ux7h6lsBE07Q2mi0AgmHA1eUs89AoNEYizzTr+bZD6gmtaTILWiBPtSdUdyH
vZV+CLIop1afFHEQ3+vpVBvNKeEF+x3jZdgfIdCpn+m11LnrC7Y66Q4jirVn3dzgFS4Zautqmv1X
W8xhqciSTELH+/u/smihE9vty209+jJFQ3n5sCf70dNbOy9VVWGuuxYpOdHn8bZHEZTbKKZ3pSfm
ahYaWcNuxVNYv1TP+rQOSQEA/tbRS7dqGjeaaLOih4LPMchBH1a/fGKaemnJk71ur1swQaAHSUhv
+mC1TSsujpquodVD/WMDcbzc7jYQFCKjPZKbW8dL2DASc2NaCb3Ubcg3I2rrwNvcoc969GjlAfOj
0RwA3nB2h6w/nRmZW/wRmh29lkxQ0atxGBaP5z1TwrjqjyKaRxhRC0tOaX5UISlVAYDuKMplPiAa
8ajspnssWfNcCoLZ0/wSSj/EraElt4CgVkGpD38SRioxz6WOZmmLbGW1foEdik9pYd9C9/FwLGuv
e9CPWKjFO9YLN+Xbl9EtcKMkLryLxP4aimYspjNOSY0ga7cJxiLZyasFRfXhVOKh/LzBJIuxcMRk
ZmKzQyDrCD2O5dK6ka/SLW5oS/pjkXd7+IswhF2C403Cl4K3Z8pq0H8g9yJV+vUSYNby+BoLtXGK
ew/+wQEwcmv5KkmW48f1uUebLjsxCQlIO/lbwlxfWQlyNeAOMr9oA6DcxRNXbhjhq+pJq/4NtNts
rbO0UbOo7e3KUqeIV/2IwqRdxzoX3IpCP1wgpXP/aeYEaYICOVOD1AsvMVWLkP9ehmcZcJpqnMrP
1zMreGBknEq+UB9JSbeSrv84DatJCrABN8JXvhlcadq48bGDx4umwZvJipCXSFZc4GwH+BOAuOxb
4lFjDohoxDsWkZWe5pePDTivWHOWPXEsqxy0sOX6HJI+9L1ze1h98PcwbQZfVPJcYG6lzRDHSfQF
umHs2/EnS4ODZmO+DpOW6QdaqXFAHxH1/dMkwMxwcxfog0mFtxBNDlpaUPdIrBRP46yp9Ybr2bO6
oZdx6uKEUqTY99Pq/ywF3q4jjXlEKQWbHgeJL/RhjP60yTazxlm2EaEre80Zxb7EEwHKfLX93wnQ
0IYu2wWHd0nx9qGLBwWC/+LR7zLsHeYDPfy5z/PU32wO48Hphr+Ikojvk+JFIkUqAeBjZXJ3Unw3
Mw21SJ4UihVTYKUdvqIr8DelelyE/vpF1enBo0BJ2bOJIUZ4h2PvdYybsTbwrM+mWAtJRoFvG21H
f24MCkrHvkw3Cqm3CWFQUrNEK512Mv/UOUbNyXRY7hFWQAxI/Lff5RRou+KWRr46bIWaBkbsFGM2
mWAB9w8RFTVDq0ecZw5nqcHTBGSAC+UhEVbmIS7ZcmOTzPewkfwxdtEil9f5JJLSUYvHbHQGveae
uICP2N/jxSTxUDuZTqwAxS/7JRFhNP02vyycsgl5OfkqljOxBU1Vlh6SOPQ/AGFffsup9oVLIADi
8PpY/Z1xVv4CiiyqgF9xaLFMfG4YKFW8VMbDeW135ndir9/CwfjXhbDPGlCJADggkuRYa7KxVj5m
B720SrFPR+TqSC0U01SOsQcHxuWP2ShICjwEpGNQFx08BfGLZ3HBzvPSBOh2Spwnr9yX3TXiR0o0
VVDRZ5Gh3qpFVwESjqvq9KS6YMY2wfzy1o38mC6HUtp3BtaZRZCaH6amO0+Eg2z2X6cyaDfnSfX2
sShYC4xHWcI1gf5CfM2/HFXLaNsFrR1xv8BQs7ixUFLRBme4r+chv0jX9vQ1AnFCT+6Ftido872l
0lL+R8EN2I2CEFbYLdkY1+zc4+Z9bC7sJuuLEZB0SXf7J9hyd4A7Qn1hFqkxCfGTOETEqCNezFkb
1l85KIH1DJgVP3z+p76PmT82YMfQUDc1oNSaDFqORdMYehb5nwjXoSaiowBDEi79d93ir+omU/0F
feiaIMLBoFpG43X3h9smjG+5+IKms9ZT38ZTsAI8DDgfJul2xfmoFntjGt1yU0WHLG/uq6cqEp1c
FMOkaGtSnFEY98YU86Rjj/ZIuXTLHiLjg/ghE57gHro2I4vE6uiuCYw+IGpA4+FajeoTXOTxsGTA
tnWVzvwjWZO+Ptu0hpd27onGa3ilWYH5GztRJy/EFnYpt9tENmOHhbbPa8WzOEVDMJkA5/kgKMvy
DKcxvcDKjkv/gFpetahRZ5RKZTaHOYfBaSdEXDsvavCfDLfcMbzNRC41PoWPW41fG8SUiT1YnGEv
BiqehFNrWYE67jU+PcVkkrhhhX7GSVK8P3eEF1xt40pG9zP+irsvs9JtD0QRtGehLcBoH4qfmJlX
nv3qKouSXsDfFO5F6HYJVirMgkbDba0Gga3VKKwPdRu3HjNzAYix0/aY+CUzuqV5Z/L0KcF3OTM+
I7h7h+VqyeKnyId6T7QBdKzfnk5oxGMEqwiHWsdMEfGUlEbk2kKUakYr+SmnPj1Obj0rR57kEE2I
uYadjWtYJu9Vr8NZL1JKBihbJOAMtCzUVZmNcqO0L8vbK3WsRn7RZ64ANP+TDwwcEQR65uBZPXd0
kQmBR3gdF7nGqDu08FCJvZUsQYq6PxpFwtXWjdYa2Ijn+sQvrVXNpUpH/raB6r2sOkHEUq6DDHxx
rW1gzn4jgwmcljsWPE/cm/oD/RoGMzkPx2oQTz3N1Yih+mCTMvvJQ+ow35xiNC17Di9+Hl/wSLws
5CJlwuIz2UKbHlOOyjMgvolzMQeDtf+1AnXGxONeyaWRftErsu+VevWRZKRmaAuK5ng6LlvT+0gD
LWEPgFeQeauHn7sj++u2PYj4XYA9M9ixUN9wBn5mtnUvR3rszWC2xgou/yGSISQ2mqJuky78yyPM
7DML2sWUi5ddpSCiRfKKjQYem+iOw3gluhImTQgf66/2sybcN1+pO6HodaH3zUEGla3fb1ZBsOLn
bKSAc8l6XL7nMWZxmQHGDlfmuUWwmaw4+O8Gqct2p19sePg2ylYBn5irqIklpNQxPVwDSnx1L6nY
lFqT7mPDzFpOFyz/zVpFjFqIKk62Aye7CuOOweRe6nvF4vfY9lwsCGACw3afs6pHYH3uMDCb887n
rjolc1zBahLDjyeHmRz8WYdS2jpK1v1VNZKQBUeAdOn36WpvsZWqMbZJ7qQSfq5HFQ/QQSCUxX4A
rU0yCDaDbNGfUTd7Jtf3OybT6jLT2nqrDC3iEQK6Q++4TGRU98783HDNIJSR+BBVl73AzlD9JeaO
IP0H+HfBZKtcP6vacADbszxB5w5fcd6h2kx1nPuqCouE+Gtj+F3gE7l71oYiprgwmE/1mOP3rNnb
uowwVvmRgimQNJsFr/vbAkPDgDkEyqo7u/3BWeYQvoKM5o7xZOLbOacX/j0dkSjKFR+MQNYnQ4Gq
ZyxZnVMe9SKRsM9dhK3TBRJYxrd+tkkiREPpb/wjoLD84LDrXbz9qKUTk4zGF6S22ApZt383HRHy
2OA4dZjshNvYU2v4Pi5/RN/0Kt9/WOtuY/O89/PKSJzIVc3pBb6Gb2pGRYVAxMNpJnR/mXmlPY3u
Eoh8NviSdPJzJJvTHaS03wqpsuwjd0nVGIpt6Bj6dzraOr5rqAE67J3PxjCm95ihk3xHS+xvMSPh
JEcDosoaGP0hq7xfufonV1dYzx9LZS7PjbDk7ecFx5ugEOtWbJAt4JBTtcVMvOoxPBrGhS4wa/cx
SIAn4yveJ0bX3yqIAOQbgqPkdMCYa7m7eLrnuljXgpn5KqdKy+N83nckgI87J5tCyFhlYjg7MqeV
dfYOrll9UT3Q+ijbDDTliA8UvWCIfMVr0JOICmMw7sWMpMFn9BHGYSaTKpQ69hO1z+39K9HAztdM
/KJDN1RLVN3SIOhlqZMQFKabZelQWgaFo2m/PtOP3e5Mznp11A82no34BGkbATMnf4h/VN+mYsoM
YKd0RYti6NauQF4xpS7zLtTFaZ8y3he9vQbLG+QiUnWipJZ4SwOpBa0pvDvXcASVV2yl/Hu3WIFg
s/LNWKTkIXL7YV+sc4UhNWSDGI3Mu+758CXPOy6UKtQ9xQg0eS/1pqPDK6BRn+Lb7/hCsEtbIYnN
kIq+yAgJODrhiZ0iaQX7Cmw1JEwoejuqZSOJXBSPsKyhRVx1vMqAITxjQAtJ8+ol+JbEDyTcrt97
MQFxLaYwMDGXFg6xnEXS4ZjkD5hPPGNUBNYz+9dU/SKXCQF0/n7lN+IWx8oekujALi6ZthwzAPaC
hTc+LRhnc0BGaM9nyUnZ4S0x/48zVJWm/vvD4W8EP9+va4imV2x7vfAikMNx6ahXeVVDDB2aUhXg
uDCNju5n7MJzrlCikAxabZbeLB5r3LZ/zlNIH9rAbjCqvvqlFsxPTMJgS7bKH3yZLU/MqV96HoRO
TxWTTBlfFAk9RjOaYAq19xzyUgAp8y41JHE7x9AyZ/0hjv2xmFF8OUnb1As7hYf/Jp6CKznjUecq
TZoH+HkO17WULiLj9MGApU+Lp7ibsf6e3DbSe7x5ItsluZRiLnu5RomdzsQGyzoHQJoZrqApO2cr
ukY6vlK4tpfH4bDgf0vEDEBBeT6GVVfXF206DwrJeZ0TwFH9W9s51+Mw8EqScevCPz17LLKmcP2c
StlScvRN5dQRAYSG3I4kqIb5YPactSoCeuQHE/psMeGMrNsxe7S45BWgVECDbFdCtyY/Jf1I/NDn
bsWDgjVb0S0Ggn4u4o1IZbEafEqpM6rOlr5+auJVpMMhnS2gefWL+JWxP1Cl5ySPoSpGCFlh4+/+
g6DT/Pxlbz1gnPDO4NNEYZNwnPPN1QRfZd9Cel9Xf1iidGrUFv4uA40yb3y7pa7e3lNbW19r/Ttk
jzwfQohpGMEg6R5kAuFHvto46pL2sgs4gG0G2tKvuAgcSNF1jn8k9C1WjUc+nGQb9pWMonwTMcYz
c2vUsOb9/rr7/aWIM8Tkz9AfH7xbBkd71cziWklshZsVYaIJxSjBF1BsTphunOQ3pxMiK1x9WFYc
nf9rN/+9yK7CF2MAr2DOJNRECmMp7lWH74N4vPKJcX+KBUChK0E3S8cLLpqGETcEQCviClNFLwQN
BZ+2CgK+OvsuL2JRCiRUVORuaMk9Rmek8RplRdNquQgjdSuUYY8cb+FSsJOL9x6mhExJtZGXhtyI
8cnfuMLthpd+F3LmooI8N0OVyTqlApoOsyuk5hJKDTI2GR8P9NRJ5Z6m723+zIIdKoiqv+QJ6h1D
iV9VsMUMvcHTI/zJi+WvNmriWJraI6kjOZFyn9cV7T1uqvAPL4wtUoLLgZUbT0AOxffSBvBs7Eqa
CV0IizOZiCwuh6T0bTo7G8bpaoPX5OzM2FkTu4wWeAYm7apnMvbbzIK8HSux12+RHiTLcTOEBxqG
LOX0DUZcUBhYum3JOps6ClRZTrQEPez8sWKnEDVHMAXgod77ysXBJnNFku1wuIcIlEyu9VvLhwGd
4PWH3DzU1pH7OUgpAzg3L+Jp5CaGGEQshxce+3zzOBR9+mgV1WpBXlsLl8OQ3tk/e7i/11DmVVbZ
XDpDUOwBhAeZFLTnj32WSVUEkWMrH5seaSp4euS0n44dOLrs2YFnxHrki6Kchy0/Vj65kbSg1stZ
n5DW3BtzmV5t3HtTUM8IhxPpoF0+nd7OOCtxS90xs0HhnRrdRJNxBsOS4v0sA5HRKSm4voJ2St+u
KLwD6mEoGvbc6BqY+uRnkYCENtzXOB15F7BkRrOcR8jGqQy5rr5A3AwhwWRVOSh3OlHEk067g8Hv
Adg5WM3vfuNXiLWIr/YH2bcfjSEnRanu1n5LLdvKrCOCyuVDcDlkHgCaVDB67QdEhUflaTbXWM5R
/to4HVtX0BvMZQ4Vt1XmASB1DZCGqYAkxUJAYSIiOSbhhpzb1V1p5snKg3FqKPgbzrIkXxoQGAwx
0DJ6WxdC/E8zDzkyChAd1dSSBcqpb1io3XvnoPQGEKAlUkzkwceixqzNDTGGOcuCe2tRyCOUVbr1
xid2D2zDyuB0a1rkHTQuRLfjoJ0ez3OrnelO40c2TLWhSstMBmTLXlFW8KYT/GaCNwVFWkWm9DWH
Ffr1LmjV/NXaKdfuHwN8TchdFvlcUr+4WqVKRhtHhb61VxAossuew8usHPHVOzSjih9EryoonuZb
QyGdKvVz90xb6KNbxP2HX+TLYq6fJn0/dtuhDeRdSLEfOgdV71RfIi97G9kOQO927W9PZa6kolMB
0pumFw+uEy4+7a3fTIyZjVZrtXNW9yvCytQ+mZpzPsjuFmM+Zeox1JtMTPMaen7rq8EUkdKjwm7j
P8Z49CfAWsATT4tgnYzJvWJjdtx/XyidorvDCaoQeJKQnqyhvdnqo/HwCk2lDrpDgVgcPYQr6SBD
rZ5toy7aT5yto7khUUPc6NZcReAhugiWEDcrAbRs/9AxqfUblRWGh5bIgcd8mOkHVdPQutxuvNvD
VTzatqyLjcNOp31Jvp2LHndyH0YeXWVfVRjI7DEzpN46gZIpbNkClGg70DddUKTD1hMfEKEk3fHo
BaYR1AZC1x6OCB3ow4DBw6YYI607ICdZNKdjrU/sZOsqUnIkVodDCGYUxdHt9D54vRE6Otsx0XZo
jE2Qe6EMeJK2aCLuzyoTBbzI7OoEOUCNO9GM1lGyI5f/NWY+slsRuFP3Pt69hFYArYTXRlO/5Zrk
TwM+q0vnl/pJrtdp+HMksO6RC72Ov/p4mzkWpVgwsGbQdRho5qfPGVncRvMO8aEKm0DVaGS6bj09
OgEUjYYxXpIdK76m4dgm6oYSE4LcpaaemZKOtcm0v30QKSNK4ZXGILf1mt/81ZAMjQjMq5OAN99X
i6xPEV4nOYkxicbbhNGHrTPR7dmpJRq6t3tvmFmZPKa+uBqiODm7ILcsHBlJ54q9sQE6gvIlAG9w
dZ9izhs+PuDG5dOcWueN4tVlnm7paiEvPDeQP0kJFl3hiURjzPM1wZYpLHIxeF6GpKtRnRV6OJc+
OBAtgtUEffddQuFl6FBJM4hmFNAxyw8pOmXq2O36elJUcu5VLfrb+xIis+j+3+tUUapeOABZJkDs
uTzG0Y7jYdbsCSl7Esg1yQBG7veqfyjNfnVGhDmj8N3OHCMyEWSQQzlspiLr7XQRgzTaJao47FkB
Gp14KLT2qmUsD/iCNCQtVZx5DZLCVee8f1maIyFxU2LtFIY0RTbXIokxHIjQRvbmMsWByutOd6uq
ROerA5m3zMHwQgXEAiQjIttskSBlOIOlNeI+4EKFBx6H1RA0X50Xm5G5bc5xtVYIiOIhPw1BbdU4
cCHG0Q73o3UTYAcrzULUkGSuHcsuxhr5WIDfVIAsrxjPalPq0RMuG+dbaDBHYdnKtqSZxK/rCJD2
2RaI0Zn7tTEqDEHADPLXfyAMYHo4qZ4kjm7lMFfMHjh5YJCB1STAkDomRyEatKJUzVkYdu1DXeq8
DxKdMxmelRu2lWVVvUBfxWHnRszqcs564hNGVDmi01eIBkcmzxHH4faMPBNFHNHjpDcuKnR3sbbP
pi2ubLoA2vjKHGERGRVn0LaQlTps56PKCnuncb3CKo75Hw1fWJKcbahF778VgKrRY8S5aUpLBC18
vPeWGfOQfD5hTbYZJkqsyShsoSbRTXoocrGMIgGbazZG0UQPEO3ZABxxpExuqlW/x7DaZcfqezD4
ErTRcnlONS7CqE08ZiF/gCE2rYJ8ADYBetRL1R4XF0RkJLoEGHS52em+st07Y0YOeP0yrtdOoMb1
kxw78/vHKGVP15MVLWkB/2nMGZo0sdkfO2zXaf1woOnpeCh/AB6GCv2VPMmXCQprXtIjvsNp+RFe
yYV5iKH5OQzj3Wq3N+Wk9EdRy0Jsu2M8uMSRW2K2ssg8zi/amYthqBHqmIg7WwJQ4oBlYMHmc3ZF
GtU4AXzg7I1IWtrvJjNdnnqlZ6rX3kBdDAp7SFa0teC4smhnfnSJkWNMM8BN62s7SfsUPh/Gk043
aI/96VdZjlSkEAqM5ZTwRmt57Ig4d2FtFgj9AXy+jtqdy1Qn8BE2Kmy5bRtixexhwly9OcJPOMSW
/xdsGzJwj5noJDc8BEPmyEkq8os9HS2hUtlGul4BqQFppqzfy1z4pmJpkgEXBoYWHJvVlqGvvSLy
3tSHWKOr3WdIBg8yGy6zWK/8f71KP7Jqn7tqDtTwRKzgYBgMJOk0mbheLjStNxVokYnyMSZOA/a6
MZudzdnAu6An/HYkp2b1+WVR4rhPBJhfoqUMZsjsmFVYeFM3+80uvYA4BNyRgtRFl/dEHxd84Xxb
TuE32o29q8p+YylxpNjhcoNfH8gAhTlYzNvJBY/2drozr8ohT2aDZyDUbKEQkTuJo2fJhgTjcuIJ
2n83O66cyK9ke8sKnxutD1Jo/QkRSDXgqoF/BM9t/Yro5nDQBMhLSDrF4dgqPJJSMAeM5AN4Avp0
c4Ne+CBGevUk4LT42AM54HjfAevqbgIVK80U58kGuChrEs0weAYJX3R8kzdkfhWI4N3s3mObQLhW
rIHFfuo2WdvZx96xVmei3Y9cpnfOjdPHYj0byHI4RCag/VFfztMl/XDHxSdon3Vpug/im/W324HM
Am+jOBFSs5bgz6y0/bKpd2VwoU8T//Ij2JyM+Vr+gQvmIamvFPqHixQGYVPgqO8gjWuDP3KoEuoz
Iy+MVU20dLyvlz67RvAgiSuUwYoVh5ydFpUP1DD2PwiFrvmZsEi2YZwhOrsVU+ld9Z2akKcMRgUA
yX6bvfrAw/53YEnDZoPRc24idfwhrhwAJegUvEeQ9msM/txzJI70/OJFAM9rrl3JaISVeW2rFAfe
II9La7yHoPvBSy5EVqKmqB1/aXhwmkShwpIxzJ3PaqZlkAmGs1wPsRYA/OyC3fDhNt88Zu5e1+5E
SmKHOiy2i7bX+zxT3FkPlOuvA6SZPcxVQ9u1m52cYAeURpnqQUkoFWpAHhcCOz9XfOr7SwUtQq2h
ND/GYDiK7E6nukzmzaAHLfq8gE7PdFOV6QljJwTGVEzhKrZ4j6DW+8trdTaYw80U78iMyKLCSBa7
FL68FEUjK/XQaV65+MUQAC7mCXGk0gNGia8lWv/L9/UzCF2EfgW+JNOQf4PAsFzmOsN0ItMBjqnc
Hj8ambiYpVk1HbMnyXYiFFz3IuZmemAU8p0HaCsRVrLyZxmCi3XJPrVxFJ+hwd9kQ5JNPrA1z39B
5fYFrjnWQZ0fLDY5JTGk7OqJNUhYlBkSCLpMYzq9EOG4xoGpo2QR+swp1y7F092IpDc1FDJOUPcF
5govjmFFBupcfJcXl4EgMJsAB13d6rLcNMipQn5It11lw2TvMJ7vfhxJoHSgWAFy0wUyPFshoEO6
nC/iaW8lqp1edjslqKHq2Gjafugp0jIwEvLQdViFwowhko8HprASHDxb1guOLY+DRToGkILQjSzF
ocd4dfe4MgDlJu2r/V11jRp3/VlD82EfUlALkRZacw65po2EneqXhldAXYHeyTyCjvlqUdwJiefR
YIlgrO7klt4I648F4ec6tH2iIx7ZyVYEw11Wu9B3h4hYWcF/H6b29dok1j/5ASNt4u3idaKDhqD6
mbuhS1oGGD/+JIsPlvRjq95KADMu6hBu/8EjTOnqKyEC5NwJLvSP+x5eykX4LnjGTqFYyhdg8Gt8
kj/860QvZeh4UOfvXQfcLi6ljzQVwaJ3DkOEqR1uT3T8ZF9foLJJxJjjjdpetMiE+WZk2A9VlGAF
0bNrPZKp48DFXqdHsAokwMu4XI1brFxRwkLMJTMVZcZnK5wLv7JLDkg4DgLtpNz5XFt8PeZt52hG
SfIiQepHylz+mrwtZawXAGJ1SAO9XsCEBVoV6egNmFfB6jGxecXSzTo88CHFTNHhxCE0y7PzJF8V
QbuvIIkbRfuB/BZXFTiCNW+2y3oT2/xLbgl5gc5v07SpjGs9917DBKphYjOLPPDJeq2z408HalWc
4bRQRw7Sa5MnvrOOoizepq2sjrAOjDpvR2vBNAxreNUFmYm0hhsVFUtxrpA4MG/dCDZ3PhOHubbo
3oUO41NkLrQ04NHSDMA76owdG3FVnnFORP4+2vHeC1m3+BvmwI7p6/PJU2R6Bc50CrLyaAzhECSt
UYMWP0zk6ZIGA4USBrg3AmLdlPxdexXI7d2rd2IbxGr7wuOuAyFLh7GT4B8vEEiVMRGtyMWEe6t+
DV3pEwu2xW4ZYn3AoVZf7mujsJGB4GMUKgW7extZTBwWuosOGIjBou96lfOl1s4ASoehZHwA+Yxn
dB8xCNATmEYGn53N18UaDmjQJWlGY8CvVDh+oC9+uuQJB3f7QuzFyhBISgRL/7SRxUqo4D4d61L1
JBG5BI+ybr+k/ne7tOwj2UkBfvzvgth3kFXmThichU5qxw81tOlZUl46KsXr+UUi8CkDTyWf9l28
PBSyfdNIllZxlIfBw7jDlI3s+Vj6G5jvoJCav5pFAdHenyTKNWTROeI7Vxwx0x+TAz3/Sel2pS/G
e2zen63Sv6acNVONIdqSI1pTViLlZ0dYSoU+nvhXY5bTTVc3xRPVcksVQTUbBJxM+huSoqqhQh4Y
+RWJ/5EVOEgYGcG+E5f+HNY0KjvjWM/0BS+FnXIi9BRPgTexpQjjncUgeQv/HsVqnd9BZKNrFhB4
/ThoIieC9w75wBYlOK1W8t/rHt7KwVifC01YEX98KqnJgr18URuhbAxbjklaa0lT6uNEQRXnTccr
iEiMAx5hrfYPwI7ZPchsmyYsMLdK3pWfdunZHOY/U5tDYHQqkvhouW5o4iGDiwXmlvOPtjOM2Mq3
KiajicqtGGSNjJFr4d3b2LvD+/LcPctP6PvCrlMrohgHdXvSbKapGQHrjM2FlWvm9R7YAaZAiD+q
4mKEjP6Am85QkmZriKJzxE7wpT7uvgOX0ozmg9E9yCAgh/GhsNq1AVl0isdU+O1TcH/nqVB8eWM6
udyYLY3sVCqujEUxLI758FCg+tSoezWtcLe1TGqkdTpFtZXLwPhrqIramxs8VAadlSmyvPkYC6u1
dnaEBENXtvgl5Wam77glOl02gPc6aJSzSDs9R6Q6nZgCpB4m/93RUD+fwibqA4VYuK/P7V6I1WsV
RsPhbHp2fyqCNk0uOlHUTgMl/kOhDWUHqZ8L7fsQw0NVcqIy/XtT9J3EKM4Y7ne0alOYYV7rhnva
PzXt1vL471skbeVp39XgBFUAzskZAYJ4yNCbAYHnp3rg58LQINrb03qTRw4cPrMt0+o5llSg0XkW
IcjQ7UA98bfelMFlxiMCcVnQClg596OOT+fXEw6+ObY9NJFUc2ZHP5MjHq0GsQaHJOKEqZxnmwhy
jFLO23CjwBTtAskV2aAKH74m9fWAXhF4hT71nRz3Gd5Q046itq3uFq5TPqUXNE9CemiDCbPNI/YG
0z81AUKYC30dxdVNLR6IO1BRtMMVD0dKfD4g1hzpzBCH/oWmOK+7NL6XcMS6wWn2TUcIzr84vZCf
mOsYGypRhHS6NqKPHSSUFjlk8SpIz73a+RjHz4N0uudBtPwpTiYNKraoJOkUBMnZEBhVoX71+Mek
t8hiHGM4VGfANHHkeXwuJHOavFCpOpLiHzrvU5nsEpmuaVIxkO6psEkHWo4eYWRxdPqvrx90hKZZ
HyFULFW+4tkmnOhTEQQ2mn9WIWRMbLqtb4dA6WHejXozjc8AJxTqYFGcQdsWd1/OGo3ZVyl4SM0M
NNRCtjNIF6febtyEbkuvpfZIlr2HHTBHTvVzAWQPcGdD/eVX2KTgh6fMyaTcrrS9HV7taZ0KHtyI
xw4/xcQGauu7efs8qa9SCKudvRoaBrUf9UJjbjLtQjJf6XpPoDb93VoQ9dbDZSG9P2fpttLH5fKj
IrBmEBjZX9hXDLbV8ZikfeJJ2tpukvA1f/AhU/3oC2FyhuL8fkRdZFWjtyY76RhxfLEXybyMf6tc
bMWia9StmsOAoneePn8lK4GM8Ypg/sDTlA/Y8FH5GI1KoZDF8cJEFB88ih5b8NO5l5qD9HsqFFQ+
KPC7AVGp99OhUMGNIJROguFDoLi181DuzEoaLPTzLS+4dbhMKGKz9JzwJdGk42JMvsPDJup4MnqS
ekOM7KSRati2g6gizlV8G3lfO2begbZGkvdfnbdbUvZo8l8+1HRTb/n9Q6g/sEerdUWjw8EYvbfO
luPFv6J001yI/2HF6342a/w4BpTIy8jZ9wk9ix2QObK1sqMO/nfDG97VB0gLjcYTuPoyLoN+j+Hw
4BTi6lF3QahAbU2e9vr/xPUvPwQDWXpV3igKvXNMc2eVOQBd534vL7PVwFIMjvdEk3n4Kprdi0h2
xZY4HKyRapTIsnsg4lOBkf98TNmX28WAk/iUvxYONCrur5wRJku+8KzAyH1SZaSOvcS6Pj8OQ8+5
cEtZC83m2OYMmKYppFGzCp0llXubOrL7EdRChS7lLyeoxcBbideWAcd7i5VZIsHWIjV9/4ph8zpB
VexD9Y48eh3kY0nXKYG6DPqbbn7ImxU4HnsntiOnUJ0827tYCRGUJ8h5+lBg9Dtz5q/NjNpkw2B8
cvOZJo6jDfpcqslXBHqOt/8zQpFdiwr5VVN9qj2uQX8KyL1rZfYMNDMgIUDS+vuotDcyEm9jL+yV
iqY04qPBl7G6jOXyJu59YAx8NYi2z3G263lbqBVbEvHkr6pTMQJBTCkFu9QeY0iwgEQ4ce7zoMNh
ZosgjHuSpoKe6NKLTDYkSOu0m+eDDE5wzPmKdtWs6/0QSKnLq/fwLAHVaT5vXv5E0Za0wrhmNHjG
iZY6SsULGsMTRS60v3buBvac2A0Qglc0tqFu04P96kidhuSXGuaSItxkTw89j5tN+An+gUjq7Nxf
xTkZ0MaRKsFOc92cg888k6XUE6I3RkF3azDhoCvhb9AA4vSQ6YJBTUfspV9mKvyTGN3KMRe7j+BJ
LVcHxm+SnM6Yt8G7R2GyG34jD31vthhTc4oqO3ApWm1+XWPP2x4SUVKLiVOnI+aNjyjfrXN2vEil
OR4cACbTjs490YX+PYFCVy/8rnBJTTZqtYba5OSzuUfLy3hen4f3VL9Cu/Po0RWUuIV+6oox1Ro3
hm0gn3pSRIrYY8UMkmWqwbQivSrJQ67TJJyYVazjl1ZjDXWmXKXsKS5DFJDlO+TXXXIobGaS7Ola
ybf5tsCJmUPhr4yrZIlmkvuLYM5v5T0leNUjzhLeH02BEp/pJHDVUnfz2uXp8WK8zI8cepCkd6x0
eCuaz9QBetJq6hz100JVS+C+gzH8gKX8UoegV5O5DTCQkzjOptHmFvrA0vvGJK1JZaXv20Nx16R7
tTr/cE62Otvi/Pkt645QzR2LHWyTgBNh7ey0iSIg17kvP6/bvYf21UmrvJD9onxmJPPEBC/+DA0S
uOh/Q/dC2PwVjbXHq9iIWosFe19kgRitCovoulfuRH5gfMFN4rdGqy/ToCD0XV4AxumroquEuUWw
2JWRnOP65QU2VqN1y0X0Nv6gErCSs6AfplEJS2gw+n2bgO/lJNDMdtXdvBy/UNEQDKdQfuXsJ9fZ
KnwUIawfFA3fPyJzniayNxIR9S9ZTQA24uGo05Mx2CsRUhj5itxuODibJOS+5hWIg2QGCwBr2E9G
zsUo0IH6Jh5kjhFCq/VcyFKUPEZUuOvH1dS9dMoHfuNeRRnENqumnKwa9dEUySL7NGAzoC7ad2EA
OGKV9FuzW1pLmuT58INmKfxT4SClO9TGcNyi/U9daW6N24wJGhl9Nl4HKT6gR6W4Hh8FL/vbM7V0
RkEyxlLdSDC2CUth3tEiscbBVJRyjnEbskPmrfp/KnIEST7MjJdbyeE/UenRMhjO6FKl4i6sNeAt
8JLCxYOqdDHGUBbYeEfH/yaR1ynzphvKaXHGFkz7k6U98WTw1x7yc9TmW+f+Kjzmh/53pFKC1wll
3hSCuXp3ZWYHTIlaSN4VGz5gvL6tw34GF9Xe1W0kxY4Em64RDNFc/SY4HGIm8gxFRahbkY0NFBKG
MibUUKnLZCuO4roPid6OLE/smcis2/LJ+zqb1w9VJFYlUMTCjEe18Rrrq32eA2pHrFBTS4lU3iK3
9nmtGffJQDRMZD2C3KbKQ4t1dTo7SLmp0/CpQdOUlZeqxXPF2AATL/o+CtlFzhuHByGHCC2q8vOo
IhX8EbC9AejnTFsh+kzReY5wEKE3m8sw7Zk8QulcmLZcE3ZZ4FYN/UV1lQ4inkhf2CZSxtz3VbjJ
xr3+DXTIfV7KWGu9SORhLax/hlEYzg94M680Pp3XVn697PjR0JmUWbq47MUAkoxuMYo6xOvSJ+T+
Tqssbl0eWKKbsRvp8ZJaCfflJhIBpR5wVuzaa8tYRODtIiucFoJ2rpnT5nDxfLHQakzRFaK07xae
EmRxr8jmk2MDnX5YbNjeKkCIgcKo3VU2NpvLA+YtmQYzuwXI79oJBYLagMLtCPZdRBTl1W2fVt9X
0lCTaS0JqtTQzTe7TBCxQaVywG4t4wmX9iz6trHZvWS2XwF4Np/ZRBxEqXhiqhVClFwQViBYsFUl
1oIzMO4V/RwtSjazQLwupuvH7fN2ZGbrllxF4xPRzMUfJT9r3PJ0XYZEUChMfEfCIvX762OloZ3r
B1eo4TmwTzp4gbS3CGMRR8wb40G9Re6l6Y7lX+y3Sdu0gQNAWHVZFqa8kBnIco5sfnxosFQfhI4K
36ToB/IohAghUD7cRHSI3KtWnyj609rJIlzQBEd7SvfpZWz/d8Pq1nCWgcTPZLv3ttQIagC/kUPt
HPxYj2qpcTXUND6tTFaiogob3Fa6YF/i+1UNN3rod9hynPvCcp4IEhmAd0UZZy9PbaVSSUTq3bmX
dxqdpZHmKhi2a3NzH2S+3NM7l/6LLTGP+vcwUsH+UtJOfSqXmylmcODATr9PD14Fdxurov38xFtB
Apm5vGWc6Ite+9nY6DzKwhWijDXsbjwMV6E/R/J39IxeNGscVKHeNmhHU9bEdgLOJHgdPUfqzV68
nOZCMiA2h2zvWuwPwbvqLau1D6v1Pio5MVk/eqw2IJ1q/5OGukAd2pvO6scTbhd8TnKX36zQZIcM
tiqr0yepOhvqrIz/sHR1jbUyh4u1fUpe4VIQhdNYb1LJMZLQbEeD5xRAoMV21IjzPxJfNqJT8OR/
aWbEefjZ6fKLjG45BEq+YVOL1bWSYTAalbIiONPzr5tumdNvL0hxaoBAghFgu5xaYe8fVf2ClolG
JUMapm9PSDtV+1J3BQ+k7spHDtA+82gz88nWisHT6+lrthsDfDJnENowc7Tsw785+OYNjZPNKlvh
DgrLTcoQK6Ft7mdVAUmr862N2KW1pRw4C8gUghOX5AyUtIUiLgpuZ9i09p4+t8Irc4p2qHKWB/aj
eBgEW5jgrAqyBnsgo1PG3WP1VzdSDq72dj1GRoFcwjTXzJ11b3cmLWnxVSZRchYckzBJYxccXgCJ
ePJIFxvTzFUoYGSqk5rds8b7V77El2oyZb2+/gXBN0MNzl8CvtRmk88TZ5qQnUNJRB9OCbyE7+3m
46tMMgwwDFTJPtZ7UJllADZJxkiEeiegjD2r0fIMzZBKTbXQLMBthK3y5/TuNxA/rMCdir+rGbL7
RnAqg+ZPMBB+apwUL1umqLLlWY4tsIWba31rE2w1aShMaH1uMLEyQlyiOBuaVbfWVXgXJ/LddXV5
WW51VSAhmzwv8oFfqFQWCl/8rHEYZI/sZgkUSy0CjCtNIiKY/x/joGd84hEoPIQuChMvO7p4fq7a
S0JZ0zOVj1Jgd0T/TJEkR3mPwACL03xpnVm7VvzgqnyA8xfQ+75m4l57ZfUBSpUegPnF2Y206T05
V4lwFqo8UPmlG27PHYrjvvkw8l0Ze7cFNK3qKVHANHl6xMwTS9CmsKxVf2pS/s1nZQMzw2HbUenS
z9FYBP0AMr0QDRiWIHCxQ9y20vWykb+v+FoEwDjq/SVK/QKr2tjXPiP6U8fJou4g/DP2tPrifWkH
rUYt7Ju8W3A9L4Ajd/5eGTCKHJaPdfZ8NG5+3KLqmWjtc4fODDrYRmS/LesuDaIe4Ll1q8kljln7
6zS7ZKg3vWSrSWVP0wBKUrHjriiuVNgVNlCLZ1hNH/u7kPiqys6ekNWeb1S9ZhseEayeroRkIjzA
dMMkXAfrzoBrYKxJdFLbW03wA4cIeKafG2peJHMtU4nlp++825HU6rnvRxzOEOsvYIqhl8ankE35
/xqKt8OR3YLYrlq+9pLY02Bgb/N1pqY6NRpUyCkafWPZz2ChPqpNXSNxPxAg42z7QlyjCWXkCGYW
9MDXMNdaDY0qhJWPBhxpFBcS2Q+UcYQGZnHgVyoi6T9RN9yvxTyPpm8FEzyXt0vqj0amvMKXnSTf
I8ukby9xBakQJ0h1Gm43Hh8Wc51I+Gkrm7yipkCXgJBMsrDIG07snERjy+1ACGwf8FPVbUutgfoj
rOktvyuXtmmICry6Yfa78vvZ2HoRrTEKSG+hmLAzDd5lV75GtEXVctqIxeBP4OTV63O0/apKqlOx
sjqffiPSXWYpiggDgjeX2MTkSnQZgWYiMvX2/Hongo5mCs6s6XYiamZBvTwQoqLZcjcviUd7itDN
r+RsXEPAXcmfdqE9J1lcbsQCt0jjbLLI0Xms0r0rkOsUUQHil90HUcTww0phGuXrz4dQIeDI4IT+
9m9kf/coWKw4LRH8ij+lx8r8zV7zwsAazOLFyJKR67z7S5bNgFAEk9wMpNS2E5nSnk/DJxBFCbHM
pJ+C1/RRrdTJt+/kDZulcE6H5cuuGK0tEnEp9jAIG3Wr4G5oZ0MEIvn1tZP3VONbW6fnnLts8idH
0rIvexecFUnymV3MvlUPJUnTdjCKK7+sjZ+RHOxTK4D0A1L+haxd8YrslB0oohG5xTvZt/COd7R+
CmRfh9K5XQJn3YPFhMZ5JYUj5NN1WpAur1PSykSS2jCyLgLsfQ94FkEzjkoKWtUPbCL16vdLoN+J
obMgAaHGZWiUXi5DkzAxitvPYwqgLfYwYf5zXYd0RiTrXsEMTXucQhHvxE3q+KUi1S2NDUZtuzCh
qQixykzYZUbMVYUa5jwDRAT3/LpDqGgZoA5C+OMttEKOeuB5ERNds7FLfIjwIQLh2nIhCNy0M/RD
nehWbqCTCngypHhaMXpbkaME7dteWDYsu+56hrm54jP9pEIT5N1u8suOUHPO11UI31cjsz3cLjwd
r7NIMAu0PYRciDt1qK+N4IAflg5czeO3vPKWfs141gwI9izgdIizQzfOFwU14a8s9plUyU59v8vF
VCPw2zQT2FwFIOMkUb3Vc+7rfX+mdHJyPRyKqPfHo8D4utaxDkUk0uNLAcRKbs4Gm3kC46vExQpJ
GsuEvXrRKJ8ZFgmLzI3Gn64U0OjXoDLUkpJTI6XCwuHTAWmkp9046uxRmbVDhGdHD2acGEghT4rw
6RRMrE5bVc7JBNZI+FSSBVjtj0KfQjlSSfBpvzRkWYuOaBx1VnsjPKOmwWqU7CrudGouQSMLyNSf
OiveqWorluFrLbUYZRzW1H1Q5mPaZAN6SRrIJgIAN8h7SRIWFG4Kxc/leVjir8dV+STK56eXJIV3
oWvQTX/6x7F6sUdS+cEO8pAUVS+COaa5sA4PVGQQtKJPE5GCf7lDrwTMeRA2PkfvEeFEOO3zwVcO
zJhZgoUJqLebzZwacg/QflIhMwbhUGvWe49tfsfQ+wKwIpgy4FLaF5ILqK/e+2uCeaVPMWcl8RjI
p6wUTE/pHuXuBfBFLI03j+Oxn7aB1QifU/Y0h7KH7JXu2Bk7LtYi9q2FWvJhZB0Z4qN4mQZtrLB5
m8psrKc1WDgaoX48H+N8gr+QTBB/02zlO4kvbN6owanWn0Hvi3q1SVf+lY06gd4OZD9lPVUaAHzd
lXdACjjNJny8xmqeXYTW7rs5aRyUgjA6Z/g1iDtH3sDrgtdxphLfY7POYMfskMjTfL52Qz7MLfK1
dXvsopYDbrkULN5aih1bDc3+5RDQgfog0HmWmIVdWzJXJhERAgxdN5lVGteikY2XBlQnP/mtn2L6
6hTAIV7jcxOk0QKpUndGCF4oa7vfPuL1fzyUAamqduwjcUor4YqJFVza8qNd3+M0YCEUgiYicuGd
EPWaKWVdWIvJTO89dXHlRAzHhT1oOvZKZJiH2HWaEMriLABTHXyDgctJUVjCkHfC15dqKzspWXhw
VGLskmFYT3AwTb8Xdxp8DT1dIPB2ugovHKGiXCvFVkYmkG+ajD5ublO3k6vivGzmfWYYpxSgGCh9
K/VX/zpr9II4v8mXM7HSF7sfp+M4ma+YkfbFWa0M3VHgMGjihtF6vktGcV/V2sE9keQ9mtI6v2m8
lhDcvgkg7V3ie4Y5O7zmznEvwv62JaaQEYpzdDwQCaD6gxbuWszUzgS6z5LwknSuNrizKj5wyThA
hCRUAVOHRzMnxXrDRHRQhv5lS2ARAEJYdSxtH8yzNl/CYJhW5ZQqEZWPSDLkJn2u6qaeHYRpUko1
MM+YAsUKLZjg5FOkNMrTUOm4za/Vh/zTuTRgMjB+3kU13hns7BVSz1py4S3zMuGhNDjFj48ergps
nryAZQMD9DD7bcwEQpUwTnIbPwGeoShKKWbMP72FLmNpjOkgW2KfeJOiWduOFiwMcH4eYKYmMvGq
Pie/40W+UvyJEqXngOGGbIiwAMwL1Yupy7WmfDf3kSVpimcOuL5tJPMv8rJSDdvVllO7uKYmTL6U
2oKjsP9h9LJnDHlNfBsY+oJHO5dksu5+9iXD9SCTB3Yxmx5ec66pgw23RdrQ9+uOcFesxWRBqe21
0Jspl8cn5enoAnlYS5jqAcM6mY4+oo3N7vNdEqKhGRrDeN1LMEKZz17QBLA+gAWIxo4bc1PaxOqy
NiVSYaatLDEMf2eZFQMLefP0OVgw3CXoVZdRIkHcJHijK0o0GIsq3HZKJL7G2T2C5VQbXvOA6hiO
mM6JikWUagJ5+kZKow+9DEd+7uIKwHUV/B0l1K86FaO/MCIM2okzsEzRHucnaB0R3ctxMP9Ktyr6
8237B+0HYSAAZyFMuyitd5QUcBoT9svzuEPWTDqIq11l21g3ZKV//BS4QLsrLK41OMfJ61/XB+Hb
Lijw4fKx+ORim13TlYqZLguUaDqtoQbAejC7ddyHKZgj9q9mV6v5q14y3yhHhfmmiW5atlTDS1fV
DyIJ1DY5PO1VRGoz+8GqE63PeMDUcsam3S8sMwKKF/NlZ4+5EeYU7/uy9dBSgNhQuJjlVTUOcEzs
b9KEpw3jj1Fb0v5Dbckf9tO0Hp9ywbulyWVIbOVm/K8FDbCgCcqLbB/OoJOVwo5I+ZNNb0BQ1zjP
S98IK1G7K/iFQ+4HBkD53yUsqnF5Fzd29cNe1f5OTVOWX9xK5m2b+pUlLaLlNdIPyUC/FZcF9qOi
IjYQxfdunJkm7ThCzysSEW33odDjCG5cEZolaefPpJwtHeO0BVCfspbnL3BQw4nMjw+fq/gypbNE
IXFaZl6EUHDmSIgEgD3m8mJ6ZpwOH5IE583j3aJFqSfOS+9V/mTxvMeAtGcoO4Jlhos6nRJPYCQ1
fNNnsvrktCbVymmFpDIGjAe1JOE60YROA+EV0Vv3gyF0KKzx0lGh1Jo8/cvsgGcyPXE6GwLridpS
zHRz4gFZsVTLLdoaQPLVMynLeAgT2/nNU3AoSPkOxhqpv+9iancqCsc7zzhaLBXeZnC9wtF3XKT9
+xWkSTd8AbBIkjWPZk6fxqRZM7CG5mzkOV1ZPGbi26WVjmO4AvKHnerRZVXBvMxKjPav5ZE7Dx39
Yi0mi5ZepAK6F5Fsqd5xUQ8wzYKMswVKjhZHxiIojfMt1OCB5TBmQ1EgnEbFO6U+JzLhzm407Oq/
cRt666lWztiMa+Ny6XaZsA3gCay42/xqJS0l7guMHldhigcb3W3LvSEDAY4ho39LNMjKU01l1ETt
TGiRCQd5ijd7Y4jHYUFJP0u9oyHX5lQ7X5r13q0g+0ISlZWo9bsKflRDE5NtGTHbu/jzvAevERks
X7aGTgS3LgBNk1rIkZhq3Wj/+wmwVrCsv8HsUPMgNdUBPirXDriofyuj7UPokWvmt7Lv66aobYk2
YToDswLgPtSnqh3IFjvn65WzTQCkdKjevyAIwVM3rekQhzSN4Wawcg4b6hECpBnfSYanNEyUTb7i
YN/vBSAsUaliaX7OVn6SXtn3SmlowElarHp+gX50H3lzwWPTH3Q/litUejs9UZGoI7cIhpfihC6k
78SAVEDhwYUI7EQI2gLHCoSQCx/pLXIbpXNYu47CN/e393VE5XC/5L5tAtod5pcsjf81aUELvxX1
Dvsl5FJlZkKEidBeL0LEMs6O4MRPtUs+8FdbMJdsaY76E5EpG9O8n1REcwpU3rVzc44CFkF2/3Co
5lF42Ft7UU85XbsfwdySUuqJNZ4KgAjrqSdHHJZuepLfhEwwHYItNBU8OKJolptoF8B3ga7RzUmM
7Xfa4OM3EOJabLsNSFnmO8kcApiTVVaMEZJsmRmuOcMYhBuCQsXjl/FMzwtwExBjST0xC4H1dK26
4HVtvV9B2fyHMReGVtZ/Sf124KoPbdOAa8/xL81B6+gGfpdbWnZTaSGmJmu4XEdN4W2XizQDcbUG
AItyJzScU5OSuxNcUU6e3lv3D2g2tccJ20l8GhOAn+3vIrBaJ49iYNWDm9WE5yJl+2s0r2UweZXa
axYoIONu15Yg05qLqAMO7MK9AbHoY8W3NvpPHhqrmHsJoXkM6fRN6hCmJUTovJyQs3507kOh2AJ2
jVPipUDh2UbCgsEvYA6mMl0caiXigZovXDXMhJPajd47Q0iNNnksgRFCfBNd2njCObB11BFB+eJa
1hbjtgDqJ/o7vDlcNk79V0CKN/MS++Vm9dElWJXOM8WWC79JgqIWUcTDd4zHHinp6FKds+VY+ABB
cyW5cgu+6WwYgqKrWNV1aWFFwOjkwahthK5cKHoncyYJ4FFw1LNCiiGApRzipyecPrxBeG/Efozq
A0GmDpWYwXAE8TN8fWBhbsEhDkVc00UYLC8Jdw8fj/shwAK4b4GKxt4sFuUBpSDHEOa5DXiZJ43H
HYBxzSZJjbn/lxXoWv4Aqy/hxVoHuSsbeLT7NNWc/MmLbtnFCj70yXWBQhAU/Rl0HiWVavLXR1R0
xmO8Lju8Vlel56nI7V0f575ibQjSQDoHaLxTxH2q6VPAHXyd9a4X2kWZbBtEpxxvCKuK2KRcNyaM
S4AXk8IJUywOJqFoqE+a2xydHWkrV0+7bnn81avIOvm2aQGKU1V9WFPz/JRqAqbD2wLtzdt85X1l
BRzsEMT0s3qYl3qY5+QrVdOX4vK0ZinLiqbcKIlEJKtmrw1ke7rSFjZv3Hqxss5f43foKOU/O2CB
t0ZFL27a1KDozHLOXhnrXtIuwWz47eEmMzaiUTV6q462S1Ll6pabEgLD2b//Vo/ASoaAWKOagmLG
5c96eK9rmQY8JzRvKMmpGMNrHH6zGknzpzCHXJomVrPNR7KQxeZ3C0oEWqyQWOJNIJxaCV3M9DTI
pG4BFd/AH7ZhCAMyvF4riZmY48riKtTD1/AQxPPZAweX+wph5sJzeIUs8qRnYIXHSu7WlZUCTRdZ
cW2DUPxZvaVWk3O/ZzpL0PvIpDy4Pn8gQ/0fEy/6w1RDr+ZdizG7I339goAqiBO2FDDgdAQ1NH/Q
VG0i2s6sBmKb5mcJs//VPkHkfybHynUwznlLVKYu0PVyR2GwS5XwfSo+Z49CyqmjleDfN48ZxSaN
ymK528/zTBX2URZUjbfOVLNp/abLduLb5WzIaaBndo8tW/dMPB+w1K4lqGsbd84ZGQyz90L9LaiK
IlBSbahq3xlcVg3TWhTZRqvYzf3sGGYnesAPAaXn7TE9Mdn/lBs5wEVhLBt2+aI5QP0wWRiqmjtF
qJkGabf7SO6RmQ1Emv5I4DzocjlbQHNgFpTanhsr2ZSBBUt+DxDk2D4jPyug4g889f3L8oA/Tqdt
OKBn8hZ2G7SsAtIljyf3YnnAvweGZS1e1ElBlmOMYMMnHuPNmlZlLColgbhUcCTE66z0F8UTLKIZ
0+tEQH36y4XjSRUrtnUxqwi3j3Gn8DGvBG5jO+0tnwzMpjgR+UfLKYnw2QQ7/aWKDB9LflfDxFEn
GytwuEJEDzWE71ZqwkLSYwDeGiOetJI1eaxFHWPD+o0UKcpL9y8dDwQyaIBUBCVdX3e99JFkhGoS
D+oUjZEYQvw7ax9HQ/Dh0rtBNE1pvHsywSfJXYdeXrqzas4AA98TtRd4XBD7MemAE+CLSbfciuAu
IyU6Z9/Q/B6CcU0KgYNBdvbQksnMuIGeEDZ34/nKAOKpl3lFNXlnhnMmlzBNnoW8gYP6hqWbi9of
wv0V0HS8TMs7MYU8dm1Q516UdUjQwWmUS8lEDUpIxZ8BSyC3bRDb2zD31M/1T9E/YrbSem0zbMFZ
4vdfCqzAplpT4dsuYJVRPzGfLk5fxmCw+zHeJ9IBbz9xmKILP3FpUd7rv/PZ4t/sV+tb4JDnWTvv
Gj26onpjvabyA7B44OPLR+RcOWpIg6sLPkWtgIMEm8HPLt3D+j7xZvi3P8iCLB0mE6QijTkRyRzt
aSjhUnH7nSsX4l0XLlgBNikDsxpCgBJc2LN1uAOv0bjOWF/3UcAlOv3K6e7C2wEXbtwNlAVkNyed
Y05FL61sHV0zdzGG8IXcVq2jog9xSCvxngTVdc8GFBo3wFm8HRVhvwc0ROjcdnlaB4xHIsSPSzfg
HexRK7Mh/d9SfNK9ZKhVB5vS7bc4xFTFaLH6xK1rCiN8//v8CKV0/rQYVHnW9xuwpiLes+esEBoW
F9W4eor5Km2ggw8abhj/f/MA+BcpO8VA1wBN6klDgvZEdDxW0Ac4c5v8MyfWZJEUai9KUXEpwiRS
WPrvSSob0yGuWCFgeu4TvJnjV6TyYSfeN2F7tp9BDItiUt01sISek1xuKUo0gCfIOk7+onSOjWV9
ANUPQ48cy89mbDBqZJe+kegTPygMy8K4FQzyU8ciKDP0i3pVwk0je+JsWD0FWTGwOn4dYEaeXOol
rziJ6wr4ItCIbWQ/BevK8RNVoDUOjU3HbsLVbWkMW4JNE0loWzIjadI5ESG6E9JhDYuX4FlwiOOe
aYjZWXIuXvFek03RhsLcGLozGVsGw5uluXV6hhSaK4DxTMSFCCs7uI1HHzE/+4Lzj+vS7rvO/s79
1ygpuXdxvb4mEHwJOnFIj7g/MnNZrEH1ystqNNl1Hw4NqHPhcessAjBuDJ+6s2KPGHNegxI1trBW
tZ520sji5qjIcdR3pmnRSwwgINLhZBe3KK+9R5UjVdMh491JZVtU9kVRkO6dfvrupV71PE4MlTdm
Ef11V011DcMISm/7ZhLYAAtGkS0RS5wlZDiKqoUne1EvCFdbHZK7TgSzmaIXv+zH/2gDLlMSB5Ce
RYUL/lVXdcA91JUECiz2uqz2gi1VOo7EE5Kic0W5GnwOA3s4uD+SW32NhkZavQKfO+/DgwahigRI
ORevsa70wbwtS0tDuNACl3r/MFS3KyP/y5WQCMToAXOKGb8j2TCqT9gbK9nJ2z2gAZJvsXdJRjHy
YLCU4g4yeyGeKMN4Wa4UoV9zGggBZv37Gl8ee5X4qvLno88/SZkO8/VN6diORyEf26G6qg3aol1E
fAR68zIN9WmR42L485k2CLvon1jbfm6M+AOkAIkIhGCgMnBAi1zRrEEYa4YiwZKSxB4++2ZtipKG
AdYUHBU3bKPFAVLbploBjLLZAmabyh0kyboqRYldHzwks8YOTuiVvC6+F/5pBBwUMFa6OIsZWsXM
tKfpa/3z2SjUSPiy+rkyMeBJiqgreEpr6LoFhLunEPUw00AdaYx26fYm6B6OnVv8cNcbNEUsdW9P
jPEgFPh/pAgDxCD0TDWRilrECOatc1k0r6dl8I0ezlccStqwrUKI+NV/fum7C9k9FxtA7wWYNOfo
ySewRgORT7DvPQ9yxnhHTq1h4JjLGnA5Zw+PMxZkIBXlrGgOah7HnfV3QJaslKVnbjGmQ0ghEN2U
gDIeM6ZceYQzKBr4TkfPoOsuNlgT38Juef+9pmI9tgaQL7YCl67rDB33kkaZWpH19Ak0XWlOOvfl
yKXiDPiIGJZIoypECYHhyFgW5qBZyNU+BVRzz9xv9V9D7b4bkes/RPnIWNweiSDin3nZ/Fe9AOZP
AXTJrZUpstHP54PP3RJCa3GNj0gfsT9/+QhXKGbt0JSV0Xu+QH8Fs/Vcv477SxafAq5hpASCYmJd
MYkmm1ICEu9wN8/CMYjJwCJs8Ab+ut6WqyknvEATO3kR0MoikOPIFdEH0MGOgXnwUf6InTpflhC3
DnPclhab2Pn/tmI1vt6Pu5mf6c4bQQqwgeV8tIylav/onsHuduiVmSBmxMpl5kBNhTwb2tD4MH6p
g0zclFA40lRBelrMxYSZD3uEDYLhCR+pizYkn1D4lLKlCWyobwSRKR3QY8raGHB59vN2EP/Rbkqh
HhfqJFC9ROQKwdCeSIpRFFLVWhG+vHOaqHWRjwO0NA0CEEYLgr+B2qyERGWT0ufNWAJjqRHnDavz
u4Lveox76KqspATWcVOE1QbQEEyUWZ504bR9OD3mp4to1e2ehM6eXR5VvW6FT0bd+lR9WPydNCt/
nrv7puYYXpF5qPTT89kXagz58fvS+M1kYoKefVimCxJ+sWP99TqGa4Ohi/asmGgNuSSicRjGEnqS
2wWHqpjDcbIs0xgSaLCSsyZ+dQC8WHwCWa41/hFMsmffjd8WjSalvVGOjxZRhW39lucgJ5Y1QAYr
f677+7XrSNdU5WlVTeBv+Hb8OYztmroeRKTzaU1GqLIri7lH6iP35iqbZZh8Zyxx8EDxLDYfo+1d
yEEA14gUGhU+z+NYT1Q0whrJxZk6tvRt1GSJcnx88jMBILeltdQSPQs82SaHWgO0EbtqRcmamh1y
uHhwglbKsI/6WXL52lLUlvzx4nDnKAygtO+hvzr50Ytlycgi6osT33N8awo6cKMttivcginefHob
+gR+wzoHGDaauU7W/vnQDPGuNIlTNayuLwXlkiCayLGNt3qw+EcDdl5llDt3KjpX6u/ok1ir+cvP
ws+T01rFzrgt9kmqrqVjGGe+i+FC5YokyiBz8yDWpOtgwCftLMeM0V7E85YVZt5BaXUKkcFn0oH3
VhfVyfRh7v/13Z7m7sbP9yO03kBO+3b/kweDsxonU7+WMr6vwlsDQWzR7xICK7kTOv+0bY92YPpY
VE3RULWeNn2/sBPkGkRrkuPObXRVK1/++LSPDTSwUPggPtHLSnH7N4I7J74UHzAqA9axDC88+o47
r3XQUkT8QxyF9kWEy5/XiHYbyExo4a4FiD93BxM0GaqTkzyhxiUncGhwQXxYhRWzLieT9ZJp0e2T
u9rEkfAECxfN17qSKM2fAgLYoOH5zsv5qf01ARcg8S/raoF6Btk3DOKRHOU0hCEXRFrJh9xeqX4r
8vhMvu/SOBI3EEXatGOxfe2y/KTdlrD0+BuKIP5pdTcd/KR1haAK4jM43CTaAmaDx/Nw6Ay/B+p3
ZblVYgJRPHcCiGjU0IlvF/edSflSIEmYOTtpH9jFEmW9ZNQ7GELUQgcrmprr9Nz+96pi6M9I1dD7
JLWLatkCRao6J0PrttBamHCaOYP3JyC1FmJ/mXBnMlLUCz7WzeL9SoX+yYplRS5N9MuK1/y4LEwA
iFWwz7qzbTfA7D2l9q3F6zOpHzN0N97q/xFXIh9+km7VI6WGKRTCj+UXpuB0ydNI3cm/5lZgyAkv
tgifQYbiQCQ6coIu1Qt5ucrFGkOzqPOwHlXbfE26hxDn6FdQo3evpY6qUVw5yAxkAJyOjse0oCBX
2pWJjnPM+ZeJ5JQAoU6XLnwn86EpOxUSfYSJC3cP9aoHKtELTnKI9Pw4vv/CQGt8gABysJc5SH2U
hONYw3INJvqQE/0TJr1dPO4cEd+wbIbi54Aq1CxI8ln9LRZDvyrHr6GwABpJG0Bvr9jJnXxKMNWF
KPN/8d9bAWi+7iJEO17gt3XPSE4qAU0vo5Y8zyob9w18U57XSPfPK8aL4/qUraiccgNel8BtNPYf
IBnuH6cpTsfsL3K5yuEK7tlSkbM8Bqzx1w6nZeh3wiPu2dDfYbWgNrQ5vrY/qu+VUB+LurMPyMks
JandBna2iebOGs9atmntmaA95tuBAyXu70HV8WwM1H7dcq+hEtWQYAqCHNWzObqxyiGdHw8JHVAT
84qhEfKd6yMtG6W2KO9b8TRRCt4s5a6zcfexIY5ocFCqedNPUHZxA+EpA8XqRVMN/Eqg8mbWtLmm
CP3myPRsnoAJTeu0kmqV6sZUIIYeXDX+4HGBAGo6OCrguiOf9Ploutuughn6e7WZLVkLxGIgDHgy
PNDKaoqkgKxo2Xc1tY/N52j2d8Z/s7M8vJELi2C0GiL5Ioc96WAgiIwYfsyLqUgLYHtlwo+qg42V
zEtDNa3+5KcOSNUYUQ8g2Ue2tUq6mlfs0071iqbC1gGekj9T0vh3u/dxPq3I4iN33fZkrPJ86KT0
MxuE7e8xMgXpMs+7lcMEqgPGtcgDP1oGAH4Mj/MHz3dY1Bgr3c9jMPI1dIvcRkj533iFZnW5C4TH
vSu90RLp5/FcLOdWgLHU4DB5Ar/ZZqETRHUZ9/Qj8Pl7NniXvzpg2U60OqH8XRT334BWzlyf5YbH
3tQuVpiBCg0otHApXunS0zaUkmeyR0xL/ff9HDg5BnBqWnzdRuUIuFwZPDNCeHqSzzYTJ8jz5rVR
unAp7gxFMFbw26IjeStTLbLSYPTalOTHOfKL2QNir4AuOaKL5nzyJD858mHwyJgHUfIr0zV4NM8D
dnzfxrn4ZYXiBRxsYJj2iQ2dri3fhpclyb+LEy3atp3bWKfN7ShR+qRi8lAhcPy9Dy23ioRA1haW
ruvAnxms/ez3vLB2YrbWZG8xV4nBGP50hjhanzp5TgYdbHt7OOJFqnBXndRQ0Rn4XeSE5Y4ZNErm
xS3QWWyZsrSk7DbKjjUIchEPpl6lwhRo92tzfx7BsKMapOri1xYfvBAxgcfXJPNfQXZelUeHUovl
GTqckBIRxr1l8Pw2zTF7cMybR2PhPn0VryHq+7uaxhr+Hfr+8wVDp6sCW/7p3K0YUH4FLwlRr0FY
ccuEg26WCru0leRQ+GL3P9JtCSIRm/kHd85CaS4eJQUzPx2Yfx/ckkwrMiLbAmtofs0KI8iL6utR
NPYiuYJGusQ/cXb9pPPcOkjzuRLypKieBQlqBKW5h3Bp8n0qGPeCHkOr+KvyMlO4IPzCm9PMfC5z
2DY3xR/anZtmK/bJ7UGV1cJu47fQwcbtl5z+y7YdlAAD2MVv3taxzm+aI6wnQxGG9TajZgYrmTZY
ViXS1FzjWLm7uyacvSC7DiWIK6Pu0bWxc2WoXefu8OCsfgZZ4FWAws0wGKfEmob+9sMhVAXvLe3f
+bYIH832+mMuo7m1Hmepd41t94G+T03kziXciH7I0gCLVPkoki6I9EHVmhH58nUcpOn5vPB9aKJ4
/zH3iTCHqGh/xSrXKN3Os5zC6O183aJ6Sf47KtUwCwSXRNnAgabol1FHrrHjjUDgEZkKMrxoJhG2
ElTfhkhEkh6pSrQ2q3hWw3PLzt7ty8vAZfhXOySAbmzH5WbgefLC0zGgTVqr7h480n/wXPnuwrnV
QHaM3nk3w/4J3i8fFChzwFKb2fQSvdliqR1tuC0d34qdBoOOlwod+++YKN7nffKqnOUq3zSLLd8I
rv9uuW4HFe4H9WmR+6byYE1SVFXNHM9vYdqFYVUaZJI+V/8Ux7+5vpLYhEps6/mccu1LfArRIR1V
ndeZtTM72AlQhNDZRtmxOwI8UWltKm+sdOhLshiq6ZHKi1nBUjAOLjNSNsZhmTrdHB3Bw3Dnp97a
+QyrKqYh+DSNc56Jesl4sr84/BHm8YfR3kSyAUpZoz02fkGLF76R4G02OCd48unfX44OvlhPteXv
7MdBd3kl7B9o+MYTUZkNRnMCsqpmz0xL2OMa4VnrQGrdRV2T4WDCqQz2Ps3YDtV0Ru+BryFzqbQr
GS6lhPLacOfJ1hsSZ2oS7iVJYs+BBn8FEmBG08leoiB2Xm4Gf/dyals+O9XJM5nDBt+IGLfPolM1
Vu755DBFjXFSz5n8ZeXWTxTWhTjvupzrcDuCOxdmMsjLTfxKfWmRTjQN/Ot23v+OJGN47jBEg2bp
53RAqQBvJccn6UhKbIiSvTGnfHqLdkpfIqgZQ3IhapcLGO4x9o1djrjL+ojTdNkQNnegxRtT4ono
MU5NMxOomKC4PCGHkuBkN//sjSAPVN7CbKKcsV1qmwuczCxs8X3kv/t5v7U6cTr/GNoxo2bVdtkp
Xgw9XoeyGZYvrs0eojVKPaWHdRvsO+99AP5nA5lQ3z4VrQDK89ckolZxIy7C6YiaKAiD82aDTeKP
vStbm8c+9zw8Co0ASkI2nAR1oWeEN4jumxQxdKpU64VrhUJCBXGILMx/FrMz0I+LcDdZ1qQsXUCt
zf90M7fj7HIR1KaXTIqV30mZErdWz5dTyTrp0lMTYh3fh2pLX8nayxvfjbjsLh594+tlfCVmPNao
5E+gfeA5e97d47MkYZyduKbdAR6PDqpZRtev5Ra4QAnSc0hnTvaTIZrlLsW34QdUi4vR2StcPJwi
K0ZhiK+bhVefNA7tWrKKmX5LECErHbghD63N6t+UbrZlPZfTWWaX0L4W8FP5LwPdaa8g6CSTBIPt
jZFZdLEBigPK1f/fbra/7oel33V9ML/7yH2RaXR2gv8lP49pd0eXJVH8SzcW1SxlRgQ3IMjscHG9
05CXsIagSZYfWNoW1v9O/0S+6UvLyMslLukF8HGVIJKKGmNSpGR1bOpzCrwKrpe3mNGq5ix6P8Xm
74YeG4MdRQke0exA6trD58YlXqoMjWD3d+TfwR7Gsn6WeW/8DJ8pEyVVuuV1FfFWrRd5zGhnBUhX
WWzI4ZPlTLIShDcebKzTCBlEfTWftI4ktl3+vsSjlSu+3VpMjFetEln3Pqutziwd70uvgUiiR/Hs
Ulh+cY5Ed6c4GfQOLD92Xpa0ILBP8p4zj+I5k9t70tOtSqNfzWU4FwpSFhnosJibdTiqw5ksWV/C
B3jrnbt+ULHVb/2khwf2e9IgTa8wHkTxyFv1G5FOF7rNK/MNwG7o49vWq6ykMYyniVHXXjj+Chio
5bvOkYTIugX6LiHPJ7c+dIoiI0mNxJxGLNzCBPRNPAynlbHOpgIsELcSa0wWt2BM3zFxalWh6ZM9
10bVURp5vYebmnJ8aKQ4o0bhW797xfrpyhtj/VQ49Nq0G+eT2keoH7uj8eT1p9JALsx7wup2qOg7
OgbkWFY2d3v19OycrLAFkEeYT926imXL3ksVrFFPqIFf7el+h9oi8JxURMMMImnQTAMITxbE+Mu8
W9+pS1hAFhRc8oEvdyg2HfTZjetE+mSvSo7uRIG1RNYduhCWFhIW9eYpTs+g/ldxM74cxOY8ZtSs
aQDFTB/sohexVyuAP4oRHbGtuYVBWm+DGvw3Ism2a1joKvpq/sLA+4cCED8oEIc2/f3kJ9PQqStl
QHKy4RqgYjukmHzLmGrsXJPBzyrgXA4r0N0v5IMBQXAptxZCG0gHY3jreMPJhLfucK8IZcvFz1WJ
Uh+ZtvZtM1zbM8yq7BmnLU9tqjnjqe/JdAMXJjiIoN/8P+egKFmNAOc5oFUj7ibnhqpR9OBJRLeY
KbpI8Q5zWVI2bKwAAc71jABGSi2OZU4swQcwZdekET7RONQHpGuH9uL4kqRKAhGCCXyEjjzpe7uG
C+Rqf2smnXSmHVQpiUHGRnmL161Gp/Px7/HE0pkuK5CJ6MJwSFQcL9OzYZMZSbqtq3MVge2tQ++E
szcb2Qb57B8vMiWo7M8NWmfHperx3fjZuxRgddqHy24BRg09Fuyc3+58VHOhftaA0JlK646c5bwh
9gER5nskyODwvN7KPtAOzll4OhDZ5Y7ZMxZR1wSpWrTTsz2W/I05w3dHA7YkMwmYnJPY9mmnhhnr
0JLZKomus1UHZ9vj77dfYicd0Z4cwAcPQ1d89Yj03DPg31ewyIvYPeqHmXDvlgUlBstJBswsDxGo
x1ImDsLQbfTNyUIgKdVO+WNZSTarbq1X34B/9F5po6+VPMjUyNW3mvYUu/poCEnH9QQZPjbcL6T5
gs5VAMMS9PVW7MyHNM5nzhwuJLcDeDFy0DMikCxfgAgH/wUZF2zhhM+2AmztBw476v5DOkJOMOdK
0HlyiMo9V3WotfUlQP4HUXdis4RWAShxekQc5AuPKrDj6rl9uYgiGRCZ4B6RSecNNW3mjITjVwOB
RvHBd2gi4iZIAoqeX8Kl7Mo8mq6mO0LTVKJza8ujwWHtnhLdGv8foW8BgcsuVj6VcK/4zpP5lCex
3CKPZ71873i1nPqgv5rQL8cEyHl2LVptKdi+OJLn+Ph3s6BZpjGaixubzYQwsUI6H2vLAlo7Y9wa
9H5UPACwxruL0lMUz6p1wzxGSUgpmUaZ+qwU94IIH4H9VWpFmjsCb3HRqWkmqfCjENmHZDvgolHt
gT/n4c/C1RAFNfkpEyIyj2zYuyhpFhIWX6WGaczzEhqfuFr3NmEe02skf67p5eQcBi1AcOroBHUx
J9gcpgw83A0Cw25djgm2nJN1RWfZrDBxazcSljogoHXJor2ip5IJM1aYKRZAYCp0V51VH2D2IXFS
Oh5Kd9zHuf6NhVOI5qh6KLWAc0z80oJATXcbSRRWg3xBPetjfZVEATiVbbMPB4qSzy9qz1TKFd1q
lLblh/feJZbV/b5M6/HYD2lfRL1BiKfqKu+C9Pksf04cOPUTV3BKQWsJ6rDtF+HcJ88GELQG5T8l
DYVtairbeaPlvgLh+pyFF8oVMhhp9+2k4QlEyjUGttrpOs1cmNm7GuUvViNXNN2w8Az25MsXWZHD
P4iW3smWzWUVwNU8hYc24urJvv0o+uZgnESQaDDobmi/85N1+Hf/U1UpZ2dpajUIrVN2tRT84xKu
z3SX84CE8VEVDSerub4iCIWBqyBnt/TjE5FhZfKldCiEItKOtYl5J7cZnpP3QaKbCrAkXLEKVBIB
N/9fRvAwq7v0eWAMlrwtUh/z53PSID8KN9LjZRh0ggzyJ9AvzyQDfHR3ree5LhrK9qfRHr36i/YU
JujQof8o1yudslWb/lKLi3NnNnYzvsuE8Dgv99a+UAeAEJtBEiz6qiMbrAxNdRVWeASCH6It7dRR
171CyzYvUr+/+pH2/C52HZN/ZVI8Fga1xNCEZAm+uGdFC0FnZLq7KeWI/tnNybr4Ty/xvDjs4rJJ
JDsibFsQzHN8ao4HD2/IsCxBgb+yjy2uyWsKUoIVodCs6a45f5ejp7g/IKJiuMgx5GO0V72RMwBm
MusrKjuZn+sWlR6gqTPjJv+muQTAPtwhuyo/76ZseTHBjoUu98FSuOQHMG5t0532jFr32DFsaJKx
bMs04h9I79itvVtwp9eqjvTWrJIqh7IyCcj6LUDnY3RxIhOpSjvRb4tH8eh4wWAZpY4uLZ9uq+ol
4eNHPBhtEp6kmy5ZFArTmcKy7LRrv1sVy+wmAB6p8PrLsYo61S4/yM2Sz0KlQkDu7I+rEPBKYqmM
uEmHF5acxyXOkFV9fCxM7+Nmung0TSXjmP9+pK1lgyZasJAppCMQhOBuGlrHMB8/ZpW0nSRq/HKP
8pQvY1bjocbK1Msv3WBDfhp/m7f/e/wW3tOHryVkHKlwhUmV8sfn7KQNQZxHj4D5VUdUqgvg062p
/vsgcYxs0JQvTrc8M2Kiqg8RbARBLnY56Rbr4vmHz8yZerSZnUis3pbLF7fYl+wB87z6CHsaHzYP
eFvaCKNYV1x4yeDa91B3GttD6g/SV4wDX6Ttav24gntYYIg7seEJRDyVHxaAd0jsB6E4z4w64LYv
Jx/txJTa6Ruit5+JcO4UEoF9n1DYG6CIn+ELVV8bP/5uEMbqDbtU7IIGGx8j0y1Z+HhjRHq4KE7U
Nj5c9+ulQU56fc9OtCqkk4UcSMXBTkkVyyn9jeVBm7T0GcVJgLocktFREfm6jGcpzBYqx4zK6D5k
KXhaaHjYPyCLLDm2yevNGT/5JN6ZdbwpWlWpJeqEqBzDXWd/08wJ4RjKd5nEg6U2wAB+8HZUo9dz
QVKt8AweFGgRXmzhcShMqO9zvr/5fLW1timRjg9U2OaQQl2CPMWo26Qhk4+0FHvbiP6AgibF84TS
6ZpS6L0TG0q1eht3ieRYIF4aIh35EUPFM410M/zZ7ZQJZcETqMVYPZHGybWevnJhQD4JWreQxEOM
P4Wb6UVlP+1dmrYmdCbDOoiGZ1oYR8qeW3NyZejq9HNzYwf1i94a0cbMBoVc/JCc2RDfhjbdK4v5
H2ROMiywGY84Sszed1xFzoof710EpwDbP9XLePmjadA1g1FbJ2NUVEfPlwM5POJT2y6HndaLH0w2
3D1XLZ7XCBJV5rTnJ3tzWz3XcmObJ0OSzidF8t+ehDwuIcLcSg0F233lPPHa4TF6OkdC2TpIacWn
xlVbeln8KS+yi2GuG/feeYVEj/h3J3DHPjW4HX2btK8nkBKKC+uiDZQU9XOsWltjhjcd28kfFLtL
czRzjofXB9L30iCaHYNUhEfjcpIxacF7TJGge2J2Puh8pIzjkOQH8+1lc1LYIKnJhocKEJAZpZ8i
4Jzx4SuZ18LI62oQ8syWhZ2Edp1K6XEL/wsvkCB+089aGV0k0l0Pe4+Z///qoufCJsIvV67YIdt6
ASx69xlKVMq3WJNMKbmulvuxKn7Lw5Xh1vnTJjwEX7gG8oGjmq+uN/fWAT4uhdqO+QSb/mEEtHDo
+av2f/yKptkmpoWDpT69dav6B5fC+qWt8An6MJox3w5SxVhkqy4hK26jJF2jqPxrsJJ5A5YtGelk
1NjLFj5bUt/ic0XqGH8jPGWBR/SbWL3VfEn797zjDeObcwZrLgokPIQJlrzVdD3Twiw5HktKmgos
yuMizoRE8bIZvTQ0DE4Ugg2dZbRvzWFijthdF42lwJIzmq9LZp8NQcPfxsbADxTmYkTqGxFDoosV
gBya8l5iM4la4P9sP18NRv53CFcEtcBWA4remdLX8/JVjWHRnwZ2N2hiZ6nAcIHPQDtrc3Bx/Wov
eowBHeHXPcRmZuGRHskWyJUrRPyuQkHmr9cIuWbMa1pPZ1SFzwXOSZjErMe0y6E08+pGXuzMi0ZF
34zkQdkOk1KeFklFBXzR9pqxqDkUGsOSX1546Feyog8K01hafYt90XKs59ZVnp5jn1QsJW3sZEOB
e0Bwtntlzln6iSSi0meWup557yLd6G2WJuSrIQ97MsRMgdrM/JwZnVmp/z4bpszrLy/Hjj8k8gpw
siuYmIGczyGPL2xmZ75anE6FCB3EHI+ecIe3GLD/8Ym6ruunBuIDBe51Rwv0PuGBR8UQzb8DhEjE
imwSaZLj3C8LNoD3dl20DaX9s2ow3zdNnMqtxL67BjEdn+JXJI5XRkYAxgGKVsSwGrl2Yss6fKc0
IHo95HzJtEGLkQpEtZOklr9wVLsUy7KdqcYGpatMBojVHY6Y1b++fIg8LFPzb45jCk9WdAeO72mM
76xP9oZaIZQwvI1Wzxru0zDe5A4Ht7zRAWY3mMDi0HXTxoOaq7r6k7d29QpR6DbUdcfmltIGVTlP
2MmkJATqBaavZ+k6hw7Mwup6jzXuzHJEkfXcGeFEJGIbg+GALejiYFUNpD1dzIDMIwCOuuuhmzLl
CW2wUpCC8AtS8GA+0SaFgVFyBACoXPGfymEf1NpNvDbbxSjcOFikF7GcihGcqqmF0zfqM2ZJ03Ya
1W0i3jW+kC1vIWdRrtHyAxCH6H24ClYiHUFv4nIZDRFVDd4EY4T4VuVrJfMz8dkpw6VPeN5Kh1MF
BwZA41RfgbGlKyLpbZFTOwBe9rYv2QL4KDHR13Ed8z2mFR4Fe55R1POKeAKWRbfM8e1BkKKJJ1Rx
9AgaQVDb8KypSAjQyXToMao7G0HH1t1gO1vfmznl2pK64sxpCkLKoGgEBAgDV1M7mgfAQrr2MYqG
x8KGUxtocbqftxDiWrDklsW2viNJn3BLCXsq6RTcHnGdtvy9bn+e9M5uq3Tlt6/7hCaewDojDGrp
xTb9Mth9R4NjqquoNd2bYYa0zEwC3tc4kFCOpLEdXcC3DdZpIg8D937tA+hq8ZqM2AvB+/2JEGfg
cygTZObY3oyI5WfIk2jMmM7FhYeIDoDYZmM4ilnp09tPdMbO0DTTZSbWhbUdaPF5TQbeXRb8O+fJ
U1tA3UpKhIIThfA+85P7Y2oQClJdqBEC3LTnwQbNNkaAR30AgWyu9ExynjL+WvK2IfqYhMB4WzL/
/BKOEIFWAdF9DU0BrPrkeMyHLks0cS0zcS+PJpn8QSjFa6PhWg4v+rCo0HRhdkMh69cw4lHnL8cj
LVU7Hk9V3i/K8UzE91C0ndYMylZVMbqswTpC/NOMGGW5Oh+1IaTWCQ5/3j2h8JckGNsjNSnz5SIQ
tg+WG+zVp8QACgi6fDbDgnw2iPc47dnCcyxiiK0dnI9xdO5umllFA4CvYezSqhKP95z0PL3TFXty
MAoZ/1yT7ehX5VN19PSzhf4PlFyIXhGdskQfLp09H+YpfHh25ARDN4/bXZIhKKhioyiBfUY7O9xg
ZX9/Uge5LyJJbK9M/luW5kRzs5sJ7Fb7J/nd0cVSUOSEGzzGnHvj6xH2zkd6pdjadhl4fT7Vw78J
HhD0QOADfPggIOfz5NTWCUQBMvx0GRWCGfkDcF46XIGHu8VF0T1vUVK9Fkl/T1fXBrf5JNrcAand
BTu0M1mfQIxjXLoyMdJIK4uRGoA6bu8wAA/4iL2WUW012o05htfuxIiTcSwTfVJ5X85tEyirGwEB
O7R+ZfBJF0xQDK6ix1xUEwz61KqKgRulRJC/8WRJdnJMuGq9ee/1MGlWHXJGLgy1vHfLoPCTsYuC
c0f5nldPoiJHEeXjscqflAx5AQ1vvnj70KsjEgT20gQ2+P8JUj/JHFMjYyG+ogux+UgbOSwGt+F8
7sP9y3xSqK6CnAO9OoxtJjOZgI0ivzgzAXuosBr3AjPDNgfCqQRKVVYo+KPdApQQpW4BCfy4AUqE
VyqACHYaJYb7O2Oj2h1Qk4854jV1a9H+QoUHBYCjVoYDz/CfSk+ZBnfIw16fAYEiKcHFwQVwanoS
fSGM0jlJYhvAKL8xgCLRj9cLvMBp8NAK98l7uQ+79xKcdIQN38dz+gNKu5LQM42xAlESBSZs2RU4
bMXNhA4++b7TYmgS6E0RYRNLNRvAZWjngviZQdNLJrSZgTHzMol+FY/8JF/pWsLZF3u7Y0gUvl1D
h+6LF+suaZ3VqIzbqnmu3pfeSdt6xq/DnTxErqIMkYqGaGc93vHyKJQQTwMeNJKCoyeVyOIaYW0K
7lfS9YvXzsInU4DZ9HKbsRZhmnPyuSsO3A00ieokah75Fiz7uzDRrcoiCoJzPa92L6JeKzr7Ufr0
vKXzRfwpXVJf5CuYe3CAcngxUkxbyxA8Ak948ouquyUEMFEbzxXIl/7brEfXO8jFFyYMX0KvdMXP
Abrg5pQDrA+gaBmmvPE5WGf/AfUyZ2ySrzdmytnM+3HxCHZ2OsanBAESdV7eXCldNC0d2JgIAboW
/t0TrdTm27FFPc1Jnm3ibHEfmRFi0SSMJyjnijVJb83O78VRsg2Zh6WkTFkgMgsC9CC2hTX2Y5cD
d+j4lIMw/D865Csi4FUcIOPtMhcKpGOBN9dXe0kpsc/zq8QxBPtnvtgILGizRAVlzmcMJkY2rRvD
dcyTDmrN+gAcpHaLx8Zp6nQDr48uSHHL3X2oOlh4OYauVz5OXS81+RFQOeegN/JNKV8fPCJrVoTX
E+9RKrUBrx3kt13gAODE0hjS5C0DwS3gOoPhlB0pBClfa+sZ1DfsKN8DJ6IxCNIGLCdqaOoeo6EO
4guOY4p834z4hYq9aIQQ/pa2DY28zApNDoyScFZAembb6kDxK0hA8Jjb54kHZCxQ8DxMkuVf4rno
PXJF4x7C4JyCY8/tDyCCoZm1MY6xMl/Hq7pMarnPVQ0p/dCp0Wr2kR4y+FFP84ojL7oZsh+0u8Kh
EqAe6F4P+Bx0hwUjG1FatrkccpWTAy20E6l8zU2hfKi0iiudlmwnvT5GNWuYhhXtVLJY1va1oV3U
MN2tn6iy8Iw22yUJ5EAUlLicNDnD5wbCA0SvMwtSZfU2SDBIXC5/YDnX608/uWF8Bafz2Wu063QW
28ZCvkedjyuv3pkLmOhpdxw8PfdrNKBCSakRm6iR+kH29+ayhlQSP0JSIt4dyT+Ji68XKgo5nSa+
hCqkfOQ+jkUlT0ewJXPIYI0FCBo2pNHNAeyJXpJWRhQwZJFnioVpO2aWJQygUmr6Uhv0MzgF+OcF
Kf25czBtRggT9WOrxXXaPej0cOZTsFH+cBFdnBrYtope/SP115niiUD2oGzR/vyEiVKKh8klBY/y
2I6qNv/DzzQNhtv5o9neG4HGCZ/PPSVSItJm0YqkxYw+7ynejV1M5xO95aZzuLKrSOel6CccYdsl
ahfu5ODS6VEjWq/xat4spKnK0Hxgwm2soq6MULGWC7pfDwp3IU8pzqZ6pT6mtRSqdZeBwm28Cbsh
0yLglYz9Nrq1ZguORLvOCCLgRzoCWbkwcgG2oPHOxE+OQTTiW/+n4t0K6lm45a6fxMAY82A24fX+
LZNTBk4H27gaFPXyju4Xx0TfhKQdqtEJODJn1zP/riaawjKKuhXxG/+6EojO/jkuOhgUXTFGA/xP
sf+LI+ti+Vp0iDKJ7Z0qzfflnqG2iqYdjDe7wtFvathjHyxJE9rIvh5bpiwR7Dd0rQ3PzS5QsWzM
afNrJ8Uz0LIZP+QhJ+P5InEOBaPY7xwisJuS1ljyCO8nuOpxX8YtRtSP9HYJS0IuiUsx0CJSeKUz
ZfA3gLIrwoBk9N2iblA0XjJIS9mpOlosvSesMjeNgeKeXOtaRMLRcBr8LA4vshSjE/srayKaxJs6
GVwMMqSgFWg1AU0+t4JOQgvq2939ZBhmC6VYvl8RMznPGzrgJXIsDvGhNn6FP2x21aniyOV4w3dZ
XYLgbTtv1oDXCgVW/unZeo0Hw02aiLlzRczib2jkLHpBQ5I5Fkilsyb/d1RMB83L6srceep/MUCT
rCegtzUO45JnNAAmF8Md1p8HEyRtSJ8+Q45SbHHPTH6m2ocJ9WH7Ek+H6t6SaBqzUk4PGbOwiRHF
6m2lv0MUJtTzDPQBm6hQdZe+H96dIiDaKlShUDWFvEOIO31WzTG+WlE8ZH/ZLjlqFuSbK4sfjOwd
cdhXh+MFGnHoyD42LD+gtSxgFAcB7kaDZI6GhznfsXnKYQ9pIVjvysMMY5xCykxYs19wfsMl8+5l
cFJYj8Erac9wk52HxF21HzpGEKWCAPit9zQLs5KSaUBrtrbuIPmUNX9CZr0DIHarVgacEeT70gWp
E1nGF+0+A3bg9dVxdN2LfNVKgK/Pu/0ADuk26f31lkqfmG/UHQHPhg0D+PWk9NZ6C+aJYFaLaLDP
50yTqxUwUNLrzoAVzTf/JD29vlh0SeFlUjIL820vdTmYABZuy9ILZD3Rqr6v87fTmDJD5gq1wcT1
QoH0S7Xsl6Umi8yeH0TukT0wpFdXmThMmipflovP8nTYqJlkvyWlsqZdykL2//yVl0eFg9VZyDRq
I3F8kPEnvSiPxTyJMVT+ySVwAuJzTNIAIJxXMPim4ncZ6TMl+ndvJ9C3eoFe+5dD9VxUy21TD+1z
dejZ1/7DMfohH2k98mX4isaHgIcVfw3EZZxSO9DeitKFKcH1a/xt9qNfcrVUnF6uX4SknZylL44e
Uk5WUc2JS+RuHxKZLJoxoTxrMC3zFJV7aV6RApDOQoP0pM0vY7n9Y7l0Bu1p53/i9hMahPKOt0pp
CrNAKPS3RHV5usy6eC8xDCZHvBaNeIJdXB5KTHpKHoSEh5gj6hnjuDfdusfyqKyG7a7lnmLLf+Do
MqgjVctF6kDujgTfywxYeFj9pE7Qvzo1qBJClTfpy4RJVGqdwdkNDiyz+vUpO+XTLPXS3kLefRTk
9JnzdJpHPxvCV4qZiIytBzSoSeyhksrhhfbTejQ3Wu39kGazz703PBAtBVLGa7ABcBwGRkeZCR01
FF1EB53fy7BJnbQ332qtjFicWPG19Fy40TsKT9JQUSGYBwo+b3b/1jdmHg+koilh1ueteLhVRS2p
EYWr+d0jALaUn72ROjt/iDUMtJ0QY/5a9fpFvBRXdCCMSoHmg2RkPAIQsFMyoMDKut873iDaMsjz
Kxmrj7cE95DfSXZOYgYsgD/2LL+MwJc+40iBRK7MHrzzvMxPYp8UtRdWRw4Dc6mJvjirekgF8OPH
9ZK3DujdtDyZSa6JaR8PZsOaCF0hQUFOZUsHJabdlRZIoTwQ6t5nv2U9ioMWVq38AnaZJoTmXY2d
/4ymL4YCMmq/cThatOe43YJYwy2dz0qU0zDhZ02uxJiJTotUEqGFrJCmBnrNrnDtaK0PLK/3c4vR
gS+RSFrE8gTG0SxeUBg9ZR+nJqvv09q+HLTg16Ab524ZtBeWnDV9DIHexc5N0t1LTwEWNCktHaVa
LqwW4edT8x2L2M1rnUqNffwYz2bzSa9tDjwUnYRGBvWlv1WgEYO8ncpMJo+K20imrDl8GrWdJyXY
hVD58f824q1YEAsk9zdGtx0kVWwAONYxTZYZ9ub5EuAj3UkX2KkE+eo9Ozj3yF/BkdZfprmaYb6F
aUD1eLT/fJlUpczOzmgBxP0VFtcnmz75CNdMygXvBwmWPd3fEFvuClilA6Z1XXGdbMftbLy4cERU
EOzwFaIx5918HlllQgxzvQGpSgbL1Pr7GhTnEI2hosUbbJSXAHPyp0BxOBfTuXxpwUxxjIICVCOK
Eu8JJFg5Y1Cgo9LBAQTDSHGSduQ8Lfe0yFaSNDZv/AcUtO50qLCXX1+ko+nhwzb3rlPEtPmEc+t8
5xnlxIW8LpN2zqBf36QGJjKL9m2fD5t7fmlrqM6dfvL1UtiC4O/2eK0IY8UYaguTY6Y18XIGtWdi
IjoD6gig9lGjXlFukqR04WcwoEhyrCYyUUFC2qUljGhR6pH9jAtGtrVR5CctQMpB4CZgAOhDizAj
3ce1s6oBRZFDuNVbjsORw3Cgj6uNeYU+Qzx7X0qh1Ww0R8oDy873GBjFpos7BCttETVytEclzsGb
Eyjc2QCuUznhLYzWDmQRWyc12YGieh8O7Hf0u3aBy8qq2l33eLNQ5an97NA1OeDhDmh3uHrb81uf
nOtecJehEcD4lN77IZp6hMSCowHpdjbJ+hNsaZyszgXTbaWI6YtqmwR3YrKA7bPtAH1EteXzu2+x
/qJymu/oEMADMz84j2JwZD+2O2Iwpr5cig1QQFTJntIJmURvA1N4UKO2hVhS8l/Cki9E6kBWwVBI
EE+xtUC1mfprpGdnblBvlmobVb9dPZIQTXnIB9K30XBlSaqm7wIfBONcdXxkJy4EyU8eZ+1u99uP
utdqpPfxmK9wMtBP4o6M3iqsr8r4SoyQukPDBxx47F+2kygG4jMwlsPRgm/MX1qnSqVMzAUsUuov
3dWn1GPmmGwZDqDr1G9j8CUIsGWTgca+/3totU5VP/Rj+vTQ0mw7JmftFlgYYij2Vy3RruMtKZ5j
a82SQYuddJXRNEqbCTnuOGcB9JYWri7zhJXo8/7vlnmo/SWYc6819JEfQ4wWddDypSeu1Lh1n7AG
+Dz+k7+DAnUeUMI7P9caF11bjQ4J+QuyzQVlXrlP423CLOEBmk2UvpO3SWqZbJ7Bjb+tbtUiwoxm
xdyFFAm/rYPa/rNL5Cf/zDQwfbKKY0pP8bKbcrdD6AtRyOZcfYAfttGxz7tyjWnXx8N7uJTguMYZ
x1iaPdJ0TuY61C7Mpyw6gzz7JP0Au07z02FsUUfvENR/PQCPUOkv7K9c2RAL+cO8N2gNk/6ioONX
lzoCY3RcAorafuMDRm/cmyZtgpS18kDtZE6korB8d2C0Cn1n4SrECpMmUvUE98tW+CooBKuUel0j
W1TTltnwgRv2KvK04ZqWdZoo+6ok7u0qlyJwl3dBLWsEqAZFnkT8sVRDBTAQ4Gn9QmeMNNqxDLl5
5y0m9uaj/zTo+/y/hYLA2f3UW/ttzf8NBNIu/OnmcjnIL/nPrs3Fw5KAWmD8GecrCz4C1ff9lQbe
PyfU5jZZhVKOaacJQ3lxNGLgwZ7Dw6990bi51bH4o1+tqouXQO6QA1sGW3H7Kz894xr8PTBHKog2
EQACwQYrXFjuHrxOQM3NAikeRtQ+FlO9YDS7S9WVdUbZ85g/GQIbtg1tfs6X2q3v53Hwfy9IUlCa
ZgT+V0XGcbTjp75z+JtW+Vc9ENm2ztdPz9/gNUGpV/A6mjPT6Kj3/5NuCJnCHFCHxRQbN0NmSwlI
TqXLjAiWGSBzLCDlr93BbBctomrSM5gs1O2mw9lctSVa5AT6HhYDNs9BbiJV9DDUxZ8D139Ga6G4
btMweOe4bYJL3JZvMosZ+hGPyo5k9sNacLIkHPH81KITqgqD+lRP2ts+RD2A9NDIoHQWou61mjzw
WF30OZTB5lyX33kWolw2vbCG9j+K1UlHf4K3/7IHUEWlXnewptwByYo0/+lKTEXQEmAFBJmCzJJD
iVA4II6U2P2QHgZsgnGA98YC9t5WmA5Qvv7UlncQUEnDvpWyZB2jStmYIR92m0wiyrZSw0f4nE+J
47S06YccYQVcQtE2phOA7QKqajrxWJSIfYmMKEVp1gmbWrvfSMJLMKBs+2yziCqp3buC2YtwVB9o
NGtMr6nLjau9qthBxX+H5YwrhVEAwrD+/tf6gRHPn1+wf3K8R8UtaqZ1ROukI71SVwDstmUxluHW
cDHb9iHvDL4rf4tePzbJqMMeinYI+Q3H0VhQfN6j6YAVfDq1Ktdaw8sYz4Zs0Sfxr1c239EuQBYC
kNEv25LsGK8WtupbRzvdmaCGn45l9/IOPSukMuFq3ou+e7Fd1i8RbRtYt+woar3wvqltin+CkW39
cnYYPG7bpS1bkR+BZm/jXXkAGtR8/sMqeb3L498Qm0844Gxysu/XNUBvG495BwgJDpuVQd5QmZcr
CNnCv3Pu5rWE4gvZjn7ZUXVHXLEGEd3bEbf7FEL4BYucLfgyhKDRA86HHzMrC1DQpfmLpwg0g5gV
SZhWuyS70L/0aBsAL4btTaIYOTpFpUF+Q1DhDQ2HUcGIo6NGivwFOIZbhmbaQsjDuXbgwsq6oRMz
YU2vfu6+rXXeX3KjjGHhn8WmlPza4Z4G7vFl+aQYHtm4ZlUObRfXTgZlmG8CtQMXmmeXwhHQ6gOP
q2B3ZWAVPp5vCst7TK2YW+yLNuV8BrCnsGjI3MnnGMMhXnMYyc8jy4llzDFwDma/HXu3cw32dE/u
xOyRUZ2fekm3/1moRxtaxgnLaf3J5DeeUYlytOHmYt69AgmezFGhYKgTl5DI3T6UXGPeHRexH1rt
fRPEjolQExo+Kjy2QwHyOTDJcViP5M7EDI0032KGstDh1l3Zd0hLbIcEPM1TQJydTaDuQxZz/Bb4
WPWfXrgIrhXGCdKFWxLCRzxJWKFc2XOke5evK6l9mUP6lMXm4eIQMGlc+6dugVqGgt2WKMxZtCIf
a7elKeEccJQPktfTm0Qtd/V9eeHFTjBN2q+jMBFnQcXDdJMYch3SOzaz7yVRGv8UHkPryNuy7IWu
o6bDYrTLfAsebDFyA3OMykqkVNWch6htj72HRBV+QlFONefGBpTsHnqORvLylFhARhK36yMYbhNN
SF0+JFKTaOfJOcicDwoKh4dbQHnWSrFSJu702xHnHEt6YEUuuJRBM5iFrjE7IuOeF9RxsxXh4HfH
7jn5+dKv1BCyLajLRx8aw5hQFLVyAfJKyfR94AKaWIcBZaX/6RQpWLVXwHmnUwUvnkgsrYdQ9BlG
DZXPw441mR+bFlgRPNmBibU9w8QutEIzs07NS+4zv1PYqeRZa7HLxefUh0rimjNo/EueUy1T5XOp
d5edINQh8o5ZuotJPikfxv0MBjaOTYvKT4lVcqwUlT4wYKBapEq86Uln3rovWqGFjdgWZ8j3XmkT
/8jFkaTAVniMIYOXjFV8zAXQgBxMnNzMph0WDIEiJsNyUCzzlsesZNj1CYGPtWTYwNhjFBp7xljC
ZyhNPJKjGycj+naEH69OHZBAJGYQ2beXwd9GNaS8xFAYaF1osxAFVNc7WGxzwX3lXUA2C8uA+6r0
rKt09OUAiAT0W2aTyRnanxSR+VjO60EYXwL0iHMg7koEkrYeptmMkZQBOdCmQEyfkJopv9TuD0lD
eMIoUA6FuYrjX/wOR4SXnbPH3YrOolbeC1HhBQQUnfiL8wRZdYiM/2Gc+tqHu8hoOVzb/wh/7lsI
eMoovCeYXytx6oO7Qor0m7veg4HPJManzJ66sku6SOWwPjOW1Qd0gVum7SmEhbd2Q0P63H6gYG3n
7OJe2QzuO/c1YbaiPT41NXpjoiUu5hw7Nq/aRSKMheQfNd8rAe1+M+lJvc5g38qmjvXMfuI1bMNh
pB7MC37ltMWlDo/wTACFQQ8/fvO32l9y2XRl90UUePmGWFuaBoKqg6ysVL7PYD0pPk6Hsr/eNMys
Gcl3OWV47bQiJ1wRgPcfgYjXnUm9DogtqPnOrwnaU3seUURRd5FrvBtfUj+D0/5jd1K+ecy3AV7k
4HjoiimURtSKASHj19M034+HHkz18fFQZNY3uDmOtCE4G76merhOuEueXRQOaUSnX595BzJ9OfK+
lIbWNMqBgPG67gL5KkyBRdteKgPdNOBVgTwC8djAqoPhJBbL2Y7yj2/iZ4yI5GHRvvhEM6B8BFjn
xJBJpXyzsEyWx3oxa4xsb8KYFn7ajXxSuoIl8t3mMyxRDcQ2UhvI3eKetSm4Pp2ZVV7LFQA1SH+e
/TmhYmAY5EFfno+ahvrBrN/zRCQSdTF+Zg6kES0JF8MSrV7/5t+3y68YIcq3jsvCvT+TCtUovG8Y
SWs2BsB8UP47nWxKJy8PxbLB140Stfcg+g8yQiHwlDVL02uzVJ5rcEulUpLPMVQRaUSUu/Rpx1UZ
ku0VjJs6Q1IWCPcOt2ccBcYaY3ko0c3ffUYxXkgl4FMWUdr/kW557JgetHPEsB0KQj7mnxsmsdVM
s488WRWBQOuVofZVPLwe7/pyCEIODkLNGpJDXhh6Qi1j0pK3qX24JTEl3JYaJgFTuarjK0aRwAFt
rrR1ZznL3KC6Wpvwu1VtUZOPKTjzjHW/D90jDPFNDUg4y4GtsNCH7pkKtXytEk6e64QI6vBvfUWO
IgnEenigsuvLxlpp2np+6m72YL1L72CsUU1ZxlvfqR/HTQhsAFbIQ7o9WeG/9AfYxmmvDS7/9MTY
snf034A1Vz/BpASr/4V2hqThuZtwwoBBEgkFNtPpK2POmR9gKgibPsiPK+EzCYVR/ge/8G1usSRK
/ErZ/stXh/8FsYFvkgyOBu7ygzmCapD96o9JkTjWEubgLyfu4qHs5ICHTSWvVQQi3TsTb1WCEZfa
N87K3+DvpWqtHvumRCerPwmI8zw4g3y6H60kNLsXX0CmlFVHa/SwxHTsz5wBx74hdH/jbDHh2Q/k
UI6QobVI4Un1y4JWPpfzV7Up3TTm9OOTiLursxZdxCGIFYjsoe8WVBD7i8WJggdmXuM+Pu+GWtfd
CWtzo4s/Fb5aGlueiM+G0cO84H9Yht2pbiSAq77YSfntgClPItYC6CyCC9w8F+whKCgWnwe7S0a9
YVAzEJ1v4IgZ6V4FmaTjSo7DcvuslwAkfe+MvLOCcIvZjHfVlAIxymHoQHvJ6QRd6mv8JsJILKrY
2Ea/DJPm8ZoJmZc4PGTsd0FXRwnNkM23fGUrVq7T8x4FZPxyH2O4nHZ7J8HHZMfE/p/8GH6KAoip
A0aVDti5rD9Mj17bMOIJ25SK4btENu0XHnj8QNGKihvYV0BreO5YM5p+/89A3CUKS4WM3OLzBKbX
Y3dNZ58eGpC7E07Rvg/YYHKJhNcYG6o9LV8Q9UDXI/J7jy9PMomnT25am6r5H8yrtuJFsh0KYxy5
RRJsFtywKPW3AdGshbtXPadYxeDhojsmyt3K5/Z+JDsAYfwtWLuJqmvdwvM62hTqs1WxAh4iSSv5
j1Xjf86PaXoqeVVt5cxKvvYp1VYQw0S2DdOCMNeiPQWn2qcisOP8/wvEkroZrT//tosmP4hkQL7G
G340F5Xn/Ia4iZBN4MF8PWjcC0cuBr8HAfhD3QYLRjfIWLo0nz+2m4XG0bamUYE44AKj9zqP5mV+
JNDOHyaFSPO67439sQFWC/BulxpVJfXlrpJG6VFYAmzP6G43PiyUTRKVFjTkV++BudSH5N4Lj/x2
Cg6TVsCBmdbJ5fdTVboHa870VdhDr3Pe1iiV9ALmWgkUrvWwq9R2HrFyJ23eACBraQXw6vljoZxM
4WZ7V2eGOrh9xR2NtauMM6qaQ26VqJj19tOCRhuMNtXdxssuctrHE/kDXtr6AwCMIQeKanWkuNqw
IrOOiF0MuAGUaTOVHtrVpzhfKEge/Bnwi1A/FJqbrhRoYrUoU0FhQsMalH7QYYdFMNbtQWFBzPdR
y4kiL1fCjaLT4pLsEilBHRMT9GWmpMZFiTqZdoww+QR3VecTtPAI0S8Nz/++6eX5JMfZmSA6WWKw
WI0Jogvmv5xh4LMGaLB8D/W7daLinHBCQqqpWBwn5qQwKdj6EHzXV3Led8oZtBkXwdiy1C9ZAzZF
mJtpGteS8bua/pvIUXRhsFQh21mZRp8nanAEkOKU092xPgRPOJfzz5AagRu5RZRkBf3XWTlYWT36
/J0cVYRAvuzvjS2ZuCHDJK4Xp3z2EiW0c6kG5r+pach8hbg32m6WMuC3HNGch0HeAXKjYOjMgx8S
K2PU0ukIoYq8OId2c/I5KgBd+SCKAU+n04JMe1Hwcd6Y5DXrBtqFeNDVJnbkicvxRf6ZaVhNFwB8
B+Da7nwMzPYYnxYy/fvR1qmtKVPpJkDuh0R3juNK7J+EysPtuNt32crqPbpi2FPOzcSg35PTC99T
iB2U9KbWvDpeLZJ5xgf7eAEuGpGQ1FSTGxAvdo2zMccFQrBR9Of9ODSstszHHbudM/xZyCRQcEAc
I6wIvE9IdCqfXxnhQ2PE18hm8koU6hV+eiigqb8tqGm1c/FyOuAp270oB/Nz9+PvSciheQLdVp7U
dn8xKjsbj0AR9PRAuncOt5vVMcYbyrZdEXkFffACTMXRlpYvfVtoIW5gjFXzg8v74X4tHP27xzi1
43DVrNTwAx01Nvtje71nCUmt1L56eo01FUSR7tUS2jdwGty6VbvZNPbgopXZXaV+AHfEgQtDO6Jv
7FoVwRGH+Dx8p+4OLNpvMR5IcI5gwpJkzfyY2Ia7f++B+dpysnz3Tqwc7OAF6so9grr693KxFvuP
nslUcWn9CTkYgLYydG7j2CuFLEnG7Vz11cp5FvlUi9vGURFNuD8OlYdj9q7E6dlhObOxQcIfZWMA
SKI2sd1/J1KY5c3gGmmki1CvT6ER4Md7bbUbTsgyGlFbfExMCi2rHQiKduhtKYrSCfMLKwXkeZXA
yZx5H2xzRoRirA4B33fyBt0LHioUrWHh3BnxsamFszBgIT7P5xnvcZGLonLkHdaPjUK23jvW0DIz
HlJwly/pmt2SSqXoyGhw3ohWExsWFQ+V7Z2tBqDTfqAakVyKKwe4PXppVq4OvW6r2Hst5wRDppf5
DAC5ebgciV2tvXqHvWp/nu3hHA+XSrcftmior+CrBb4K6/PnBZGt0Fv6j6CrnOzKKxf7XOMNcoFI
FDe1JuvhCMUs0hCqQDWlsY0O1Xrt6rNjyCgLPYgXLXzCT84woc1Jjl54pZPuwnKc9zhhNqwubN/B
4MBHKcXpMiXI9E+JP5brWMCZQ5IoQNk/zrC27uLpRDwHFiSN+q8kzTxyO6caWNOzWda+hOQffCjv
uONoyeArFb5cE64tAAjf860OygUr9UXTy052o/MKe43nFbkFaB+aa2VNLy79vQrGym6zyoO0hH9L
xscLlKjmcvnRWOH68lnwhohZDQeAbe8G0garjOpcoHrD2UsVgAsRtosA4umh1xXj+aPbRL7JZ2c4
ZTxH/LomUvxPB/69lpM476pSwzoi1BBNzVhHx7KLsmZRp5SG/esq+uGCqT2ICT4SZ0gds795Ldex
BPa0YqQzqHn6gBNxzn6TwnCe2JzWWozQYhNrrEr57zubESTTBLOGzm7CyLUPIcZQXQL9+BLIK6WM
veVSWIyT5aOJx3ntlcDjcj645lp40UxYNohu4OsRyvGmVQq8Xrx9vu6rj6HhDpHoRkCsu3ehYGoQ
9NBiz/aDIIy/yJOu//N38RsK7rmKK8TBb6zMN2U+t7yVpG6NLrXCNUnjfArQFa5D7tbnqgXitFuZ
kanLfJq2vSunqfDxVMnMgWZf+6aVIon027Zxu4LUmMgElxvWT768yhJ1inp+cwU9O/vhMWWOVUKA
NqaPNAsa293KyZ/Ps8/32Kc07JLDPX4IL5GR5MTg5W2vV5vn9HhVbRlnkmCESk3iWTogvgMQGotM
Et0FGtNf2o5zNM6EEvzBjAr01gTMM1DGMxFd43qX+ivTely9atYKxB+A6eFHlP/1s9jGelRROtMk
0wnMtzjmclZ0gz5BxlgPRovGUaljZWxjMM/X9wdrlsPuQQ/7zyyevGwbHCgAejVBPTStM1h9YQK8
cGj6he16ZKJ/+ABqgT29RMxP9mg2GJv+H0fMXZJi315xhijoANUBWaepzGPGQNuuUiJ3rEbRnS57
Etb/zEzidpzi9KzF7QI1hjWQjHC+OWHRayeEJurOJXn5hd4NIBd3BpMxt9As1hQ1lZCvF/aXfanM
oeR2my+R2N9YJ8ij8C4wgLHjxy1E/scABhytOPKSc6oz5kNR1CVUccPTv9Gh8DiujjdtLpVxq5Zf
HiGemcIIRdJWGOy2vTPtcrXz4QolED9PrsZM2amQVk3ufXMbsZiC2QcP01lny71iX6yUDwTZ1jKw
Kve97qNBxBzef4X0QQPalzn0CJHuTdqRAd31EkFqCEkcp2eDNVArCaFCG3aivilZDWN5UCP8rfGD
N2KwrPGFsOmKqwBUen9qUHwXur2bvtmaFBOw2oGkdyzgisyT0l8YVu5xLE4MCFk+grbfbqeziSit
Cg04nhPqj5JxPy42ULeqq4gdyXj59/q7NOA3PMDkbr4Ax/sysxqmHAfQM21eTjqITGs7Jk1RFUem
coqaaYHYlunjmVjqlWIoGUV052nxD1uDr3B5+XK+LpNbTbC+Xh/AfaczMQfW/lNDQkJarT2j+CkZ
BZNEMTA4d/iqbnU2ldQQN0N9YwYw/xslGrjABwpwb/SnuT6NWw9PjjpExLESceq6MLokqBTDMW9d
3xSVpuJsv3riu+YT1WKyvemapffSJrDUW2N39Fu8EZW/vT73PeidaDJ4+4Ls2+EbhvoDYxmUSQBo
8MsJJ+CF+ox6ASWNrl5DEPWAiZN1fJZKQCsk2JfjoNU1IwlHCw+kCZhBCv2OguRIbeFbXjizVevp
w1TXkaBvrDpWsw/Wn5e1NEg578rGcZeiEhHSi5WJtbNMK7q3MP+/Amf6F1QZBpBsN7zTXwkmXQIf
izTmDMfUkUa+kVAmigSptvnfSahZCJNYX7B5JJaYvUjwato3nzBOAYc2+BsFTQh0tzVluxk5MiwN
Cfin9UieAcL4EML7KcjeAoPLJfw2pHGF9ffCQEyDyw4VVttY09Nv6Umqg0zdt97jt2GtTTVV7Kzr
ZMmLgIECDVec873bW6rvmijUpNlyE8g5qP4oq0l821q+fc24tcgS/TtN/CI+oi9z9S6rj1AJIHB9
x1l5//dhv1KfhuRtR4uYzO0ewomrHjzu1iFo8Egj5MdQ2jQguDxa1I1huYnReIXxC7DvenS0Pmhv
is8bbgcqPuTm6empGm9OAaypARzRbVmweQ9T+khtBVCFW665XXjb/oAedt7dILH2aOiXHw2X0Wx0
9ndYmrQKbYrdgdu7FvgzhHSymjWtq7LaPHOJmLH8H4/b7NgvByQXSXdWtZbIS3NaFDwVIPdKeQY4
qRJhnrBxfaSac/QxKrcCe316fwRG/vDjHmROHgpHJe4yc2P5YEl9H+tYvaZek1JWw3u1Nj8poAmX
2jh8bg+KgayjYvm7iNyWBVkfYjGmWfHEbeLJY8JDVZ7FgjqrV/5X18TGD+6n0DAZULZ5C3KSG71K
jsI4X9Wl1ao+XKPEsbnwslKrbPVi3s8BODEKdT4hzbp79CcwyP0+lOEjcZKgUYi1G1kAe5Wmt9jo
Xvjk0C+K6XbG6+R6ZYSIlfKTzRcy2/BXvhpyp9dhFu1OvIJpcyGWKjZCPvoo0l6r76XU5iGF4D5o
kO3mj3KsTwWoArX7qroIX8erfLTl7Wa7jCmhd0ig/jAMwodPGY2sIPBhXVxi0dxPwRqp3X7Pgppm
oFPPbUkHlM/Uk0dphBLQdc+xuoCOkq7ONe3r03hbTXDWi6OSVwgxRc/8SQ1EtYjBMB0JaNivV3T3
00zarO+Am09feS486BPu0Q0ql0UQVAx4a0Xydij2aYA1eBZNAo3PmYxr1jZsUvm7Us0dA7kl2won
eeeBObd0QWS7Dak0Qlmzmo2B2iFHD+bz/nPSqTgJ6C5oEmomJ/LNJJFcwFYwZJb1UtVkgw6WTXmL
CqBVwU/A9JsBKq9kdWDzhxaKLRQqyKSD7AWXCqL3luY0W7kBZWo/aLV0zuSYAfg2rrorh0qz9qqh
m1RAnmPm1V04IdU7p8lBWbHukEMpEADjzZUEe+G4XbyYJ7DuBDvH0S8B6JK2Trd5GypJEsdy+z5O
WCW73IxP10X1iLfmvRc29+HB00+rGHFha0unI1TgEwjZ7o2NtBZQ5jo6MtpWw4gWTtKPS3R6iBis
inx7Z6Mv9nZMTZUXeUjirRPLcrDKqIG9c3SCjUbzEflVGrTol4CeP9OtCjH5NILn3D6xy84Zpvys
njmAjJX6A25aSw/W6YPkGyKr32aRbXjY6n5p56RlAHY8A6VI810WmdM4NlCxHWDwso0RzMj1UipN
OZnrGAK2v7rOPBGS9Gjig39MW5hNpGA/yyVKHRZkX3rqTn6IMp7YfLZSJDa2YsvaqHk0gLDkGK6o
UlkOqdTSJiklrrt7BJnxvwJhAiama0iAllYR78Z123EIWrMnIuZTy8s3uQOqW9EWoZ4eA8Uru17K
aL6+MBoadZdMgDaGSB8YwHw+Bs+jNyxZG0tOP5kGLnf6V6w0l7EBOSarcYbAf1apAdu3F8yrbxh2
rK6+n9JNFzuQPI21X/WroMXIxO4siBvz4D0zrSz59TBSq4G3cXiRueX3pWx0YGU0qpwgWvcErE7k
x4ZSv5Id+amfpi8mDl14JetvSf9h0pISaiVVefJlNMQzrNXoC1YZNq4EphMmWK7OocEpBENG9eFA
hpjccw/90Vd0jWqRP4psbcUscFizCIklXInrw3LBDU/V+Q8bmLoXbMEpzNtlIg9q0EJkqg67qExC
91juudAARpOe9aN3aeEMyt2tp1FBTEbkURkYyNlIhZhQyloTcbx7stuaDzy22wcjgg9ET/2iokZf
/TglfU/g2IoLFldZLBUBJWH0Ant7tVBDZrPmx7y56YkQJJZ2sL4sM79nLPdW5g9IGt1o5mkGFxUs
feX55KQyziCG1Ghol6pYBNY58E7AVBaAIkCGzqJZ7KxKkohwI+DsyvxWqNgRi/mLbOtvAHOfbsl+
sPumpcsfckAjClHyP20ES4LVsc5bNuEYckslIb4NMwp7Wm5nKgVyPSjL2URE9DCgys/92o6xAeu0
rmLWWPv71e+1VhRvAVhwz4G7E4Fi3Ohend/b1ZP6CjI1NRYdkwf2zLzKaVA4Z60HUlvbMoex/rQy
h0qVXukmvVliErL0WJXkTMRrDjxEb/NbzM03jv4pBB9ER24c3VDIIqeAbO1kKp14FRuEUY/Y/EX5
hNdufBysmdJHs8FWrXkqoZuhI8WQ+M5JCCcvoYt7jWW9O3WEwlEKPaxWXWTv5hMupYu9s0vwwFOb
uzHv6VZRGmePUKDzk4TMDp+aZDXi8H0yqOf4/5pfEpnXgC0YRBz/xE9A3Nlmg8QcJcr7NPW8FDyp
SSSUexMp9mfqNrdHK90skbb9/22UEbWF3h5Q5XbZVjYsOURxBILRUXRb63wXwN+NIMqWCb0DeDCX
y/6UQJ6c74op/aEgQlz0bXOX7OSn9gqSGBMXTqCLdgbGUxX+FvalcWeg2FFzevjv4ZbsKdpPpuq+
ZlQorVxti3t0mfx4h00S4ya9pxKISeVSiSkOJunoB8QSeRlHYI8WspNbnLRpPdfqWUOuMDu3I/g4
t1mAdlpp4aReovo5WIiGwhgCFl7YiGLdyHqMWiUCFtN/YWVwMlcEVKZEfvBxEJKrCr+NhJ7ZV3/s
IqDnW+0g/iRr6CGTsRMGKiVaenTG/CUlZx9R1Qe2By7Y7dGJfdGEC5IRtxzWOPgue5cD3jG+BIcX
tyPkQBgIchvWVYwgimQGduPRpk0wAWP8cnp5Emy/H0VFmxNk/kbkiP1vnRSFMXKvat/zDcd9rvZB
5skF3uv0uFzJ+GarDlQ1UuZNPN24OD1Zk1RV7k3VlP/r1fuVASNAeD4GQVHhqBiJl+vUyYCmAiAb
deEaIMVITkSdCQCBkxCfF7yqQ4A/huMboNhXfki2fDSPXDeaojFTANZcx2cMBoBbt+ittb5bX+rg
tEHymVh2TyXgYt1K3tSkSiS/6hvts/3lBsHPrjWz7XX5Yw8ILJzgS5BsQlB2mIox9dqs/FgRasQd
UZx06fAczfN3aeVptcH9hKqehF3Y4BesFf1D//VTxVTx5eMtpnAKwvNd4PUOa4wluh7gG9kMLjAI
2R6Pu9ceNXPQ1zib2wm1MkPyZnuvsEoC2p0+l6oGUimWFJmyd/79wY0cijrbs1GAo1ZnoU9V2kdT
lNvxLM9efMRQ1bEmK/p667s3AOonFCyIQ6tB8szVBBkbgYUli4+YH1wMPgkxl0cuXvqPuh6yPBra
WeqH8brPjm/j2zuMD5B82ytLWYP/GRuWw8T34cM8OzUQfRsQdOFyeyNNTJHyDPQba6IuhX2WQdF6
6xuW9+msknR2WALptAGMfZ8ek5oA8gRM1kpXZ1xyX3ug+Rb6oNgSVkmYsmaTlltCHSMdM0sQs3GE
nGT4Mjwrop4L+wcpdRUTzhLmdYqqmN9X6jnIQBM8PraK0uFHg1BbqNXk4hzZlqfRSGttTOKJ8aj1
6z2NmwXhGtx8Ue9dvYg39GaZO+rTzfnYUCCcDcOMVMHRWRktFkc2yTteybW2eXI7jI+KZFaDnT8z
OSKxPHKkJhg7i1gn2HdMG5JxxLxAr/jZnn/ddsNAWE2XcfOWR2V6RK5+PABtML3J2OIb7zqrRrOT
7IT+QQyFIun7YJXDYrjCwgUcZk1osuMaCJCjIH7C4jaXzuxPXNbN6381EO6d2+Cl6k8750aY9nvY
kks0TY05ywZ3W2S0Auou+iWhxiWfioam0bc+H0Hy/F3aio0CtjOb6E7XJHYo7ijC6w5HGanWqa/W
jOK1WpXXqFh6i3wEYjjoVq8zZxXFW1ZoE++XRaUh+3yb/rpa/xYiIAgbzHP5tQziE40HDlenyrww
yrO2PesSVZqy2zwD4xxLjIsduf3taTYB0jLDOCs7K1qcEppstmfbE45vhwZpm1Mg77LxwmdvK2rg
0gmEez6rZ1HuF44l+B+Vj1BM5Aak8oMyClldzj1j9shCHyFPRtrg0ZihCjSfg4NprXYvjpKKvikL
sr0ZWqsDFTiq4LFmo1GCKZU8PKSynMYen9Pt2vCObjqfDntM0sFm0QAPvobM+8tBbsYIQZpq10Up
xE8+9kM9/FWBgBqCml56ZOryHUaX5pz/aAsjW16AWOhPq4oU8tJOg/b6AewR+pQXySXHTrkwyknc
kl2Na36I6UUXY0vXzV5UQCgzbMk89VCh3aZJtsZ8H6pZjj3Rh2IeQL+QdcO2SlKu2snzVPHXOs96
RpHOUHwVNq0truXGASLCrVMfOZEjXqPX2QabEBkSLb2dUpXA4M0baxRMkxtoEsMPu3RRDhwp0Pxt
OpZfkl5wNhsIq33jwC312KJwwsyCnxn4Y4ZfjWD8qJhWcfymnncqowBhPIxieMSAabTrd2/sd1fh
FLkGwz4SieHhlNStLiernXo/jUUmxtiIhu8ivaWngZS/cuF3wL1ikuCWE4YFTX8R8tFRPZdoz9tL
AGddp+uyHh+IIpBqnuUT90+0a8tNx+j5/SYH38pAXug3mo5zkU0gfgyNC18PMPUfWrXeSYeZiNSG
LqIK2uTa3a28jzpvGW4OYyzHP3e5rxLfuCL7gMBc4uJwmZUmYN9rfAbthYLh+jHXwA1oyS9pA0eC
1EbXwwMBBjyjFGvdAOqWEH4wGIPi+iS8Y6//txlSwQIHCrP5FxH+X4C1Gk4Y6bPzU+Z7HTyR5B3+
JDkTvRa6ORXJzfwoR4LT6WVczZ3laFraN9woeF4nZMjkdF1x1h7+YaKo6v71MvChYYHyNWyw58H2
i86b57mu5Mpm7myMxe2rHW+tuMfH1xS05FD8rsqtIOS27svCw9QuzK5gc9HxPLWQFHocg51smNig
ogyKsDBmBE6/cnF4sj5GXV2PFp/1jlY92hJH/hW9WHUr8W4hwaiOGuVfQcH7zAVF6JhOuqC3StvR
Ja4xlhTKt0YMdXR6TXK1ipKgE6I8kadpgbFZw6q78faypyDZpUu7J7vSMJIBgC3+r66X6iVH/sp8
RVWajqbHqsCC9qw+SZ0wtVTIloI5z2OR7VwTWz4b37jHZKbsg2cKTGe6jJABMfkIDOp/4xvdfC2u
mUtOc7lyDkHqsj2lsco26ZwPzEZEANAyBeCSi60pV9i5O/e8XoTDYQIk3+jxwNKRyhxX42jYffop
L+OIIFA+P9hEUWYJY0CeObEVp4mLk1DrMA3kZITUSuTOKn32I66Y2LY6YnaDN/oOJ7o2GZQUZAyu
j3Bwv/mdXrmzMdBFZdnj6w8hm3z2OLGDJm4xM7Lm46h1ioB0GFxYC2QxNy/lWNWwW8JSU3msGVzl
K4XRv31q3/HKefi+KbinoeQdsBhptdVGoUvyXEP9Iv5uwy2dvtjxBHwfrRTqBV2FfMzdWpEa1B54
3XjwJmC9HDdvI8Lwf3nm3Wy1Evp/QYrHs0e8+/E22qs1UDFzjglwSY2BvHR29kG2MsSfH1kMzCOQ
pH4H/x8KAqw/0DT0Mp6I35CwHB00VNQuL81bZGqRKaQ3lA6pX5wGAqZJWtozdVcsNJgfnmprKjCs
uYIlBaOR0982Sw5BqcexaTYo1OoogD/x2MWb6n8zs7BcYXASjkXGmxu0STpTPJXX8OevkYfGbUH4
XHICBbNrF6BFSqdqUeQradCN4Ul84wnnXtv6cKc/Nj8bMhNkHDd2qNCwo6MQbZINflDM/N7o1cTk
qqbc/k6We0BXnwmBwG1BxFkymYo/O9LykHM1Df7OyaQe+O/1yNyZbl8gY6xQRJa/8eQsFmaQ1QaZ
Jl3xL9FvIkglc0sYofkeEM26e8aCCNOsD2rkJlJKFC1TuoKUxK/Vj+E/8JWiE4/WO4k3xXt/VXGg
TEFUi36dpcsZAYI479sHtAdpirWAlWJ1UqETV585m8zQdul0aFOCDrqhOn40d1yC81DhmrzcVCxU
5lrQs1Fh4ZgHc70TkCEuUTZky6t9UdULUeewcryylVYqNiKYjMwVaFaT9I55C8MvPkQh5gKv8JPd
8BQ3sVYJd8/Moz0a18TE3fFSSurAynaj6zD9Y9Ylf8YYO2Oq3k+dAiLKl5l4E8U+psO3JkM7e0kO
2Br19KD28Li8zdzhvOZD9zsqheojQB2z65aXND+pbKfOTgxjqgF29lASc2Z7HQpVV22dmpVKBGyK
0z+uBHRNRKz6JD4ImGdTIqakyO0Ze8076TGs9ewMmujTGZegP4vkwDQSdYvOew43F4bH2VWG+h4X
gGPoH4owMKWKdREWdSOUIsBNO7AjuLAIAE2ETerxBalSBCIttX9Uzu27z6NFffry/B6GqBCgbk6f
WjF++2+4GcxvnQkkvmTG7lrW5qTBIDc7ZB81jdEVhyGxflQxQOApxA3dv9G/3m5Hez2aei25ovQu
oS9qW8wWkqsdSIx7dJ3vfhC+eyfbGJKHxqjCHYwfbY39WyaqfcFGP90ezFc9XeDWlGE3xnzM3Yrf
JL8I6cmrxZ+PqvX86Yd2AZZJc88X0qc0suQOqrNfO1giPuo3Q7f9WmDydZ0ucUGR0NCZ43BVXBha
GLLhYyz1bJC/FodXzNHhz2zO3VTiwSW1WjFwUMMR0Y0QIoVnGfrE9bOfG7JVPYhZeOGxUMqwEhkf
kwE53shvMtCnZoogng0d7n2YBfOg0QNwjSMaPuqsPj7QshXJTHXmlmfL7U/2CgotdCgbtZDk32W9
t39kJB7muMIFlyW7TARiIri8TpQtCM95ZMpYvbo4kr1nwFKzoe4VFUFJ+MfiKqOw4lhWWmM6o6OK
eiUeTu31I7MA5FndGWr6SKLZsvXfqCPu4y/mJTYJXfcR6/e9LbNHuyL/o3a4NVgVzyi6JybKTkp1
t/+lD0WJatQlF16d7EH2ftwYv8+RXpHRxmzS6pBxLwR3uWraEIWmfRlk1U6dKOWiE7+de6eUT72g
V6fgzse8skSR0x0ZT/2aMPou2RB/JCJiiy9iFDeNnpIje1PE08HnmmaKQd7KymgTh7yq26QAeBuK
k6tvS9Rz2rceOO8/Jnm1PiZRafMKm2Cw/jZw5OIL23w9vv/4iut3CZEQhpmQh/uPrI+qAKK3BgBt
ahrxSeLRMExTkJl8Su1FaqI8rHtWQ3DrlrojkWTD/1mTqQbj5z8OogedFmP1oTJBCjlbOQaiWG4G
Pf+N37R3k3FvFHj4eNIRzgaG6Ig9TyygDAM3aHfay5Z0NBZfluqom1KckvPChmk6aTdKDbDDiT7g
6OlJyqEU2M73AAGf1F4RcqfkOicJF0UD7MjbzZ2cyP4q6rQa8Ttlkyi9jFimepVlt5UBrDEk3KOb
N1b4cWFw22iprnSE4OLiSORI0aEDuPnvlPOTeLGBIUCNnrqS/by4BoWhofydqi6SLwWc5Ub2CDVD
9HPUHPJzlcv4i9zeqxCur4NWEfpmOe7E9Qmygj3cTgIAf5Yn0MhdzzgsS0urnRnK1P4svmsXgZ84
UTy5ThdzFYyP5aRtyogIsoCnIuGEB8MHOkRiuwdABqEW917ULNbLijVgk3No+OuNHPqh5ffm0ZV7
u5R3eF3eZPt0JNP4dbv7eIeGm31R92QTh0idB4dvZoVucGpEENBdKuoLLCRDQOIQGTFBXH0RX68a
fqiyL63cJIi41bt9SHjoP9QHd7XFqpKsTXG7cethj4fTwSL1baJJQ9xLHb2mD7+ZbOAiDypBLL70
kWxyA/XCEaB+1Z49NHnouwTcMxQQKOhoHS+SAw7u+GIu2wMl5o3+q5LYlEDA1lfQTnzeeLD2ULDJ
VJZPye3PnrfpPuIE6C1eYuI5+pQloIKnP4reJGV24oJPpU2Kgcidny9HbJhJ5XaVyqK7Tqpkns93
sXqt7abp9OF/n3cjp5h4F4sRIMxYkWKZlzm83f7m+LWx25xp9ZC0QOPryF+4MvzjXj8c+Swqs0c4
Q4mhiHbOBvN1TouTpv8ICZNf+Ku2iho0Aa26x7W9gVQoF7OjXosNX5GMwu0qh6jufcp6rGuEAjFn
rLdr6s3eBtRHv34LIptx5gLmQkxVQloysE/MPl5VNCbUWEGsEvej/XT+Q4n7zXB+0v5mThQBpxzD
EKE3mz6iYPgQbmVFgk7zUQbPpXq36W8qfMLRfZOUyOZpZyzN2wvqGECcD+khbov8UFgWhh5jj6Cs
w+LxBIsm0JiR+Wx0O7PPSz54u8hQapS5KgZpmWTpxJWEMjc/9jujNa0DupO8bj9xqBeygNmNQMfg
LBGvMps+P6dFTPRXhbcP2JY4JZbu9vJ1gCJBCOiZInmtAVpjLmG9vQ+LS4/LTf2177000wwi3l1e
qTr45zC3qTkXHjyRzsUzZJi+uz3V8o4qV1aOVYsY+N1jEWM6k5TMF4uE+Bjf3Wn7AMB+U+kT7mzH
RPVgXMdBqYEelN6d39oxszgs4WMet7utiT/SY5Aty4sRb8MzDksb6AMfqG7Jw8SP9oNs+9Q5TvOF
XRaiio/1yyXWVO0TeHBoROh/XZbaHEppkETTA+7iTaI0gTGwNCMGcJjvVefuyiA8l+WgVEvgrFz3
7ylw3Tla4nU6HrUevfvBMu1pmKoMN0QNo09xAbo8ddqmjWTlhIIQ6M8YG9SnqzzIY+07CGHQJ1Wq
fmMYdJ8XOi1JunLcUTLPSIxyx+6InbiVpfrkOKMjROpdgcvDDbdsBYfh6PJhKbKkfgYxq7GofE3q
dOe1r9EUgVcKWUpkHNunqgfOSjqdN+zeOv3nIgbz6kVg7jD/1gPHHzqgDY1ehZqmKe0qAtxvY3Qt
swzpUHCm9rxLnLV8NrL448bKYgQUpw64Yjjoah22ReXqXIPNC9AokA78W8SvmbLiM395l97F9jyp
6hvV/nB2kkBvo/BjvpDHXJQ+Y7d3iI14gXGtiECj/5ZW5X5QxRK1UB8Qisu7/PRBzSajusb8ijwQ
xOPXomaRFG19LRi9qZP9HnqdR1/3ICGXLqy3HXLZ38chPZU6AQoQ3fg3Wd036JUtTIHJR9XI8+RW
ZcSfJVPbzQzqoVatRU79FoGERk7Fv0iiZjHMwQ/XOmqIl0NBThy9dddhO7RqroJ6mvMeeXuKZhdx
dqDQD6j1Xnb1HvIEXclpWbvvKLR6yLLM1RToBU7o+v0nf6fruyA59lAJUjw64H9Q1l47Kl5ikudD
Aqk7143rgAYuRlOQ34ZC1sWiSVc6RI/5xldpS1qhr8IcaLuwYnf4Ld4EzgYlUuTtUpyKDqiCy94M
Ro3IswPKJrAtM40BoxFDpRb7HdtDMttOFJ9CsSZJcztEIZVIogRGpa7ooN5zKWsZGpI5pJCvbaul
z1Ej/aoRkvDeshbrTo5uTXEX0zwxe12YCpmgVtX9d/pjFbMxXXo3z86oG1+6rNoxYqRLcvA06ezG
ZlSqDpaQfVkg/HJDT3Lic0gQrf3GgpMCDbb6xxuGlM+MTPsu2ag6RQVbk49ofudI01ZOENu7DbVb
rbiONQ03uZWlPSSeLq5p9LJBuvOd0SAcG7dfrf0QAbCvhHBc/CL0AkkPF7b/hFLr/AT4PKSgJVQj
yZi7XJ0ZPS0QDA5Lw1IzBXk3EqVJQFB5yXojOrKCpmOG1if422zValqG3SXBtODvRT6sgZdQ7T3D
f9+G1xkAx2jkk1cVjU7BhCETWnbcw0EdFwk/Wq9XyEN34BiX2DTzNMaDVO3w29DIWH8eIcB4Qg42
LQAMffd4VdIN0RBHlT3tvRM3zZCHqZwczv62ZyZ7dNAyjmcnjQJfxYoN7kdsWSGFu2Cf/+ZQxp4u
KtXetWwWYYziDQa98W3cKKm7oEfmLpa+oPwB8F2pmhOCu2iBIsjn/gjO539hr1NATZVEaDKoiWft
1BfCMmDnXTgYhLplpzmhfV7SGuwxHvJq5ikic7sfEkJqOoRm+HQ2ep2XrlP2Pxi3NyZRE1fdZgLx
NhSDJqxDcmKxhwIrNWley8gK5f83x3v581MMghdrm+vrM0I3041azUF4rFHH9Tj6VEO81ndEgYJ/
A5TFnNi/nuj4ozQX7/eT8I+O0/Fa6k2FMtfael0ckkHtKn3finaj8t27fbbKxFOhMLhj/OEJC/Ac
9rlyUKKOpUb8Cgh36nphgfutu2ecufa3kNtTNaaTnqm7fCLihGFAoEVz+SxHK76s1tPbjv/oBX9d
wQWCnfYuycx8iL842vA/tl1aNASicsgPhnLRB3yCvn/u1hUKjzoTDwpgXdm35imsp8KAKNBAb5qC
aPSyatQNqPXiFsdVGxqKDbFEydMtayHw4t3EC522xtNe2RstBpRZ/Sieqn6VzX5Fm11tjJrqLqCo
723Z9S9bbeAERA9q1++exsgQAQGUgUjXI366vbLs9cxqMSgnn/upJPIRnaemwR28yv6WflHKuIrE
yk9trkxPql7mdWcIKOS1ZgVq/9yNRJWQInQL3gvWBVFypXm9MDw8QyaaiVBN8xvfmk4gfmuc/R/M
OiTbbbXaUowEpF52X+nL5xo3jUgO6CtbcDeTNJ9Cuf8rX20N3c4pGy11zkuO1k+H1fZq8bS5aDPp
aavR9HviUkUp0Zj4PKEtc0F3H9rIRhqC1+g3h2wHV4VcMx4H3ezlar9cmwLT5OLFmAS+VuYBdhMB
4ryN9U7tXwUM+sXHcCtNB3U0S3TsUsKR/6bYfKQ3FBfEE9fU72Z68Upo0asgzHKr1aezGOzBI1Qc
RFQwqFBTEJLNCTb9HbNFS3UDeIsQ/Rl0ImU3u0IafZLjLmJODiRSPsGwiU+dIABKF+sRglIbvep/
gMax+zkGnmOXWGAcpM9vCNIzNfPXis3/FHQTARKovm6PLl4JxZ/C7hFMzm/c/rZz8XdxX7nD/Cbj
R3+j2ePedOle3xCFBbLAHDNofm4sf8zDfSPY8ZwEBt0OZ07wzZIQ574XWhcdZABCwJv4jPdz/3O/
Oei9DLxaWNnTO4gdeDiB6cQXgGWRGa6mCxES7SzrfMm+37Iv2Ijtc4B++Y1LCECXIghC5+7m9cAA
pFhix7l/ZClHp/8+9eXt7Cmv3EZnf2anqINx2ww5zEeWNRKrJqoz40fMkMN+V02VbKYJMHb7JZ79
878GWUr7T9fBsT1nd3VMa8LjWOzdlv1jamSN8tv8YrRwMtbLFiN7nrER49KfMgG8oZ41laRZRKoR
DyarzOIQffxN6Zv+Pg2b14kM0/ScFJl/xjsLy0oaEYU0R49d2r3/CJKcgXc9+zKsY0mHyJJzX/Fo
qXkLF2OkcbhnowbFi3FYINExJI24ud3+B/v3XtqL1KP+nmnm2JRDjAXOG4WvpIGuuqi5nYbx9YuH
lpjJBMp5Kvqu8/eE3/48CihMJSyL0PfKMCmWzsErJQSNVuPqkCL+ihWtMrlKDkQtzmQbCjsDx3Vw
BPinkuPO1UGVCzO20z0tJtZ3cscxWg8/YpkkV6/rQn8mzOIxyHMYMuHvUiciKL8ILVLIY8tJ21yq
PK4kmLuDkemLsFfy4lLQsETkjAfQ8rKnaZ0exWS5MACVakc+bFgb1CeJ4o+EEzFNTvBvJZiO7jQl
pXqXJRjozbAF+QI3GyIc16c3up5dPhR/quAUO9zRTUhij6IG1izjtla3RdiUb2jLIaUZi6ML7d9y
DU6e9ZJ058o7lTQ3CdIEW0YfjU6kIvmI8OoP927IhugySo2cHn7sSXGTy8f0ze5YJTXIY5TM1v9l
zLiLns9KG7Z8Z1ER4aVUMsFBoKKzfmllj+Sq7uvljuu6I8jexx6RiMyAy98Wc/sLrnZ0A3dJO19F
TMS1Kim2ZvSmpaidNpL1IasjND9VlGciVLBrnaMkyGzywh2F6OMMWQ6O/LAvGkdvE7VlzG60t4YY
+DMXrrz92jzUt2/DX9BYAtDN+S4IaMCtNuwQB09hNhCMQG8kOxtSM5SnzcRQGYmciKefIHDDI7vW
EzOZ+zk8TrFEInEcqcZ80aVa6+zhTrJ5/LBA51+p/PsZWCbx7DPd3/Hzx3BFb1NmnKl//p/1Mua/
8POHsplxx4vy/DZ51d322x0ruZKr6kFWdp5vVSMupycMucscUMupEVngvrDR08ld1NTD833DobvO
vtViUx4KvKMRu017dZwKhHkguyo4tJv2R9ptJX+DEOUsjJxt9Sf1W9Et/2mXxc0SdKRtJTyEwV1Y
9hkGleZefGStRqcDn/svEOwcSE4PhvcSWDMjx1IvK1GaYZXTQ1BKCBMvYFz7usoVP+05kx+EHzAt
T7nWaPRqLsBohBWB7NVrC0e2uwgSOuNSkkvpxcDxzDCZP3GEkiXnaN/cNnpg/k6B+t6ojKpFghs3
TFT/M1xrgLrSZw85X+5LdH2oitSp3I79dnjBOSPzzVniPSuZYrUOlGBSBH79dQYprv7iTFo+dcjO
tEJlDWgsPRDcyywVD+Pci+fOEBjXZQcp/+2W2OKn7ynccISMa1FoIqc571NLGmbsw+sLQTzf39kR
OCzPIlWyY9R2TF7rUy9mt1DRyNwzPN/6Vu7Wh14Sq0q0XewlFRWRqLKT3Jk+V8oADklnYuLkox3Q
x6plvAeQqpEZZMF/+CU/7c+OFRsyLh8TawEeShPZIxYXA1mNiT1pwR9/23h2Zr/NuD6yOLaSgNnn
zp6bmfSARQZ+j1762wxG2uEps0URuaOmSdAXw+AoSF3N1HD7fAyrbris7RtTLLXU4ln1xx9Cjsbn
a/3dZfOu8ZkcQue4UQAhSn+WP7J/EBQaSwwVA8oKuBtr9HmPw/KUrt/MLdDrD0BqsGamftzgNa5R
Hw/sdc1tcC2lTM5Xr+l8/r8qm7+aD7D72JJ5t58T/fDzoYhchXtAxDNBS8FhwsSLnnJXpBhd8jNM
0C07wz5Qp+xhGcf/dVcDPOOgM23XONgT0IRryyTd+s7Jqnpib4MZGXCT8TWJ38bibO0y3D07YG7+
IxVbi0n950fiHWk6tjX5/QkZavo7CfgcRlM+k0SGegY2mTMjV313SAvhuCAElUNtebj7XZxJHjBR
8eQTixFORJGq/D6ZuuQoyape7T9LmgQoYz/39vpAFYzttbod2sT30K6Tkwzm7Y4iNmfbAPwReHBd
wkLXqkB9fzZcYsHI4ejVEX5td+XUl4fws6b4KwpDHECU8dGsxz2Fm80TjJEzKsLuDTX0ugGoZ1Xu
2nvq+TJkeHt2qbv6xEE/Q03x2gHMSDCYgtkd/7MlIFYSjmYCe97j6u2b6p7xh4sZBnf84wH9+ydu
83PxOh+2mXP/BPfrrPaZ+MVBpskUIy6LHjeg9aGTHi89jdh3zE/oC844MGHspFh8wXB4H9bdcwqF
XyKTCEWPS3Gsh3iOpTAAauvZIgg+w2pR06D7Mi/ErZxmVJnvPXqbcswTTtzVhaKQYcy265jHYI9S
qKWX6VudZEKOlSu+L1Zs58Y+o9nl2oSZW2x6Hl4c8gcyFA0XrDU6pf+6W7y7NhoAzXM8wDfS/0PC
Wj7DngcBW2NdcQKEUDni9tSsDIT6dmF9l/NMHxlFlbesDvYUKYDwzW2lKs7dainkV68Og7zjd76r
22z8mKhePJ5sBQ0HYsnJM7m+x1Ryp2jp0Tm+MM56k0hrdl2tqqNWsZ04cM2kAQ6zakyOcnCgrtYz
TtgNJh+9A0vBiTg0Dq1ZuwHgH0xyXpLFIShbVySjaTd9yV3/CnwGdT/hM2rEVrib96SxsXI51eFP
TxRv86Woa/quhPtNXypuQs8emIcmu4Q3HeKfsaVsN2xWjNY1ZAZS/xMiWzvlsmxRvli1vMUyYqhm
UKEcECBG8HnHpFdBfUsqUBR0SU287s5ugBaZh8uOXm5jQPjNmnxtJEzIntlQ6SGrEWiYWsOL1Ao5
csllr6k7vThtoUTzyvIvJJMTFScMtJAUgn4WEpwjM/L/nsQ4c7ydnFgi4rtF2c4g2oUE4Zvxv1wo
M/devFO2SHDW2rtzkPCvPHZ1ZCfCV2bhOEZv3jFoaeah3uH+PoAmeMRANtK8MZNoDWy/zFd++IY5
s2HEP98uiLsqZgyo7jlDHVHJFvHqHxcH05TA3NxLOazpganb33bZ4iBfAlc4DNt0RWSYzsjLbq+f
lethi0YVsaNOWKMhb8LBk62nI8tTKRN0LlWsl76PlUe5lMuUOpsUaXIJHdllYosuDRVD85bK2OtK
1wWmaayj0vOhgufn9D1JsBaUl3BvDrRu3t6OKNwCVgs8PJc7UXFvhjRZ43TZdD7p0CQ5ScMYw4XB
G+CNPkLUO3UZJHBY5CfaEnA5/6src5bO6QntpvcC6DK45bbAM7QAeO3ooYf5mt7M+NIALXGPanvU
SZ11zdUlGWPc9kTEnaG2lrP00SOpFP2/tnPOenSXpWSiF6/yonrgCtBDTreNIUEHVfCTlRMtjX9M
DX5G/qjVXIwvz0wvjJgpAAGvf9hj+PHeW8sJ/RrKHkFXPaEbXDoKElSpFa0vRkpW/CKckKRyYK/i
wAaUYPLbk++fijcIl4PVYHh9pt+SrLmrmhOE1pEsvRZ+nT6aZIFASKjUAnPFOsBIY8zHKVotjZSI
LaYP9+qjF5Og2ZtVhzZh6OuIvZYvvrJ6M1FWVgVosRpt2MTItS+LE/UM/2G9NxNt11MN2rQo61v6
jDSUfgrR42aXuTpYrbCRkLftPHM30/gkZ1T41ylcmU/b+xF4Ukg2wBdnt8KfnA7Dms5/ZbVC1m9X
FkLfODeDQFypxMRF+w0tZZJzeEI0RwjnGZtt0BFomPCuAvU3KzcQzvmO+6ctLfuwTjZnBjWMpLHY
4szFfGsCH+OuVkcyNguB50zzxFRM51arkQb9IW2o5Gifhn8/J97RVsy/oedwicpzyRJRdd5gcQQW
eUbfw5ufjpuN8zVqkfMLGhVp7mZ+aVcKJ4Sd6HaLP5WwqtKedNozfBSWUOHfFP8hgWoEiXSCzQJ6
V2oYtg6n7JA+RItkYmR2ZJ8f1TVchNNQEXDrSAZXjV0aPEUjcUfi7tAyTvPfAokcRHtsDOcm/yw0
DrxvYNHuI2WJoF5HqWTW8B2doiOwYJLUUj8aPu0ecwvDG5j2e2dQ+EHnyhQKplRcRwT2ZmGP2DfZ
ghajKAErR+/sew+drCeCGL4I1ETxJ0/XckKH6evvo1/6z2Of1KiyDshQlEIv9BMOrTaH+iO9Y0oo
WD6gWdcyavVz4AdarOivNGUwTB1uO1olkM1glhOCwY2Kxm020fMbeXFL9R477uF8cr+We7+FJq/L
hWchyBlHqTAw/Dq4czX6D/NKbmS7T/ftI55NVOE4sunJN8gdLjLMdNDmQC0u/a2QDnmphRr2VuUD
dHxtqrArKVkm48z9m1yWRUZIVPKhipSbUisIXnXsVSd2pEqoVHtWArcHrivrIGe5S+fOtf72ioza
3Ihnq1rH/xZeuGP6c/uyXoipxLXwFQ8NKasDM66rG3XKsV8TqSCf1cKwUoxXKya8G9JG6k3bTo8q
5AF0Dn5fXuzIa/vCmp/tVaHSQgEiTxMs8KkuQCVabWRflTG9TSi90HbqeobBJ7z5Fw9gAdZ76Hh0
sUYxqPhXiEUeSgnUO6lDj24iT7OJzbaGcyR8qHNNbSM8ka1CAiphq7p7fb/b1kFqrMETv6L0HvjE
WcTTmXvC+pPC0ED5yrOPaGoJzctMQMEzfIVIvN1qa/OfWHRtcwMF6dzXsn/NR38HZckz7kT6oVZy
qSPXM/hsYQdY2PHz+GESPwCUFSE+D8c6j3xvDJHqqDz8gsRaEgmAOHhYbL8abPiDDhQP2X1lqv0X
QLd74CszqZgEmIZ/VNPclMhHVHnPY2YN8xsYFm1UGjmVc00gJ4rOzVZcam44jljA7/VZkdpRorHZ
GGaOAsW4KdNpOAf7E/BNjuZ2E5r0BcCCaNu25IYiwXMQ/scUNVnfx2Fl65CC3vjIK2lbtFZ2h+dN
R4HVNHDZhHbOGx0z/3Si+350f/NZQUqM6qbr58APADoGS7GIneSYsY4mJb/jUHZEIwBTopuzGOa5
6ue/pfWLzFHqLKs9ly+8qQg/ujQ1bsZx98MFUVPEPv+b+PIwdeq7cTMrkUOSWw6HKxuGnI3TyaoQ
EqP4/6fu9eBWs8mUH7uI3E4zWIZ8mRL75RXZlZ3WhQvUNSDy0ZfuhRN5FlMHz8z3BE4WBLPEvsI/
wLWDaZmqGkAZf/J9okbao4NwIWKyeekLtIPi4D+Le99bZsKywtVeTJT9HBsrvBsiEZZmxmr5EfqV
QYD8T/djhUSclMpdOfP7MostF8ToaqYSeFOrrWehXtKlPqLvHVZSwnMseewjWaL2UkjMM54E5aLt
LGZc+5PjvaOO+nFTk+nWGLxAJW/cg+nUFDctWvymVQXzBZpWpuIFqvQoJUSm8M5oj/0EV5rd/Cqi
kQzaxJcpQaIhZpdrxCsOpAex0y1lw/aEuaAq3Gpey38RJ0eSXkDxBlZJQCmI86qGZrweGiZkbH1v
I5ySOsV+NmPxCFBkkA0DpOr6TGqi0pvhdLqAzdPVjngbjxgAQ9tepSBxLFqqRbFCG7DZEsZK2Z+I
nGGAjZYh2G+Rrpwb5uOKwivYfb5hPi0uSSve3ifYZGqajNMZj/0+/DuCBt0T7AyfXni9iQcpc6JT
5+koN5h533/0kXw+vTmxgC1Kl0wnjyWg4FyYHsyv+oTOKzIy1VdU+t7CdWEh7W9dtrPrsP/RxBTu
yUaiH8pSwUpfeXk8J7/VxDnLPUBu+Lli65GsdLR0bnKUUTAbVImD8fG5vUbYijtNHaDZUdUUD1ad
gP/rC5a7zQdQ51GJq0NCD2oj97KM3mam1UKKtcE9gIe9CUvlyPYe6arIjmo2nIM/UDa5z3DV3kNL
OoAPT6L0WWk9+7q1gLQry6gesNJcyONxgJMM1Z65sh4g4p9XKonrNqZCYMpCrin1gm5vuu7z+lS6
q4YfDyAEIkgPClntwJ7q6hQ2HHXajTl0xUV2+3DsXnJAPEwjaZdyfdPnvp+lOP6q6JfXoX81sUZW
VmHIVpzz7sVPXSUPc+iYwez5/r9ljkBahowtuVQ0iiAeGF5xJ0Wyeu33shCMMVNZz15L4QbNsvQH
ISE10bYZEkx2naTjdD3Zh9pJrz6oLB1M4Ma4mhUheczG++zE5oLCtdntYoZRPaSBL/Eo5Ad1nT9V
LP320BKsKNZMd5UitroeGK3fTMArxJHKN5uNMa/mNRmJcf45l0KDRo8Rtnsf4FAgTg54c4GL5YOf
bg42Kz/d4ZDI06d9C2nILdu56Rdt9EIdY5199nVQYeTNf2c+yJSIULI9iSNzgdsN5ZlaQPiftzVQ
RiL4Nu21f2ADxp8FgGPC+A4aIyD72TZJALL7kTGWzljAiRS49bOjVz0X2OKRKfRtsi6WWGzNXlXc
xmHEDaef1TIR+QL4Ahsqe44lMPK03a6EmZR0yDfWH7IlscynnxkJmHSnHdJ5h5FN2qjPMh4S8jaQ
UAlocPO6RIUegLaCwKdoXnzC6on0YoQkDdpE8zhz/Qdu8n97FNNDxXFvXA1LNSBR2KC1fBdSj3oH
k/WqQrJWwSrz0nmvnzT9FaA2+cHXxGZmRKarNVwyIrtWdnCXQXA6hfW4S3jD+ZRLyYP2fqRbrPiQ
0u110rtMuzsLM/we5o7VsZVWL8btPAP1YRQcbRhgGBITfYnsEQas77A/OQYwaR9JR2iY4uPRHc2M
y3hNjlhrorU9UUF/x7IOGyjHds7/7Hej/EUMpgI7oCpDKVmwDwx89VeScYak/tkd0aVoy/MQ7aQD
ZLYPPVCLQiuASULtUWT1NGXzzWuPP6vS6McVIiYg3X9t/sI5Pmx1/C0DP46019QrpyXJJiqXSs12
zhQUpcMZLyKKGroa5WXuK/XRr6psCm5v/OAfH2mLZXFilFkAAA/cneHBCHTwPgvPanyv8Mf1Geqp
fxiKJ+uihhqZGrdhgHtcMjRDnYZSmDxWhnCCYbitL7j9DMECERXaCb3FCpZHboWQdzekBvVCrcsR
dSz9+QXN44X7fdoEFYylpjVwSsX510aCN5aG7J9wOvyZSppgZCshuzkaL35Jfax5Q0GsU+Wfomdd
84CwMA03sIHeGNQ9jVosfYT+ntz7VnM0cH08XH7jmONTVynmJgFhGUFex5SHWN0+J3xTDVoi+sd7
a39Bfm/BmaFw5HcdNP9WEeq0W3rxW8IMKTI7DyVSVye2HXbG8+++Q5IwWRN4D8l70KbsCVI8jwFv
gzZ/bCrU5BVJ8Pvb2MnMFANeUYeUIbRuRHbHiM4m+zt3PNYN4qNDgr+b+Ht6s+j4T3x4Z+5ppYct
zrfSB1EZLPQ19wR84hna5UtM+hW700HpCVFR541FFF2diKHpKavmyBgMFzBlRGin9gPDQb08WGGj
Kgkn7F2ZcAGSa68LHxKb9u1rsBQryM0cEiSDMLQrwQ8z02XDi9iAe91nxjUEeiMm0HoczDOLjkL0
e47d94wOtwdeHZROZ3KvrdUKd/LE4QA/ty9M9jlUK9+BqDGGehKuImG/AmKYM2kRvDlT8v+JVa03
YkN3OYqft4Ae8oabQBk3MOOTBCABEDFTdq07ROUvPALBjeaE2H+Kkzy7LtQaJncqjpxwOAqBKX3k
MYQBQaIvQTt2HTNFPT//9I4jsaYQFY102UugVIc+C+z2AENWnSr+1Cqf99xvAucwDXheB6ZjBJmj
/HtA0oloYuFh8AS7uzFINk1rFiQQ9eatbFnBUaRJihWwRvUcIffzfekVAtgGPjf8vJGfrAQzHZzM
hz/GXxPPZjQ1/xUIqZQEQRWSi6T1cU+Q0DS9cOGfsSnQxAFd/Ol3BX1ElNWSzwbWIyemXNcNJRFR
jPek0zxsPIk/X+XlZe9Xmmb0SgwWJOUvsFxzLCe/XgBCjkFfLoyM9wUMxq3O1l1a8sKvPc+qIFys
IfcNTJrQ8YoV5mxF5teUA0TIPksC06bHoAdsxPqQFpxEJ1fUn1mfF3nDEnJvkZvKAaK8MjKm8UQj
85TqMJ6hPoOID96/elEh3YZzN+K5r8mv8GXLqSYE/8XE6gpFKqW02M9xRz0syygRME3X/exYTL3F
YExYZ8EwPIe/iRaN1AdG5+Hy1pFqSHIsvIEYAHEMFRJS6HRkiz7BXQKfvRnFAzf1mPm8/tGu0Iag
KdbuICnzeZtWrcIe4mLjr2WctNxdAyryRc0oaDH5CbN/NXunOrSud+bYXTxT6hY4rAS+sKVn8f7H
2AlntWzMCDJNDtFaQWo3aZ60TH8VrHi0SawJo0reODmqaTeMnVHfczgFFejRdtml1ALm2BmVfvMi
Mjo48clQ/qM2nlPBMV2oQ/g7A65Gje7mMUVQMQe3YhQe0RcUr7cETCKfY5MS1h5wOwRZcahUO5Br
KHvgJkZvn1Jeuo8unrmJMTAziPM5RatCDKPJN+fJ0KaQD+8tTeisxblLYH5eTBRygyPxoZpD2TEE
JavxkRDSXCIu80giTDRJQSxr7L7t6ch8R/eqeb/O37RDDxwir8jqidMykRx9w8ll5OJzFwi1a8cK
/oP1XlJOTr4xbNXpZNIz1psofvA3EkEjSqEq1Qaow0hoEaZQ+HRYwQgelRsBtipXSYxHdQguamhR
L/D7dUjQEZsjakrTVVFADiV+MySI/682TiVwPnPpt5an/nXHfCUgYXrAMbrqbMs5rTd2Qj1k7N3n
mmOKvyi0QvSCcylhMiQKi42RE4EBY0N0ZxBUK7pFa40qxgo9WdB37FWuq54U2JcSjEbNmePoe72e
1hbleYunorbsporTNwnrtXqb/5y1AL89ss4fjnmuIEVSpTBN1bXcLMDvPQX3cHfSg0TTUAiwVX/X
GmykZLiaSFbABIhsNc8dHg83EBdgQbzq/7qJG4fV89oM4KpCoRq30faJckFYBthj7O56t8jUUk2e
Qbif0G/zs5oC02lb3lLqy7o6/NY1SfcyRQ1wKIIEt87M2VGRZlEfRbpcmetfcrZs/H2Y1m4TYOqq
9JyL4ll1hRVswhLKaLmg9XiYH4hDEr6den85k8KsCEzAFrbBk4ZQ5nvHyyX7sxO9K1sEF4o6Y5U1
JArcXQzrF+JyboKsGXHyk2sUdLfsam6PkohQOUV/KXFsrL25D6raNleWtnK1Eiex1tGEJbEAJZFd
3vTpSLCRAElVd3GXlj5jNBgTDbO8woXt8690vrFfevW33SAwUB5JBXrH3f39VPQByyF2Z0g5Orm9
Qm4FegLIt3nkM4+vAYYhg3Pr+4mtEdNfnhMNRUzwVW3+3Bsqm+c2l7RxdmcO7g+2IF18adO/Vn4W
7ico+GL3dHg3Bb1xrQ/bTTIYGrmUJUr0XgT45jQNjbr3mOfW/bZPLWK7OJlLhSAK1J5cQfCaIojg
8Pog5JZTq8Ge8r0OkKnCmRVUFXCLrhdGfGuVHLS3Rk0fUiHMtfGPbMAyNmBg0s0ampu1MUMkDhdO
yreLPkj2JAIm0KbL42Ynvw7V+rWHymotaLqnga11kum2QeF8SQwrzXibE9rj/e0Yo+y0AGgdSBeG
wTcSuta2Umnl6u7w2dWTMP2fopPqTdP4PK/jb6gontfkJAoDyJcBjvfc+R9rEEz5snyXgmXD9bt9
aOazdLpei5np9/tKRnIAV02YP09eACl2T0ZzcUuXFRa2vtyGczKiuTAYQ88xy+thIDs3aKF4A4rM
mIbc9tZCo7WLPx0cWl+m35/rJGRPoZHBuHIhSjNn8kgXrgGBXTTJ9oYPhiYe7JWXuIDIPZJygDyk
uNZlF6MWaVFJhHdH4IHtYJX/7nQTvkp0D7mu31YBmzcqTRY13NmFK3o727/Dn/Yt4HnqAqq/zkWN
uKxbOs70AnPfdtxuH4eD2c2PKYfAQyQQWM4motWWM9ifEmtUEyi+dPBK2LP7yDmQ+sFk4xiRZ4AN
wmeuKXTZ7iCDQbIcRkCljnk8p/HqwLBwxCPwKWUDlS7j55PgXZR63nM1oDTkvUuXzxrzE4mEnbpz
gA1yUpLaKPssaNBD9J2AmhS8SRaVu8Yfdno+ObTVjzTtBPJEsXbKZmj0gl3vhx+3xvlyO614KSid
tEN9Y87T2Ci99daTpoFL92lT5ESqswj1OK1vqPz7eWqDdnM+dV/5A97v3GmIpljY4iSEdYp8XmyG
mZpqKK0wNMmNkbvdlR9T3RcCNAmPFOYcyQagyrnra7mr1fdEvxXYeU6giigmI4OnWeWpyDrvlL7o
vuWPt3uem7O2+3NPXhIEoRyQr2vRhS0EK/61NXKjGB5nWNNgRv59K9z5IntkSnUqpZLfnYCsJWr/
5erRwLadTQ5BP96CGyTAmZTzvdDLIi3OvvsDaYVxB5Wgb6KM+iRg6zGsV18wdguXh52jY4M2PH7J
jmMTFzAtNDOI9Fa+jBVi3btmmwsvrJwrLvVWyOIJi1XaZ6xTHlxVjh5K9FZ1Lfy2kPB8+3Hc2hC5
AKr09dagQETUXlazJHVZbEfOgrGqXoXsyQf1GGrB/G/q5cGY7P87Mo6rwLOtNu/Ks5v7Is84+5a4
iawWko7CK5FQ2out00iKNfTOfnAsMHVu0x+DB335Pw21VUDWe5mQHz37Tx3f/EkKrnABtzwbUT/A
T48e43QHXvJRK9sgiZhECzLa/4EmWbbtFYRRRAphx/OlApx/r430bN5bmgIdMQIm4Wx5UWIKej36
XBgVuQ1JLtWP26OF9A+aTE4podOBap/QNPdYRFw2NtmI3f8c6DcQtIaFbarGxHqEAmpUGRJW3vDE
fxqyvEHrNUsQmhwlBCJGSd9i41HpkUh7Cx/QbQSwVt616qC8H7+T+ftghAIF2NRXvI7itePc5pP6
i5iDElxU0h8yb7yHQt6rtTHLNeW3hsrOXp5xaIZhCvgHE2fMOgQfOWH/NNN5dJEGCnymuyympkKt
ln8RJHm7XeACJJwYQQig4IwDZKUwWvIL2SaED6T80mm7PY8Si2GVIPB7JexQwdXNZ07Ojime7++P
J91/j4rTrD191zuqj7E+qw2EAerXf5K1PrJ9S7fMrxc4VOK5+ziIMY4M7Z8tqXCKGkjEz3NM6RF8
z71tPZY+BKTw+P4U0IfWtzyhH/ww8R+8grwCCJOa2Xg6PMqtL7TwyDbc/Wuv7yl7aYedHMTF8s8c
pnvVdD87oN19OgDs+4mVT+x4GmSC+iZyczBBwWy9LuymJdJwZU6jt/MsgFB6o9sESSitJJH3kO+q
qqHU2gEhLtBOICFAsX+BmVp40NmuZz4+YHmkG93tjPH4dUlwKauW4FztxK1OWBJGfPUvnGriNMSf
87tcTcy9SGlSzEMgvxGcFAYK4aHoktpzYnrTcJnf7Gapy3cNHxQ25tNTfxk/U/YYhf/ph+F6NBkV
1grs/mVmzMPCo6OqwsC9jGNkRKJ9raPy7BZgs0iDy20EjIftOhNLaGZQTNW+mcNuD2XqAiGtrjKc
9NGQ9fv0QMgFBfJUs5lkIdpjqlAwdthNt9w19wavYAYKfPsiybP16LXb6LIjL0CEZYofqswWil/y
/+E8/R/PnAXBl5fs5LjYuT90d5Ykv0hv2jWstNKlgr8ulW4NYJRi0aglALtEqKwGWS8qXWaQ1OX5
bfRZ+RWP5js0hYUzk944JrJIxEICnFVvOlMTtgFinT73u0afsHRh0DNrAbPZb9Bui3pZvL/qeKF0
fK7rqUQ0Dr9AeAmY9OYE94Cj2b4ErfXIi6/PnGyrVvTSCC58PcnlPVqPguLn9pTvpaB9GD0TVmK/
WVMyROqmdEpOvXGtt44rwTkl+6Xs5ahdU9HyG7NzL7esK3Fs9ROLzXK/lC9rBbnYfAeXXx9ZHdcx
XImMZBLkHTZRGpkv4cRW0xrLdy2YcFMBdOSBhkJriY8f8+EkKQzcILwFT/vi4pQIVl8p2r+5LqRI
Fzv9HMYQI/G8CVzNkilj1SFnHlX9kSiCBVsKKHMXSpFVONaIXXGQvTHTaYk1cQvUNrXCdy+wDkNU
JVc4rQz0SxVv2pnckl5oPtPRiIR0tsh/8A9d7msNrJIMNyKsGnJMHsmbhbQq6M+gj76VxiFgg8J9
LuIQN3IZkFjIgVUVzBq1/VfI3aGqSapYOPvxY7Nr8HaiUSIS2d82FFS26EKyhp6I+klVKGoRLR++
s7VGygI1utgBrH+G4AIyso/KfBzTRokX5w4esX+RDhfcB7Wbu0azhKstFH0v3UD6y7x20i7Cw/jK
r5B7/3aohXXVFrp2fi4CeawdEr9z3qZoauGHPpsRFyxYbZevLGARea/vpS/1YWVMxKV7PtaJ571A
XIID0YxEnBbiBPFsqMR8Ukw3maZH3/5DivpDg7UHCZwHP5RZmNrzmyS5tvMVDiwwCoeDIpCs2AvZ
0ZkETtv+STum7aTslBnUjA2h5mO6vLqT1qukUnlXRwXoqz6EJApkrZqaIGa8o2LJ7Mi4+7qESmLO
9XYqvCD5e0OtpDTNhCTOU1gWNeMP2xJTtfgBaYAX3TEizkngE6omjrYFZIrZK5g7fO2uUYC8H2n1
s1qgeq5Hz6OSm5vgBdIgKac7AcngigCKOmSKc9ajb4KX1D4um8P4/Jajb7gJ4FRT1Ex+bciCQwD8
ZlQXwSMUHhkXJI27LM+CkCJBvwC/YfbPpvBF9d9bibkK0hR2B/qmeTnwEIUBFkQ2Fj0PBXHWF7oe
z6pN1zUj4/5BgD/ufQKrBBpUE0F2O/ncg24Duujw1hNacxdGyjOsLC2X3cjV9ARUT9/Q7RxJM04y
qwJ11qyLZI9zhveGZuLkF9ViJP8FRb5JGjEvsL3fwntf4jqldsiFuFLCgSk8vssYeSody7UlJqmx
Ln6tBoCi+dkCZWP9irt0WZIBiA8B+fqRqMD1mU9/nkOPOPN5f/hDqpugEQg3NVqVVNSj5v0o9mjs
81lHBssEpY7X9y7Xd+NnVt1DSrrLVSqaWBOD2ju814fWJmNhS9CP5Obm9BudjSgtU5715rH4lifZ
pnufr99cp8tTq+bpy5atAA6pPbwJyytNyeDosUWTmfy1+w0vfLNMYqBL/GZhUibzQ9dKadln9mpf
bk8pcQa4mbNCTCdvk+sTcibZVb9kWpz1mh63rrwk6N7d2TkIvGePRVWKzU/uIZ3uJVrVW81JZpdI
u8MBiw1cvbBonZGYCi+reDdnkWGtX8TFGv3SPiRwXcYv4Irs7RyWCSH5gfJWqMzKhTEd1gmowiQm
8RWlXcqq/5kmonzI9ZXsGNavhC1v9a74mqnsTv5KBFOIPdIewUrhmUG7spItBLHhrym3S/RuVdTc
s6lVIjlKRnHquxOId58QbSylocerUZavXaKFFyl+GLl1ZC4o37ZpxHTM1dV2zA2IG+8+LH3JX4Et
Kw16u1WWbWGND+dd6+Lnygbpono0Ox+WZ28HNhN5T+Gxjd5N0NEE6Tnf28iVnGy38NAjM+enONyB
XbU0KDcZX0Cuk2HzhWuFONf9o6Re0JManBAUXBhnJ4cwJ2opndCAe5fFw8Fm4Ldp/AMPm2tc+ZgG
JlEcZz7P1HFGS3IASREfjyhfnWvXf4EU189s+cT4gR2Ple07YolFQuPWVNMcKpjd5XrtZ8wZeh7L
yhJz70xDVg5hMpFzbfJXdmmo/1MkrZDApCTxewPoLP3zN0m5RatxphBiz/YLgVE1zZo/M/yARRqO
AxzJlQhFmgRFCVxqCU8Fa8wwjfxZTuuy0RdnAG5PT89TXSrQJsduSmWRQG2sVCquB0yf3kWnz5rW
U/JEwMPYxdD6hpQbcIKA0jjLJNXZc+BPjDQgUStT4NvaRmF625cEYijNc+EUXQIFRoUw8ytu7NP2
/2i8c/vYgBvUcWT7sn3lsgNO9fabMKOvT8SEwoidpQfXAZLDEf507GoWgvrjSuevimcV4ei8R7B7
7fRnXEGNfVedUO8Dc2GhEr0nPqEygDo1BpvMkPm9WsHn3XNrg0YxQ1PCVduoyZT83uP6DSMTeESv
Yjzq9c6a6AmEmO1LSCZpppJLhVqAstUT+N8phvRa8X+vRfU/16nt2WZE3902hCDiAE1cL+Sic8Mw
bj14N7sUSivvMNMZeSzaJmTQyyXvwLn53ttHLJjVJdkku9iHZF3WXoeS/pOwaYKuT9ErgMaJS051
bzUL3h5DgTStM4rR6eMg+qYZiUISy/biRPJBjyFl+lygScXFFAdAs8Z+9lHCDi7ZuKmSJ/lIywZP
TojCE/pfbKaRzm79vtMq0PbJQ+mw3G0PZYOUYjHH82yWZy0fZ5r3Tra6pRtF0yCIeBs6z96lRI+s
0ZAJqhS65mp7dKwYjou/4wWXNm1RPwbcpjvxkHN3NpRFMeSHSywViDzA0kgqQ2yqzHW1nltvahzy
ZLV14uj82vaeQXDcP2ABW0OKKgmXHj8wZTI2Q5LFLPcJ6SxRpGG0pT4EmZQV+NGuGEcwwbaAysvL
UmmnyM86yLqpDCRFZsxCVrUqi3Zfq0puXgDBud3dntZiDdCv3Tmhb0h4itLEdp/JAG+FicRP8lkG
TEXtxkmdDhe5/F2yQQJq8GOnblN9Gp8/SpCXjU/un4WJKYNurip80mmMXkiGJA9jfvEt5DQNPyIi
vNk1385P8AG2ghejp3VLOIYri9buhzhvfcHMDCmFKMasDFfdfeUVG+63WS0XL0M9tZ6+EGajj0Tz
RqMrmuF+uoi8iO+zEmGVC1aJpO8nYp9SDZL1bl7nv2Eh8z8ZFxfcc4au4wrG2nqQTR/a5JivqjlJ
PVj++5iMx/aZ+OJKR/HHRmiRR8SYHjbs1GOwq9b9WhWgse/iXhKGPaPJpQEG6readhuMkl1cvIjf
9bIpMgdQ14m0GDsJFsTykI+d9up5ispyGOLw/BRdXyVwxmzh9zoLoJ/PA4GfC1gjtyZGh8G6rMSI
rvcvWxPvPz8z9YWWrMC9NDPVJRzIXgo1VJEvDjokX5szUVxjeX0LOLI+gfpcTfg4onEbWc/dBbxN
/21nZDbrhPz/uvJVDX7wl2p/uJXQw+730ZpQuNBjQ5eTtfrg1lus+wpG2fAAvQQDQZk+G0e6T3Jj
GIxHSEgwbOdCzMewFIXZPh1sMnXnO7F1Fv+Oj0ctPBtnpmONOgogxKzvEkYjRMKBjn8KQ/kQtE8/
PDtK59dLdxMnYXjFm07mCPuz0oX5x/d5jtlxwt5QuXboF584lbk4pG5OVriRaOGNyCFmMbSzWKgI
pG2Dm51Jf7jw4CawHqb+Nu/s9odvSP2uyuJgdfXmvsZ5FeDkfeBMKHstfMMcCFag54lvkVcNQzQB
SwhIJHJzSGjUDNnor7ZDM6Hm60y/Z3XPQWDtxe2tasSFW8ZpSLjv/pmRBwhNuqALENiolBieUVov
usbBBywpgw1CjzRWFYXQg4NbSnSEjt137zXuSMLXN1sO332v87REVyPz3cws10X5KQ8mr6msZ0ek
IesIntvgZ6LSSPvzf7ljwxKh/m4qtGcQkSChmPMubD0GSotIhf1lTP5wqxplVB3pwUhSM+gRrIMf
UVou1MMGfdwFVBX6NbHDb1AMNwmUSTA6AAp1rZdhyMY7i0uQYo0ov/CMoD59yZotLDidFGoy4Iyo
ENpLEvuwXk0AKZIqUw1MtNrvnHM710FcEnbmafJ6Z5kCvjmgViYhAXLHFOZ7bYDn68ija/SJvDlh
yZw1F5B3T4S2BfmYEuyzy09ERd5eE62OMZr/bBeTiJ0flC+CB/4QvbEw/bEvcqWL5e8bQyddkZt7
ugiMCA+qSsZcO+wOyss+69TWHk+VxzSC9bhPmvKnV1L5hu9jIqOxNNm0jUjP5oDd37zVDt6O8Jm8
tZ7eipytOY60nO2Yp/hYmdwSk89dP5AkKW41ACgRcaWOTWknIU3aUSlAxBpGap2eQzDQcvQsdQoY
1AlArDt3S2s1UZta467NP8j8hgjf/8W4BOo0VMK7HMzE12R7yhHpD6ZGtAVu4inoqMvC1Dms8ehc
FiLcAPA6PzUt/29deS4rrKt0OgcQe1/+bjkph+69ZgpDScC1uG3CdEhSaGy05NiaXGU0Cq40nkqm
ygVGcP5YV7f0PKViTXOrh/i8v6mMs/iLNZknU9Z8sVc3vE0eBiiFjO+DUnnLWfP0MFdtJ+Vg9ybv
i9AzDwEtBaoCOk1IJ2efcujIfDKMg27b2Xf8ZnEtci63tALWonX0ixpuj4HrgRuoDw4ssZrRUh65
WdEpk6Pq1tNbSmJIqO/IM/InicgDs00jKQdX4AOskF1bFruMXIoXTKeZu0xUaPqKKNnN4scX/mhe
psmHSVGh4n4PYTbRVytp6sgKUVRwyzxqZM4sdkzg4GvKEdPCQnBB3ZukJNVQyjPTxg6lSbFGRoh3
5F18mVBV1JHaviY6/2ZLjxeFZv447fmxnxvECV9Yl8tr+yPVMfxIT7FUNUBRVXRZa7WRTTtWm/0x
qquyH47IkHh2IOXLK0tzftTvg2jTnHS++3BDiOIPiSoMTJ+ZLmMwKC3q6VJJON6EKZiUfTqgnoOv
JZEXQrVml/qNxHZ5GFBbNWaYIXy33cXEEcmZx9P1Uk+uRbzuxdzrdQDwwGSw1i48Gs//48DdD1y0
a/8OG8+xP2JHIlfoQBgmXX0rjt/Dtr1a62hHsb5e0RwoWU2+iJArBdimwlCfWn4DQ5hkU3xyG9DA
6W4MJRbQe5y+H9a3PiOnxp3EXg1DP5Le4MsK0zd70ZWmuGgEvmC7ZHeVFB1uaBH9P3S6FNyvkZLs
EecU05Dvkd/MB9lUz7pyAKLCFSJWWD7UwbFQABb8C/C/pwv1Q/5ZYirPFy8fL7TtYlBs5OnkqS4b
TdLje6gzXv/gY3JBhj/2J1iUyS5kdd9yYIy3MUXvoOWEL71rQ70Wo3UKWsRwAe5F8WMewrqQwoie
9RRn0DV3W4vv5r7R+CdBJTOVRCdOUb47ue96LwF44+7+Zo3bIul2y5kv6abcjVU3aTHKZiIllRHv
rE/GQ3OgU++5cJnp00nCSI/whJJ5VhJgzOQMd4Ee2UcMhx/1XJe8DzvgwaiW6JVnwSuTzkSlBjuT
wk3jQX5dXDVuSUJrygqK+0g7tXgkj67r6YA+Mn1ZS3aSVXEoSTwBWN/COG+gdRjoIpFP4x+K2fo5
GP/ymB5OCX0QnTyBoLqEjQMu2wkD7w0JhQljs3uR+SduQ0EAUshW/B+IQu8cKeXy/a9+g+RT7mag
SdyCnFiqIrcIipoa2kvC2rAvCb6UresQJmlG0f3R5UXfPTdnjWdwafGXR889ol4s3UiK+4rj+QrB
Bhfbt7LBgvNZWBL4feMUjQj3gST4AhEC3bjHaPThEQOo1tZ8yjwfkzDYcsvFa2D/uS3VolnTQKIt
nUeHsvw1aT1oB2DTNzNjbQPcEIi04DFV3K+FM5HWEsXRqS+eLluQzvjwLdlWmigPkkLmNeMuIwHP
aqxaKM+3axW3KNTlUSoZrWqoSeYH1idoOKzVWWdiwOT356PnHMrB0YrUKqyzsDx9hSya31rdWX89
B2QvHNGDQyUT/5S7917EIFxHcv+dJjklb7yuPjgEj8qjoeA75Q1kiCS1FHMVS3SBJcHGfdScZID5
jxyePP/mcwwAsCkjkzED/k4CcXs5rrzBojg2hMLGKM2wzGhXmMCdShcI8SHOIu+JgmRsaAGv5kHH
QLeEMDLwrxyYviy6ONYQvCN0K8OxWz0sKc92qrR3tV4mYR/FJfQFOcKMxrdGFrSR5mv81Tkql9vk
8Gdx3P9f1ezs7j3938swkLZBNLBUGgkroZQHTY1XhaqS4B5dBKy/dnTV48P676Uo0+JjH1yADDOM
4OUubOZD6iYpqWBVG9Z2MffwGzeCaYkvr3UebAryFkuD2qGuVcIFGDaqkjrVGjTNv5Dat3n7Grbp
6xvMN3RNtAIvbQRZrKMn/TeDbPZt1bxzg+EY9RL0wlhJ0dRmEq1T4zVtcqkx3yVVwC/gR68piVbe
cWYTtejpZt4WJ0seREqnGNn9qRrOBlaHBNm6L0kD5fN/JtjVAieIzzoIZquL30FACw0n1wlDxl92
Kdy9PHniZmfYTU87vkYdttprt/oEIjCd9LTm7FvnhkLBpMyDQLitS+eP25TFK223tYtThRsg+WOR
W78lADvARkqwgk5wSNCyRPknPrPrOIEZ8gnHaiMISZyVBxPa8L1WghCk72h0y8Qge51tgMYE6biD
PVXp4VjDxmmmmkvbmHvyjaof0ioUAOzH58vQeCV1xtWrBSm6QmTFbYoZW1xfX4PZU1rM/6tSpUt7
hhkmURGc0Fea4Cp9o7hrzqY8jW/UmqJh+XCmDW8abZqMweqHxm0WEFNnm0MfmpIdxbJzLaNAEOEQ
MmQ37ZHP+Tmd+k5/DzURG3W2ho/M+j0zsgXg/Jf7p9cT1oKy6j7Wbmrs4PQLkw4NnS/tX6Dg+AlG
LC/XKMVSetpjd1tDkZIoCfyEX5rJNYlb1W+hsVESb1QVaz8O9XRzc4BuAcdv/bQ06PyKpfkMYNvF
Wcbk3TKkFqgZ6ATgNYK7lzlH0cckodG1NhhvirEpVHi3Vbxog/+AhQYHIQhIoUiqkuViFAMpKx9b
YmshW6h/jCNUXvlVrAVFwNKSkqx4wVzS8+qT/oVAn/XfmICTdinydSqDvK988FO1v+BWlXgM3eeD
DS2ymP9F7j24k+Qm4za61RGT+2X46n1gT+g/+LG6n/RqbGuifM1tO+dD1tVg5oEA+0trbKMGwUQG
+0mnrFdrXP5o7dsCdxoNW14LnvkpAw+VQWcK7Ihh48CTiMIsk4OfI6uuBXLBBCLrrW267WRY1u4l
xjqus095PflHVKByM+8itWDHFzszbcckt/ZaZw0UtrETN4CETtHoR0PThjbhEIWfK/6mjsstlzHz
0O1dBiVYD1AmWgobAWMrs++nF7o/Zw3o9hY2VVqZSX45Ero50DmGQ8PAaKo0U9fp/dxfAvEgdQdz
1avRU3aC6kFOpJmsaji/mt4LmwgWqLXGGN9qZDeuz1OcxV2YN5qh9ITgd5bHWPpiZWJ6jS/OYWCc
YJJr2kPVgtWFiA4+4A6qZy/YUUcaVoKMddCgrOgrU36ZF7qSo0k7kGzGabOw8XJ5Yfw3UOgteQ80
XI+uElSrJ3Fx3hyxg4AOLfDOTrUH42odVHbj9EIoVppTjf2FyRj6g23iWiIPZRkRuZ+GxFkbKaeS
XGpKPOyXD3PGEXK6BIOQB5d89oT/csPUsPZr9aZTWI00zCa78JT+c7PK1P4agcoKDjwdCjVM1k9/
+hK0cLBeWB2YloDmXR9bsg4zbnhdEKLMskQXvSBfKL7EL1/weHjBuOJO5heJfLy4P5u5z0HcQwKv
gNpy4DwvHIFXA1t2rW7wDTtLwBgy2RA6QULGrIVUjMTEg17O+Tzt+2w6iynWw8j8FlmxMJyctIQX
TBqprA5cihodSbNX51eWHeGC8ndKewOOKTLJw66QN/6wWaYTvk3f9D47GOCb+pMMKdonl8cbIUhF
Nzhyob5Ls4K46yVrdNrNLiPKN8VFQKgFduQhLqbdpqKc6iWRUQ975/q968hIPQB955Q8LkYbqSES
LDZ5+tNZTF/8KTqGiNt8mQWXR4GwvRfMLMOMrdufk0nCEQYkzODJlHz3h+jtwsGnuEWezyDV8fk8
zIZ2s9YAkgvgvaqeL36qdb1P7/0u6WXvCAwEsvRewT6Rq75deFt4X6U/a89I2hZyQiTbjtN7KovI
XfP8811vJIpjmWrMS1itCF0qqAGMWtSZP2N+ZtqTZCKLmhGPOxnhgB5PE7ovF4WVmlAL9WdpuQfQ
AXSTKEZYDXjXse3OapAdlkwGo3UbaJUVl16r0LSP+D6Ej27aq/UmMN/71418kUqJnXwa4JBV1Zyq
v0YA5rgGaz8Nc6r/0yBd+HOzP2/gmW4sozDedUVGgMEsk4rMzY4kDjvAWw/XV9YGr0x+7x8CHKL4
RBd2IiZp4RF9uOmIa6o0GeZdEuhZlaoyDZuUgTJ9UPtrZ5TsdUgjYfBEnp4Cqw1FhTNsKAQgmYEP
KbtVcKJNYtIUwZ83JW0ORVw+Qit9BbJGaZg4LBDQSnVs7f6YUdm19lcq8Pg58Pkr5Gdn0N+rNXn3
a7Tk3rbxPg/NgKauyppmmCSEW8n67B2gZvW99Yc1WhUDAPIPD6qcF59ypoTc1BwzZtFZWzFxekPE
qcAz9kCh7iKUpTRaYKDNEhxfagBKRFDo6ibwO3QNrTemXHQhb9lsQCYZFBgvcInNNllN4BTDifkC
9GrwOq7ZrxxvVnbIaqiZaZuvWXK1QKXeY/MA4VPbh4jI9HiNbiHxRrvT+j2AJLkx/eUoyC9KmD3m
JM7h1Ad2q4woqbiSRJ2nSySVRn6x+sav5Y56KmCy65wtMGLCGvAPFrz812ly5hV/DHiwmYm6o8XG
yjVdHtL3Mz97hZnG718a60+rGsqO5CTwyUjTy+7WsFr3mWKW0OsqmUgks+0hCblrstiRF86Qm39O
ZO+F4qgPzpD58beEM3CMKwtedpe1colMfh0vY1tVQQxmEoh/N2w7MXGaMJkb8VNUZLVomQHh5aO0
7Qdz7tPQE9fUTnggbtevVhttqc0+JCcytQiL7VV0Y/aBDhGzgiMnWkySqbJysfmXn/ont67XauTo
NjqngDqsiF5/XBFcYPPLt2iadBS9g5/i9CHxuUNUhXPJlZbFCTQTWukDmJAipF+CtBV3P33LtMdt
pcxVeCOLKfuMtJSSZ8EfcDyqkhacaagoJDdd4bxQIi9ktlcgjIrVeXgwI8DhvvEUlMp5iG41OF2M
PgWdNVMXcjwDUDqTjQs59DwbLGreL8fTdjvXMJMBmju8w4clbCxXF74gh8pQDvCY5ZSYV/KcO1m0
c1M/8rx4ex6dWULIWnm3rMYWQuAn65QJ07eFgmzvOK1uyG/gXavSJdE+D+bhJSjM/Qv8W0gGenBx
IGoJNEDUzbe9DhAh0WufGX6SC7CyKYhzlpzHFZSQdGOIoYxDZzKnCqPUT5VLrvUX2RvKUqCGL0HC
S13NBo69HfMg8bBYLhrJE7zNYWD7OhaWWSK/mxM7qqqza/2S9Or9gFAMKtqwSknFlIluYcsB51Gg
hjrZ+jOIN5URWPB9q+WympxqBtUb60XLMq2nEvqgXAaze+jX75N14qDJ1WC0QYVFN2OWy7RHMnN8
TCICKOOu7cUW7IYkdcOZECUE8POF/yReK/ke1fHJ8+dfl4ULHiWNufz+v2mhQSakHzuyG8rkZ32W
ZgyeePM7ZC8I/5THtxSZMA71YpqRSmwcL6ZE8q7iSokpGQvrQRGltV/6uJnf6rVz350DMPXWmGZF
9I7R7Lunv6dBuSGPPaR01PyQAjXsWScYrjMJOgNcP9svP+W8xZILfxZsMJUZcR9hsDAXFTAXhPiC
wDesE9Sl5bSwZSukftsYZ48aa2UJbjGne7jIuhojScHwrvjCQlhVufVMdXE8wE+MISsr3T2TICtJ
Jc95AfGGiaFW2c9LbEXryrmpyqYK4fuzp9UWXWJev7zuySbO5O3hw4ZWl95dK7INCTHk8WpEaEl0
8WnvNHuy0e4ab6NxFovZXrr9z0remiHZAk2FKmDqVIcuLSLKPINuNddl236LyCrP2zZhy1Qs7W9o
Aetq2fmInnSjU7iUSC+9Nrr5ZgUMFClDJR/rHvUKWrkx7JRMaYJZ39BNv+s4lW7SUFVx+6aNrkuO
djw5990TPex9Z7Q7WpQGazEGC4T+LOC8+q96GL0askUWw18P8WbTE+HKMH5kj9Astov1CrZ2Un2f
wQrEjxFe2HE9829MMU7WCF2+ND0YRQN3za+X/vFXa38g2qqqqzII+Twhypg4IB+NHowFcgtgJtf3
z6HghV4h9xFRo9SHWCERtdFS0CJIyUuG1iLC5D91I2t/dwD5uDwgw80OXnH2nb16CjYcboBCjyZ8
ywtG3o2fneP7G1YS3EN56ihN3pZz4swRyHqe2ZDES/M9vnYjWqfoLTAvoI/akRTaENwW0kY+EN9C
EZ0WylIYYRIPMwtOnu3Tyd9KyW4Bu7pyUcjGAezDAsuFcj7kegFyNYbouqCfLhc6GIvvk9JkltNE
Lt5Nc4pajT0ccgK5NEvwGfAyoOj62UbNRN1eeKBCd/I0rZSLXaciT/5QEEFfHESnHY9YxRCQOpqV
Bjtkx6UdiOqw3Ym0EMcqazRyF7DDTBWKRr8ydMtsK7+86FMOBsV0a8B8OXnXOr92+/pzUHnmh6g6
luUqIETWw+s1hLKoBs7NMtSJF/1i+f8ZhbITtPNEibC9jyMse+bbQFp9MSZYSX9ThDhmBxOmfUmY
/VfrjpZ4HxJSK5NY5xTdDESCdYtyZgmFHiXDYJroEyCdniEzx63y7rDk7eJ/gDU9X6tbDjpu5js5
pXSHyk8D+Uhid5k+EXDEIZf7Zr9VgD98J+hzuOPnz9GgwWqKujBejur2Eg2egAunPAUadAw8FOGs
4c+GnbEE/QzllvI8JaVyMQ+0X5a3szd1DgR3s++FKfAdqHTZ8hyK0Gjw+xpEuv2YpIzXg7sWZ7ww
shpAg3NS0dPKY7qstYihb2rEPjAlU0n05R8x88+SsdTWAilfhhibJ2v95GlxqQXcwVwvpeCO+Hw7
Bci4C6vMRMPADOnJxiRq5+Dw9WXSQ6CTGMAo8awmOW6JL2V8Ixw1jaPpooyRrb/GeujhRgpV0VqV
HJ+NFQ2lDBm5K6uvcouPiFCl/bq1E1EI/xRspwVS+Je/W+h1oGkvui8bAbpG1plIE6ABaXSWEO7W
Ye36lGvyPzRrOr+gF8mg9nVisoTCWOBokZO7c7/s0ZDaVgcg8Vfj9P8iMRlxDFmA6ULgHohByZw2
IUk4Nt/FLj70zL+9YgtwOXJ0MueIbMY9AAeIPwRqMZKCpfl3zBcB+KEnBEBCE+jLi56lPf0QaLuD
PKguNjnrkRuy0EwxkbtAXIiwyt+KQZbAFq+U6CuWin2xaEJjUlc6BEhd/W2gk8aZfUw9n0WzdgsL
l++pCnuO4eisQ8bpMZMBiXJTGRq8BiH2//GHpAN+97DhWHNEAVo40xF9rL8njJllEs4WsF/d8hD3
WKtlZ4J8Rull+JYPbKjbSccB80nUQlee3fBZ3w2tQifYmUWA4UikQ1Z3uE4hf7tbCmduNFGL8czQ
zpYMH1Uf29BtlnU8XgOrlhqI4spHfOi1QHqmuMp9zGapWHTe2ciBtIiEYmwrjtVhIv2rzUNFbc4Z
6Gk7rkJIEo7Ff4PSwWbx7eMoAfGdrLqDlzWm/SEDcwuTChz3g0QshB24nRIxrGNC1BRAA4BII1n+
YHvjLs/wqV38ROJCYO1ASa3zCLkmK5T+oAYCDmC0U8wx1vBiqODVT+/ciPgixeDzAxWVPqffrhI5
GmSTO6JAyC2z1YGzqNmBTJy9R5+rTk1+BIeUsi8sswbVgcE48SnwwAZVr2RVVDg5rwzigOtVefru
xQXKKzBNChrB2/d45Hpka8cXQokBOAHznI1tBXeRD1B8oVAbsJyc7fr8AdTY2jz7ErQ9hPsruMpi
0wY5csSaIE6yqxYrjIXuXqsFVRq34ubXB+CAgbVuk8OKuX2Pag4ZMv+bturG6pN3jxppjM/9gq1Z
I3tj5XjZEcsLL1hFdG08Rh9l/yRIgXDfpAtNnmeuHlwnovs+ksPlI3fuPwqfMVPCIfP5TOrqgBB4
5xLuwXIJzrrsrh09MAzHF0Z1PeoFvCafo8SqJJPBv9ePgVhF4UMeeHFKh2be5QwDHrHRer5RlVNd
ResGtO3U/L/+MshTB4AomWaW3pRctEpflwlVTPGHILJgjjdoyH0Qq8lDN4e0gVbISqBxnQ/IY5D5
jv6i/fsSmJQa+QQiWtnIg9VNLMxpWjXkVPP9OvlvU7oxDqAbzQtlGsqFUVq7I00v0ESJ0cj3T/Cy
BgB04vCF2ceWa8+ZqV/6uueS4JzSQqDoXtAHeJvPrbo2NRpTLyz5bysX81M9keAUiDSq8cSp2324
vtNMT6PioKoc9uXD1d+ssWPW/cRddUjqY6wqlFGzAY23DTdcEtZBGP21G+f5Ip6d3oer0Y0M1DQP
fo4q4CQ7vK8NQkLNa7vZpzuzEEzret+TImr20vXMlB7MjB4bDT6WdD2vvvJRl5h61rKDc8Fqcp+x
XE6OU/C4kSQIQ8x0lXFNIqlX3cNAbOyZ3I40gM8CE+3t2yhtsg4KSl3tkp20rYl9e8ZyY+STIPAz
8z1G+CGs1rhdZWKZJbSs7H6+LIajP7tC3XxPEowi/E6tsxU7qj4uYHa/xWsdupAI3/G3LGjaF46m
WqP9pzCpL3ZMgCd8O06V/QVxcViOG+ShWV+i3mScAvayY4hMIgGSGxu2qU0hvqwM0iB/4d1cmFXd
RU6Jj7VAXg4ql/8JXpDqecVnAOhUPqUjiH+hz+nfllxPvJ+Ndj7IHiJ7eRNhZ3uiXACK04bynhFS
maiMG3D9Xxp27aL9Df6YmUK/HHLtBd88XNsGb73/Wfvy6d9Vo+Brasck0arPfeaoMYNMz706Iu39
nnVOArWIa8fMZeUyY0cWfugAELtQNYvVKs0msfnkpIacjTLJ4bWkEhB9RrrDfZrNruNO7hbFFxdY
clLz2XTotERaMVZEEx/V2zGLnYBhqr0AxoG/Ox4eQdGaIhYmbPtREPGKPnjXJPvrYsWg5z++14XB
G6PL/EBuAJnLsJ2oqQzLd8OajP4zWpKijXVD3L9BlnKKGvIc4fs3dxQDUqz3Ap4n3zmCJFlRGVHr
OuoBo9qSpVN+SdvT3HCU8SqQwnZFP5pvHiyu9gKRDRqsNEuLInYlBym8TFAjVOfL7Im138uvdXfb
665CeLxjCDNdA+L53/0W3GGG17Ym2khCYOIzetKtAk2gPYrmZN2/34PMDVV8TCao1PRzLrCwxv/T
AyRw2K9PpoVXSLtuBq5RVVuF1GiIvfuebuKvpwHspYGI+1jzj5WHpWmC3A5l0DPprDteoAqD1jGO
WvT57egYJ3lkrehW4RXxtfr5fF52kjUeqn0W821i16smWJdIyZEwWvQsunNiZzQJqol8jV6AUFMW
E9GXuacAmWcucfJiL/+RnYv6d8UQXO+Rg6h48xBeY7vK2DW3h12DWik6YoMiba5fd/gFhym853ek
0fj1i40YI7xsQFtKa8NWkH485GBWpbx9ce6P60Y/vQuXyswkkg5OtsqW2a2c8664u/pTlpsJ87pn
9Ap4Or1yrtc9ywSEVZkxQYN5otpUv6vLR+g4+GMVVmilZYHutHY54DS/sMueedZGzBv05/QQz31Y
0+pW108xMwzDfZR255nDl1gfcRPQX9G/SmlKoDu6U94y4jQiJtsbXyoZhAaB2gOjetVPk8W/JQyt
ZvQoz9vl+lIekTRxhmSIYaqb5mxTENs6TRbk4jNEqEUk5dc53qcQiPxF+sS18O0g4I856G3YFlju
ynxmepsunIiWQbqsUAbxtAetS8tTJb2Z4bFvTFs3LTRuaQMm33pZTta3mS+Z+YnwGqDnQJNYSve+
0t//ZxR/apU3RlsGCoGec2yu79K0O+teoUSq9ZLI276a0qiYC2qEehj67f9kgLq4OBqX6AEBQifG
5UMIUAOEMsMSMm0vQ9TEnnwNG0SHycK4ttSAnYcZ2S+GktC5beKJgp98DYlvi7DrMvcrpc0azdmd
4A8jvgMFqRzHoodqIT/GilkdIVPCLTTP3eVP0TSkNEYMuaqXhBIsps92vkpoJBXM8sbbdqAliG9V
se4YyoaQESfQyWGAc2GyGBTIlK8pPpnZwbgcn7UxMFShsyg66tCM2INVp2SBLuFul4qF/H8Xp2sx
8UhnvAbuhOcbqe33eq5TYvXzC0djVmpPveY3bPzj8Rw0sx2EvbhI4KVSelbrGUquQ2srR3oLuw90
ca+ctVgD2SBt1JeOkVwlVguamz8955x3sL4Jd+Zq+hg5VGAanWK7HW33GgF7COwkEOwSfjrIWaDd
difeDLMc9578dSjgAM+nyxncglUVVDFCsMV9Pp+9rfnaNl+PBsNDJ4c+3yTpG023Ip9cBDAwaB9/
Jt2d1kx5ZRtCj1xtTuXEnSYUvCPexpA6urXXJZt95mSarkPXkgXp7ojzVgxKs2JYNI7XiSv0UCEK
97/wfzEIm7n4lInr13CBALLGFS9H+Q8rgVSfxghVIaqgOzvq3s7lbDOgqgffDNny4GUmKphs9wmh
V+H/a+WOolwSTwdhBoneIMKIzMSJEHLzCYO1oOQS3T5ZZm1Bunufj4UnidUifHxNHNXz/TRmPygH
VM7uKucMsO6F/wvviHaXxbT0clDRNwbWSquIqYHr38XXE06eQMNSREjlhtnd6bjBlXPTg0CYQqNJ
xkC2Ar/XAEr1Ab9UUZMG/p6UNi12AjnRoMSTJEvLGMt3Uyl+jeI5n48mXkfD2ZQ4Gf4m1WmPE363
gg8bFWCroSo17en3BoJLqSGNrsCW1uY6Y+cHZindj8hduQbEnnfcRAAxp0vPbyMgKWLG6NW1xQKR
P21J5QLUSKqHHIAKJ++PkxAwohhE779L+/SpZ0RIzfNPMB8OZQokpOmnle14y66L3QErEOWqg5jf
hlboTDVZZEP4kNnBEexqcOgTSM9sb+eGNMZXJZyXX3jPKasbZzcr53f93QKNYcHrvLrFCNkB7DnP
5kQuP1ttNrySG1rx93SX5wHnXes2ZSMSshsgSVvGZWDuMeyURQSvHMDXAjSzWbrD69Th0q8jGYdc
Y6KrL1YxIJK/wBCIAFL/M/opwEcd9Zb4w3wSQmEc+QNS2LqHxmyts0JrBQssrfRf3IChDmXAbB/1
Ape2Dl9qbQha9lXoYkuBC4XxQRl26CCUfAgG8Um5F9uPdB+hv+vLWtXSaq/MTiPXtEQ3BasKzuUJ
NU1SWkayECjDNZhyQ2M8vB7dNs0bS0OJCe6xX3N382cUhKsNe5tzFjjFGqnqqrI3Q3b2MsvUWmPV
2ZbLZA6g42wt9dic25UUWasBjoiDY2kF1jnPGQVQn1uYwFdz4kxYY3Io6HFCj5YcGX9Tfjc+Nbid
uOzOcVif1S8mYTKjDCB3XXUSbtqmCiF+zYnZwcViM4GyzQZf0yp5uynRQFeNWdHfq3JwKGGf8gn9
hoVKQvsJJnbeOQMawawwpFuwCIz7WJM/9/yD/tCahTUskUUY9J1xRINYqwXIVKu0IjSvEA4xGTGK
/fZuYmhFRnMfrhRKY5mRVD6JVdTFViKFh862Slh7UP9fdZQPtsQB5sPASCsIkk2bPq2uczmCrqO9
BpMmksQrQCXZ1GdnFXrX8DS+LfLcxqNTYnwgAEFIAFMfVHkERoCWzGsEECZ/Wu4R6q5c8ESwzyaD
VCqRvyq9tmoBTt0zw2DLOwLpLJQLLFbmqinuzScFg44JJiSdWEPjMoNUiReQyBInujY5+tY6OjN9
j4WkF+6tqYutWEW5iZ8iJwJpGLs3R097WqZxFqPMFWjXBnJej3Q9Hiz37jLfUyWjcP+RJem3EUye
ZH7WT3Fy2HewXpBRvZDVUs5bDiwKlXAfiprL+u7m0TJio6SM/B01QxuqOe9XxUF+votNbT8TfoVz
8AT8tyZ88IAFgZCr2Sz8Poc4kIQ/gRVlyTk1/Cq81Rsn1d/LZhauytTMF4wzbLTllFWblld3E4JR
MZOEwIn2xHltX02xY59csD+9bY2GWnUQA2P1bxUkLpbPDQUWC2ChMLUx4weuJV21XZy70ApD3RrF
eUeHnPAonSliloyosPcKHFScypxJjg56mf0g+Dlal/0+BK7Z1zb/bTbLCQN4CVNnt/jH/C9KjjnV
+0hXGOpNEawyc/nHS3I86ypBZFNRpHxN9gy+L+u/L/hu488O/svEf+/D2P+HNPUyJLGMOGBIgYOO
ELXGBlnIJAFXZmX143cLUBZaZ+jIqWSuvoRvYv8dTtBRIBzxJEHWs2ge5s45cmmv2FTeauX2bl7b
fOoXUxR2Cp2zn6MvTQXiaDi0dKxpv8KXkz8avMUqC7MuX/28VFXqgTXxY8IPPZR0NUy6o6FNwFtm
bKML5F6rwELq0Z5b9LDZelHXGM94YY9tz4s0zcHgUQsY4/EW6Yb8cSX3tiuPMoOlWqgJr8UqxDfb
d/qUxzOfSCfH/pWT8722cmRO6lgpjwgbmpqd0oAFhkwJuRgnWHa/rurZTa89shEnKpmuE5/fl/dg
kBXSzvpO28hn9YQ7HqR9TVzLyX88iIzi9anRTFuodaeg5NtmWd8fmGFoXCTqU7OamjzEtQVCugls
ItjE7/lUEIQIc3DEN0WTcE66hKD+0GxhK3FqVs9wQuTeXJ6FM22zeC+GN03lV/gSmuT15FcEIMY5
UKBNkG+OPx9B5T1YblHuQiKA9gh/iTcnx4WVEXi9qBUlbibPeebuxBidMbkTI9pMRMM9WDraj2xN
u9/eMfWwLvvbVDKZt57jfdGYY6uU9S0TBtkakwGCAuPtC9Mq4DjgqvY3TAVh4G+LVk+p+d+ly7zX
hugtgFfYSMpsGQ3VFb8we74osebRx+PZpQeyZXeU1mmp0oHnQk9jU/MngehqHLuAaVF8p7v2yYfK
2Sb8bHDhE/Pj/EaOcT945nCJDzj9crK6e0Ue4tXT/tepoxmp/qMWwff2ECUV9TJuSO6VCnl81g4P
JMlMnnpNZhlZzwLfwocS1MyfNkyTrqWFOBadu70LXdz7Ahqv2t1lX8OLtY66XBpEuVVew/b6c5Bi
XB439oCextjDtilYk0LOHvlzcKIQFKPb0CVMOOla+Q7L+3XaGz6FXmJ8xnDkkn/5K1Jw/lf14JmW
PlEi7crGXtrEsS/u4m1fdno80BYXzC+W12ocJXaPz+lBsjSVoh+BA2mTc9OIstPAedd4g1tiXKo/
0I2tStbOLrkEHEsplg4yb2/jAiDuAPIoz3/0n08YFo+3gxZCvNMTA8YI4a6vC30AgMAAdb/gxqWg
S8qlgVYAVQBtnJU+Mko3uG4NMZo5QXRupKQMIhrWCz3hT7q9KGhAcUILP8g2FgYV2QyqkZiStoYn
23JojvdV7ZRt6g0cb0eMi69PROgGSqFsgcrK02dnvwCJNq1sK3znqMo922/mi4ddIPazGBCBpwJi
4o3v9uwitiyyNODa9OqdS23g96JMTQAnkGsP0IgLZ3Dfge/SApNPPfmrKqkFIkTkttFAM2sEvmtC
R+SK23jGfNvgHrWM8g6d1kY8qrCbvFgRrXLuIyj91PrnaxcR/xDdV3t2OHeOQdlswww6fEqKgHCW
hXGtfjCrZUvEYbxeojSHa03XjQeCAYW5SwtSAEsZCIDNVt32CO2wy/Rpn+fbIilUaLKU2pKr55Qb
n2XluLEMD8Bjrzy9K7CcgxjtHNqsn9fif2RSvT8CSfKSPj0EbBIfCBN5MsNFjjyo1NpI1aH+tBcn
q9oMHtIrp4WVvafjMlDxAAFt+IzdidMA40BSOL9zoPItFp2deWhpRudzVptR6iByXqK12HavPyEf
En4HmQLNVcjh5mmtM1HvP1oDeR5Z5JWWlUDryjtDRfmcUQ8zOhBrQCc8YFZ7SvcjAVancibLiViH
Bp8LTvcLC3dMzNSePhbnnclmypsyH2dOsXG3ON3d5U31J6d9iOFfasHUsu1+VM1H+9CuQ6ido6wu
Sg1NVzOBYdr1n3ZMM9UXzn1ePI6UKyKbhTN1DG3CbR5AsHlzu/pml+iPdc7lWWkUcjkBMeOGRiau
ASDlZyNEJLIMebkOfFKDi9PzRAoJSKDhNiLlOUcz8vic0Bx1AaBjUHt9Y6XGFeNnz9Wdn+ftpZ/L
1vK4hei2x1C08UKqKLywFn/8P7sYwQgOb7kk7ICVps+2o5DySCiF+qZsUt0lrGUmq48i+0TBprQC
gVV5rRVgxCx47QuBXjN1SzgSaoa3oF/PSfGUpIZ6ch2Q17SUDc7e5S5VBFxqBZtpmyqcBpe2NjPj
t7B2kiH8EfGAHSkjaOSqKyZtd+f8EKo/Tx/dfhOR8GWWxaJsF3yIWuNNUnhaUtbykTdds3P7oRLD
OkhMhzO1CkszHhF+djWqrYjqWE4VhHptJxRKC1n8PvpxDbv6wJ2nk0BbWBR3islLNDqr0e/zDi+o
xcctiJwW1/VyJXcgt1esHPBU3XRAVllaWegWr50zARWZYdfiWOHmm8p6KE+bRMJut1hTsVMEnH1w
IcpMBzHl8RZcXUj2BSCWjw4QvVjpVwK8LgpmESI+T6h0EI1dtiYFO5bi83kGiRm/ksk0eMp40nQn
qJMaRo70o+kQ0jDNEtDbtwJlxpPGPLa4xA5HaklW/pPGXI2mT2QKBWw+Xm/QLDhuRShLfGRmOT63
q0dbiZZMJtSTFgsSGt2rz4E9C1BRu60G374uh3j+dbDQEJlD50lw5+nh+CZ7aQQ/3A2rcSUTbgZo
3CA1PuJWNaRnHFdL17cUHGdDA0RTl6LWeiu+NBEVq4zMoJkESRrWKW5Tv4AOyl3Et4webkwMF2f2
cSNstLkG3R6UW/vxVypeZ4hwH4gfT1Zt6y/JkfTxGmcFSWEx8L1DrksFYe/r+jcRRKlQoxkz9wPc
wYRX7SKNKdNmK1khUM2XmfL9eP64SdOLqItZAJ47qeQ8vST/LyiFpqe/2aMRpch+nUpOegWadU+S
ek1Oyk1088FwXK/D3h+NCgUyoElMlXSqyCe/q5l4gR2cg8eNHbeHOdzA4aGSf3lwEVis9kaxMZ/n
O3gg+TgQp8nQfWeIPBvsDIXRADW7AzkudXzXQL6febCqArqqE3y3pnmoJDOixCNp9eiUOZaAFF/q
rkQcxJKx/sqS0J6no8Lu7t+Qwc+7g71qW2N1rzO+PelH+jcJa0uS9dCExSyvngNZ1tbFD7jNdZzl
faeva7NTbtyWoYtxbiyXgguMl48oow/FUo7vaXPfXayu1rQk3MQQh0igiBAVpzN22ubXPxwG67Ed
PWYcnam+uCSn8Kt4vMcCbff+R708Oxpc6jZWuaBYGgjQrkOPvzhnwe45m/yP2r6iHmQl6gxM3n5Y
+gbzscmGjzJcdgkBDgcK/56W+ID+TMRsg1OLOaRFXBz+xUliX5reCPEAP50tgsPqzXEU4zCtqDYp
uo1UDrq/FibzjkX8gf0A5JvORcbrWyy8Q8syj+nPJkRQ61MfErFaqRYVpbe44680K9wmW5O/EbbV
9XI1gfYldkSJimlNF5ZAVdg5X9NDEbMD5j/anVwNLZF8k20XHGwOghqd6Yf+iODgm4CoTezxNxpg
+a+aAyvh2EfR/D8lGauv8QN5h1ptGYuEYFuCVE6BeJgMVrPDEYignGBpyDJWXg0o6/21GjxZr7Iy
BtD9x5BCn1nQc4KORfJehkeR99wJ/KUpHOWWNhQtwk9V5EOBeZEzlOMPLgHOWuH+79LCDwfMiUGS
Pmhh/Q1jmqYivsAKZ39+kiagGmF5eV1IWIs1R2y9I2FHcgx1cAH0Oc+IjhsPsSn38aqTtnYbGd4F
ZDpyrWCQAOuKlIvhE9tLPc55qwrU70iDGtFLPJhRDtS2CdPLL8LljVGhBnsIfKrdjSkMVUAU+ryF
OK2EnwGxSkNBIlsraEDpFUvtdYpYtUF4ebfA5lcNbQA564W6az5dE3vDH9zjFadL7qOsjTH4FhSX
pHf3LiDISmx6tZ67Ts82KzkVj1UxBCjx2r8uilqdhmQpEhvwr+eO0dhNhP9eWnvbUAm2L/otpkcL
q53fTKo6Yb4OSHQTNxNt1EEdBWxIvNsKp+gESvdovZr5nFcmw65R2Q6bYvclnHrVkfJvpyH9p5t/
Kczbf6o6LyDdKXmhvHilpZy7luxpEY0/c3Wmffl4Pu2NVurjIhCoz2s8I0meEUSiF4+rCknBEGUj
Zz+LrKozyjb50hbHNqF5KPRpd3JWntx4NWPXJDwVOZjGxjAmi6bhJL4zlgmwVdSgyqQ6tRUGeKap
3giz57NEGpwbq5PFQhLaTpWjZttzRpo0ZkVQ05Eo/ytTe7W3iLs/8pFcIIWcZRAnHMTz/F6sc3SL
avUuqW7odu/mYTsZ3diq0vmy8c54Yf8eqEYZh2NGIT83Oy//rTXkk3BVvZ47+gS1ijK/8BH2AXiW
WSjuCMZSqwB326sIl6YKE8jSVjXEo7GnDGGXOSLOwkMi1o/kbhDnoxipNyLSh0ySLE2lcCEMIH39
mTRDXZUaHLlEQ9jp+Sh9nU8/K6r1WS1m1EpDbDadppjEYqDRrVGr6N2cz4X/LKekCIdBlquEHNq/
9rFRJO2fxTLSc/YOW4KBWPGVIjzvOitnpm9QOKyl+tLwWr74DZIkwBOmBc94BeTjM7mO9+jkY6j0
PHOTWxmO/S1dhEsz0/jY46sqyXf4/gxpU5fB+Otcws8SCPr9/eEgZKUy39JT1+aSGdd4nYBYY84N
gcPdrXBLqhivLgxb/4KbeyR5nqw6p+nouWZtGimBJS9B6v5nBz8iQClyRV9cEevmhBWji+2rpFm5
PdoW4XWDmDZOJtzngwPLrOCIsg2SGLr26yWy/G3eY6UaVPOnCtgeUR9WhXPpH89YkR2iCQWJ9cqu
m35rMoPNrGoZsj3Chosp5xe0H0/EFcwR1C9VdUlcLl+3v9YMqrSXuQYZ+a34gUDL0z4f0+/jY757
7rwXUTuasL7KKQcUI26YSmvEJdZbWCorfKswxO1OdJBpc59rw8HAOh35Jc1+PbGtuDmhxtt0Ljgi
GFVZXvsXxrm+MTIKvzkpvwSF5/NRavYsUlSIyv9L7xS/K6SSjAOmFgBJxACD706UHNeAvPvGh4hL
U7bNEvbgm6SwqB8Jn6h6cXLoNNRzZnFeX5U8FBptyw3fc98OqBXMpOSmDQh1i/hQhwO9eBbjVq88
hakp5T8PaNFuNGwrgn+sbXtZstuqqb+ycNtjkD44Gq0DujEglr8g/JLDnUGTsbj58OMoGX2g44vQ
A5mOteGoj146niRnTtqInnwUw5F/YW3ZQO01wxKPhOqnNV2GkI3gKxxQFpSeVsL3q0G/OXXul2bs
VMhJCjOT5aVOLTYT14MKAuqlZq5cFhD3/pO+3wf/jaQeQd34dRI6BiMIuiG+L7zsoQkadnIwXwRP
albPESb7WWJ3uzrO3egNLHx0Jq9MqKOPaThRgkYi+fpb9cVedUb2RtnQv4aZcu+LwTkxhzand+DT
vsXl1XBFAJ42JMwovVJ6bPhCsJKQnr4RHie/Ui3plavfJuhJrE2b3qik8Na+Fis4tvUxMCLStxoH
NLSFo/BBzorpZZXY+wPKboy8HD9i88yMJ/EhvE4NFnhWmaq0S8G27U/HgH8v6M6ExNdy25U0FPkP
DSL+1E6v9xgjoxXeuOuo4qMnRDQnHr9lpCxVw/kvcoeHnZTlOP4lrUZFw+gO0SmzVtDiNbDNUper
cR6GIOIBe8nJ5amsFBmhM5uyLa+wwGq9mRW27SRjllQVniFcJv9MJMiCMjGc370tCYGVY4oU9UFW
pF+To6dRnSCxy051lL8QPwzGS2JFAv/ZPjwET0QtZ7Pq+qZ+xbMRhcPQDnc0/rvonYSsxC4KrLOz
UcCOnuPOxqkNk2QqgjtXRAQ+S8trTlVqADQFGZpB1jPlaJnpWG7rP/42XFalXN6RCHty3bjP6Lsb
qShgNNvDTGYs7VSUIHFoqhbBT8Ac4+aKX2Y64SbNRTAwrYmgC4aK/EguW6cQaNfDZXeQbcxXsqqe
oA2LwG7kqkdPLBgw7VlmsHktfysmePXvMcB6ovPfBf/Mh+FIDn0AaOL95SOyKu59RxgzKsZP6qpG
zzHAqjdpYRhUgjSIMF7ERKyi79m36HqtDHiA6Y6PQvFYWwXc8kXapbovvUV/Qrw0E06BIlu1Fwns
jazTzzd+oOjKBreVaqMxabShtxVZRvwTm2y4JREpoW5+Qf+4hgfWc5HuFW3Fk73z7TmBs5ctus9t
C0t2FpQuIjv54hbOkmf5DcQyj685u60VMJPUGS01BBRWlK6V5wwtGTCDAVLptiJBPkDsSNT2IpTx
iNB23FDMpy1fkAI2NccUF2pNK7kDZ0zfKqPv5IGsuPxhjNpBXPpycD2yahZG1RUV3xtgSMm8aPQc
isS0GeVr7SQWBFRr+vuLYLM8UdAT19WhF9Rrz1eqRZaZiaLYhQp/9VCVsxlu7Kor/3G+OnBQcba2
occhLlnI7p2SzQnyBA0xf8zxH1GlmrR3I3dEjg8IaWNFZ4VAnO7cJKxdPHundHQXnSqngZf+mwef
cJ4vVnFC2EuLauVl3fwQY7BXOhqSRpJEIv3e88AO5e7337CyP7FrOUVtOX9ERQVg+yY0tI7oGaAC
537jbvYFxB6hRNOcWKApytZIFcgSIp7ys2Ivxa42A0UyomuSaDHKcDEuaU8oROOUTMoDr6EjcKCR
qUqb81BKxIipurDVza6JqlNcR8gZf5r3aRyWO/tmoJ1YQeFl+GpZYdnnejAexP+ph/iof319slyd
6uh441kEib0tQH854uKmxVkhqUMJQvoi102JOKRkSjHDLpppiuFYkrVJ+abIKXKrzyNhQlyC3BkQ
1llH19BSH7mS15pt/+T9emypM5fL/kf9sd3Fm16NfwLEW42vZjBgu6KVhxGoEsnnYTnSFMEWgMQh
m6N4KycZp2zHjf6xCDvb0tE8RDGr8HlyiGs4H7IQvZLD/Mlg3q528/yc3FZe1Id6eAIn97wSlsGX
y6SdxcYbpFu1jitrdmNPRlXJyJKhXQIVQjrfSxaBJHmYMJei5WZH5ki/dE8DRWdeFHDGeDNN1Fqr
4p2zAbv70IseG5RpFDRHo7Vt983d00XTtEtcj+loTUSfaoiWq1nc9hbwKrv4X8aVhzzU0/sV4HvP
iDORjTZy1406MypNDL60+vbASIieB1y6t+ylU50eBnnFxYpzeRxs/n6fw7kLzKJbgpXJk+8/afOU
WaV838O55T+v0wrlI86caHygkXSTo3ORoaIrN8RFwaD1DDSs00SWqrvtMkjfOMVBeNvIIP9JulEP
QZ8DWPtBtLGdqIBlq28pCnvfYPvJEgciwW8l2tkI8b06rcXPiqSnOrYBmbUwqGji6l4Tjg5Dcunu
AwDLem+d539d5FHPOeObcNCm/3HKbCA32+IJX6RfjJDV68AVIPHrx9G3zhCjZcOShybOOa+As5Bz
Fhd1JQPtj8qYw9iWRreuXGL1nez8z7mRy5WByvXb3ZRmnXpSeHV6emXuIfuA/PjvgNklUn4LUZ+r
gibwBv8IMBPsomaJl2GEZsjSKtIo+ulWfMC9Sb0kzpaJFJvoVCR5r6mp3DQHs47aFpww2lAV9ouP
NzGuaabyLqtnvlhp/10fxsbfrESI5318bs49E6LA0I4d9+VGmBlII8HSQsBOxnBum5njcJlHKFx0
UvSA7FvlSEJMYGOhPU25d2ax9O0PfnsKrZyyOfysVYRUPC+5fxJ6NV+xj4zRiNh7aTFyqOqIj/kP
nz0FQGqv0VjymWQ2gxEpHCS/dgvtmwcOQJSYJnlZ4ul6bwrSEcQLeQ1lk7JLRvI50Jbh1uECgw2N
8yikkdVOBUXpagBbCoaRdRMFwQD2+xu27RvULMS2WDQFwuJI1qgewhcqzlNJH3ibAmEZADBWp6uX
mlfOMOmu59qeLD21P/D8tILJPwpVhBNSpps0rumAbIZSBHcEcwjkbowKYf+AyY86/z4onzhjQzC2
8FPdTbNCpW0+pEnHO8cxm7GHpzEhB6eElVfAsKMPkX5kHHkr3iAntwPMyDbE5ALHKxwSLsCkVAWg
tpRvaHmINEKNTsHypnpWGXbn0tgv+xiP4PKGeaqTXE1j1AhIiHM/CyOcgQNfqpsfu1vVPpcTEKGU
iUErR2dplMzHzP81TtLhi6A2okf2EVQwPfc5FuSgn5MD92QzinxvExeoxnL7S1Bd/CMawV7eEsu5
3jDRpiGCLU/rFUP6H1uG3pRAsN53STUk122qA9t34Fxpor/2MP0KFSyBrlYxCL5Zj0wI7ggLvmnI
bQcWttCgY9W9Xc4xjTHawppaZZ9wmg9InnZsgiBM99KGlLcFIH1YGDEmzrpmXk1Tp5lxdclzKPze
PIAlSgW9MN+obcB2i/Bhif1EvpVW5pkxfKUxVk+YAsLvt6cmeKHu8VO08WQ3LlK8Hk6BA3o2K2/a
FcXKESa4IPpWf+1L0P1habrdUYyk108ugmVEJ7mtkwCwoA8oTvbpVAoejmDHubyLXgxhEDJfSyRs
rwJeCz423VsX3jCJ+XyoZgOqdHklEVCQNmS5cYfYbeOjmoZStIhi0V/8eczt2VNriL+zU8gAvkZg
/6xnLg14hX8bv+tFhkvEO9u6z4OL0ojepKK+LedMdPA+foVoorkOCu5nNIxU7rh08bO3ozJQhFBN
xVuaQI8T6XEXfttnRd4t8Y1j1/YxgYgBbhUWCQUQOBGEivXD1HgRHPhkF6fVpOuiq7x3SlGbDpqu
GyOytOTIEzTdHX4DaZuRpRAEo1jZYm1otZoZ4nwLLycJddk5RmBLc+0LxPn/iB2n9PYSFsEQQRCN
5hfmq+DKleJB8o/sQ4Uc2c+nKiqEvESY5W5vem8xH+na+cVj37sC35uAN1ZlcqDXvW6UlsjNbboa
DC8latueiQaa91OZUKD/7p68zPJzyYZGfjIeKwJCOsO6GZFTcs2UcOKx1j/V/TVa8VzVx0XhbuEv
7Wh2DA7j3QUDxRNcCItFNgn9RP0zJzZ896iBWPYNUe5GPlhJ4CWTW2U48UBNkCpKDT8cuAiQdP+1
qkaTI+9QKM/baFAunlgy/iedSBZv6IcRYJ3/7jBzN5CcKq4dh+nBiM+yH1HkguL4QBBrae20Gc4O
9vjOE327MkcU9BX3aiHvN/VgBZnPnYOl84DXT0YbRhDZ5WPhrPOg1YxFlqPE5CqmiAT+I995sm9O
/wS+NKkQebeYbBaeeKOFsLHYtCwS8PbMiNoCQSF9cPX4pkTbUyHZmMnq1F9So2qH/YlKQifHCARp
Sx7rcZ4MYRHKeqyc+iESd3NZzXSDTJsK6kOKhfnnpiAnbmK1sfQcq4cuLpGbeArOu4vwgrrgMbDu
bLkDlA/IVW6zn4oef4V/Rj55+rg6vbvLHhUTjsj5WPbntikHAbiIKENy0rgxH6OEdmMa/6e0y8ng
ku53UUi72NKHcNZFRWRIkovL/pp4lc16JFBjfuJxsIBQzhj1iWU1itLGofoO01/c0xf5Ch51JbjM
QjMrRiNU5unG7HFJtx8ILkdWIz1f6IURYwJiS/hs2PbE27VZgF1whjmbWFxgM1lfkXNZKryWensN
CmWV2HSOBDgSlifxNQNwQh1ovzGbXLwkWQ1C+1FZKc9Ucr2MQseD4dvOdsMiL30Lo+pGe+tgpb7T
kGWY9xXHtltB3gfFXDjtwpxrQUC/i5jMRP6Z1CrpLDVMy42KXGzrlr1RbGz8a4rgz+N9XhJAgymq
3mA+8QEU/X7yyRLa071FqGWI0a8F0z9ywEShymv8XakfyDCuwe8DHR5Wj7G268kik6xgqiUzoiLn
rCvO1UB9ZgM2w38y2BwvPkJQ0vQQQwtJ9NO1Rfk9n2EMirpiOspTqSbj+Z+w3vb6VLDQVjWB9Epj
nTWMIOWzZa85fFyxKftxKuqL3o6kPELovfDZXN2xk+iKmXRJ3TqVkIGhHuJkC57jios/aOFlHGGj
cycGuxLElJlhxs2Ui48NQrhKlqBYRIMhE4RbfTYMAlr3R1p9vofkeNsFyXpbGthg5wLuEIXbBO2u
iWommcfrqrGILJgSGvsYhmhBVcFiV4xwQ2LgsQpCbjdPsAFPLNMho5uibmTVt/QYjPTNHONlCnV4
6QGbF9wechw4crXINbYbt3TzgNSldMaBnHucWhTn9oP66atvwJJJ20o8UZhBTU+ZMAnzG3f1fyhL
AnzLJxYcS27dL6cIz12/4EDKQ3sw2xo8HVJsDlGMQ8pjqEE7ZaGx4Muwtg2hC0686AQwFB8Yl/KV
L9EhsHRlf2Gm/x9EP0NeBL7RKl/UMXGZoqG2tXOVrq3zd8FtW3zSWif+eP56zcQp8pxVHtc9RAt7
K1gR/hq+Veq4XHXXRIxeTOqYuDA8KsyLt1YOtY5AHPOnI2n2IYbGBYshvnwZDh5pwmr5aWdIamNP
GohdGoeom21iEPhaCJCR7uN+5PX9OVX02uyVMRzbbNEnYfq5gg2iCdnPMG91LIvW1l4/GOMGtHQp
cP0fGMGOF5aJtAd8yhJ688koIZl2nDBylx/JHP8wu2xc4PTs0AKmLXM0rtuAh1tlLVoixnvJoYtG
Sdc9A76DvV0qMZWJ2xAMhApaIAM0kyV84BJWkhItepMfG4zVHeadhZODglvC5jLIx4eWuZEcN4ZT
N+ixwZD81B0H2/E8KhiYxbJakdkg1mFTLIeSi/jmaGTCYha8WC8ICPqEM8xEZZ1DkVXYsur2Diuv
e9kAHYj4V4daiDdimGHTJ/syeWynCPKETCf3Y/h7n/vw69/CLEmj1DTzyjSCQoX8Ohsm3AhraCaU
v1zxTZ1pDHDOPbwYC1CxTvRvdzPaC4Vn4pkCsdrFhEu4I+2jn6acbRDYKvV82CBM6IuWMM/pQ83J
ArgZ5a8732VTGIpDd3Wmnm2MJR4+EZNKkVlf6/p4AX0q8GyMkmG0NksLPWYpRcFM2VeGrLdmire8
NKmpcZq3LFJD5Htu5mCWgvK3Byx5XWcnN4IMIi0VoZCtYQiIfTxbr3yVqx+APk9JvzGP2lZJJ3do
+brBqTJhmPL3VwMmwMjjWmeiNqOBZSXsOe+JozhnNEi0W3ULjtUyEVXA2SbjqtVHq1+JHeoqGFNB
1bgXmIyj9RshOAF73G7XblEa3bgXn3HPnQqYp1lceqTnk5L04scrTrBL2G52NeoabML0juFpUUod
MZMvp7mhGQKb+KT4lyYVZzlArgYM9sUmZRLpMXMiNE6Jo2v0NfROw0RcihxbdROeiqfLNszRRcgb
TPv/c5XHSNK+f8zF4h6zPi6e8Mx52VPmmaoXYFpRmBZJ9DMlfWrN+k5xptATnsO2L94bMrASWpBk
VIaFbYlG5pwpU77iuY58z9pMP3XPYZ8DWcbETSySjXHMkmUMgABx0ZvK8QF6jQnCONNZ5xEcF5qW
nDwfGGQecqW9ekYjBpImWWm/COxUe5+nCWib9wLH6/H5pD+eD9JtP+/wdjZQ7sp5bQDP3q03Spty
Xte/YCCU0LlS/Vmpvjz4oM8KQCYmOhptmaxwCKhjgC4r7u1n9twgIdYPgVFPNNrS0jQlJCzanbr7
y/V5pIkMG2aaeqADX/U0zyH/ZgJHMDHISbNRgtVWS4LRlpC2Hv5G8BjPmEF2wPbBT+4Azue6HigR
boeZCaeNZyCvSdDTF8uZsceVojSUZqgMeYpvytTYkwNsxtjYAnQsni1clMuykh8OITAghU6UoWrU
EJzxeYuvc0rLOrn00s9E9ai4o7kPBGF927LqDZVlxrcBYhEyJz08xe770jz0WnP4H0ZsEbThiIHn
S3OL21Ko/4GNp/0cMgHRwZPnwI5SOzKKFHhwuGbvhc8dGuZtXq346GCtQT2w9HSHP+AGSYIExcfF
98T37TC/ZaIDFFy4xeII6Nq54fo9f1iF3HR78ddWRb3FTtHNbzjQAZr2AyupbvOGjuOddNxQSXBh
Zk2JHmDVRMoVRQLJ978OQA+cgDbUZtMm7Qswf+TyxnB63jqPD5D4xC/egT1aUIUYLMwIBDkGMsCg
r/QWbRa7IJ07tJUc3aFc5zul6uhLFMSC+ZgrTRbkS+H/+OPZYIWbSh2WDDc6yxKM0qGgMtgtqYVM
zS/jk2d6xdhcyPzQYiVIBdYRINsjlx6gADOFg9310VCOxT9DHj/jnvzid9jGICGk0tymLIRWIt7Y
+GAp5Qpflx8R6L9bB/N76E3EC5wwt3+VIbqaXnmddsdBhSSmB/5iGYBkpkYEAIzj5un+xvio20HO
18ZurBBAnITP/qzLme6bKvsUeW8wc3VbPvCK51DpdF8kfJbx9bpLBdTge8vRpbaWMbI4uA7Tzmw0
f0N5/rQ5hGdxIXNglpJdiHSsD7WBZUfpIT1AfFDfxjsVsh4kRajqGo8JDvT7qS/QRkuUqARiyE60
BnRojYTwFluRK7rcdqGVZJrK2Dzt2Rvc7Q/zfS9w5iCamZCC9cU962Ld8OaJT641js2wpQX5h+Ji
K3giiQVLVmWCSchkiftM+vTYnWVf88ueusLUvnCTK0TfQwbhjXiRb54k6UEpZCfZGAVMf08on9r7
D/kCkBs1xQ/2oJSoW+Ckss+T4ogTK0M58yu1bEB4aUMHNXmxF/1YUdfLA2WlzOfGxNq36AFWmhz4
4aiQXIFs1yLhZw/ZNxhupx+3iaWIfnlinNIFCCRdl4xsyrGCLy2e26zf4ufICNhHzxwSBVFacJQh
3Px2bHg9Mcc7lIH9hG2shP2GY9XgNI6k1pg02eWEKsNLF8JFhfQTN/PKX/uEKVf8F15Dmo4xMZei
SQKLC6zuqWuq4SJmhrfUiazruPLbtnVnLKIn92MFhTds8dn7YqPKQgrFqbk1e/llcmz6l/SwDTrf
VrG9zll14Ae9skTRuSHtWsIt8ILSB/J+tEx1QBRm1eKM5a1KjwHlqJddf3w7yr5Zdtd21LbmvV04
0gIC3I2KQJ5V9EizfRXPjoqyjipbEUvcz24fxhXHLtjNcRCKcE6CabIFVw1h+QBF9OxdpaVNDVrp
jJ9Nl822tmH0Zm4uCihySDihleVLaGzKaod9eRAUVGmMJjiTzudqqHhTKr6QiuC/Wq5CMsEe3QjV
q4n7l0oARYunepfRBSQKMBTpGqCpzvSlnWO1zXYMtDr5yzl49GhAmo8Ot/awPJ5hZusYv6QBX4Bw
UQs18Yps3/o2mWoG6GR1DS+JA8Ly5KcNMIre9/Y3j4IFpQMamaNH/Dczvh97obJKt+rJOjAn4vnW
b1kXH8dwQJsRcWrGmzKfI+c3d64apUokNl8brTRF9LnAA3vBmeOBWDQ1FTe1IfdQAsvd6Qzigvtl
AYTpCiLWIix86v3nksgIxTGzeMO3clxHSJOv1GPGjqy1j2+wA5iD/gS622El1SjCELHkMYS6dt+k
4b/tilJMH/36JhV/r3nE77BpvPojVSIHy5BRBXKowvsj4ySapTVyO3UIbGHKO2nY+1hPt182dUYU
nPrQ4ulvCXCxnCbbyxN9LjrvS9QQLK6HPL7t9PLNHjoB00Y6XDKg2qN14h+Hu7F/ohbNDN+V40GV
TvA4Cr0LnGwtwtkhlViwt3R0di9ugR69TvNWI78zh38sRg7pjboOYp0HCS+BIvm1+AuIFGEg8d0N
OsqmK8bZvMhHBg3mAQGA1YwsB49GcMbD9sYgBmO7j/+GVrTn6RsiRG6u43eg+1gytI2T2hxRPVFo
Jy5kKU2eMKRfhb/pDsM4KtaMtlh4XeNrblaLZMHqrKUwYoQhGZcDEobfQ/soVI+jxUWDDtBMTTH1
UZ9gSd48Wb5JtY3QEqKu6OhxOgbN8dTAX0HzI56fgD6nYbmgV/yt6JDiNoD2b6VsmLdxbm0O15vs
BDCtpRm3D8hzr/Ex1hCk25EGm6In+jH54KjAemvV1OOXuTnhocDqngIqb5D3MdZ395t5vi4OUiA/
MFH56boS45GSw5LjNfQAzNtle3XTbE84hkM9NxVzvXQTiBqLuKLWuiHtZ2Y5HIJPV/8EJjXEHzly
WvorUgKer0dX27upJKFeshRCklmW2IDeIXqjAieWftogkruIVmG4VCvWfQnlwt6NGwfsLoJ3m+IJ
JBYB2/9Z10NYUjUTc9/rObSADDjlN4Zxl4ztN6Txc0dvIiqhuMZtXpUEkXwU7q1v20diMD4jtFUc
aly4Z/eDBCSrNXOmjswre/lWt/kaS7jaxnwdzwYFmYUTYypXm1F5FlnFBwS/hyCm5mIGLSDB80IR
22dmhzTBlG5I/VwS0NR3KlE5U5P2doC6OAO87xJwaEcsxYPcDg03t5WFPtfzow+izSgnSVRvtvPY
FQZ81YwfFtCtVOLfDxSVZl9ylab50Kk3YXM0CPpsETSzFxqI/YXBMX98hNcS9X4+Auo178lYrktn
wXqboKA9YxKODP1T4Y8UY/kQzy9/I9L/gvdA1Dc6AFowOgk3Cj1oNhekCUum6HZFmrQ2byh5n+4H
I18ArTnyB8sFzgtYI4Bd4T7HQmjOpNtTTmC7UxKRnw/428IEj7BLK02C415atByPg7aurzvYnDNM
Wo3PpQOMtn+ohxWeo7Pr5jqp6ChdpatbWfEHWJwplWiT+j1ZlvUsWFVrNfL+UgO7pC1JUBC1tklY
/I95WkbK9SzyP7jysCqkVpH2qRtPYrfuZFWpXfygU7o+A3nQDUa5s8fgN7tvOMZ9NLnabzE4vTI2
kZ96ZUch1nSw+Kv/hk5kS3w0fd1UpdL85hBUDf204wdGXJQnRphM9LmOOeUY7EUvrkQWC0h57Kqs
nOGszuy0/I6InuIsoWZaykiq1q5fipb+G67etGbY0knNtFo/kFOBk+juY9j1j+zOzJdUvDuW8YZW
OFlR9P0hqvjmDh8r4/CUwauPlQYiA8Glm0XstozP9wKxmLPda3NoI/H8T1T2ypLyYgAqscQYDPAs
uUNd07mY6LAKnizwsvaezZfGka1AdA6GiE+89ILtSfrgDQd85fhBQc4tU2+ttBlJmmfgzk+l8EON
iz79fYG+n4iB4Qut7cOQIGMtYQEn/Np/qRnOKzDwq54jAiDI5ZpdBTwNWH/a457NBTRtvYWtgZ4p
790HeADEUHMX46pDIvSvOCDB07BiL8qHAQyr593eVj6Cs+NtG0KyAX/r1m0Yfg4ISxDqkW58mtJl
SGoOG4Jl3P6UNTyZ1yzHbdp2joxEJEKSMkqjnFPHlHiJ1SLH7WfvwPYEJEwwPQyCPQG4AUytTetQ
x34kO9l1RKHGKSCjXEHiuuZksOngG6hDg4mhgCkCFLrBP7shIDdFHCgoYzOyYv0uorWfsdsog/Gv
BgOFKsILgfeceped21Zq26ZVMaYpMrvp+J5PStLNo8JGoaQUHSHuLzgTQ+W/qmP2XtI6ur7eBD2R
6DBtyTy/tJJ9cSU3lHDFNoTBzzophSokKBatldXhPduGcf8WzvjYbKvFVJj6KfRloDmEifkxWGRg
+wLIdmC1I8zVWHmVkfYLqd0kHGkurKEb3raXZvIXTcxA5jKXqlWACAE83Ba3ThJ9ejauFCtDrtG5
44VYjpU7fbVfz1RPV4AkYNVk3722iUhvlghkfLGgw46BOpUOcYv3POzM78JayVBNZiywuXE9XOfI
TvESqLRV5DuW9UpxqWYbUaQ9VdZHO14I+hJ3S04/Jw8DALDlvLtnfCrIZvISEcderUE5ldasSSGB
+FlAYmkL46py9DOew/p3/5nZYnTLHhTDPnAKhv1kluPEs4375E/qtqRwmeCaME8gwve9gPheunXz
OglW7LJZhblTG0TRd8bTqtXBF2lJnt7Jt1tVNC/7MBweJaiNcCuuwoV99RyWOzQydqXEImQaE9+r
B4kGdlMifGAUHtLGO0uIoua3qVfVd5ubS5O2HjuucJFptv3dEnXABgl4JGYwGRdZcWcUtiVU6ibW
m+dD0EZoxCljaT1VA1eLJFPsIBxPXWMb1V1iKjvdFIqqOFdYm9vWYA7Nkf+Lbd2a4gTVWQqd6GDb
38s2KrrYtpXr4vPBLOdhq1NPhqMop6P2lpGITiNz/I4OLEhUrdKQlnf6IXqEpPr2kx20whMbjvjD
/qXGsb6iP2EjNH+OI5sEKX6b+Lw0nPXCjUpeWKIE6OJ7O6tWFLYHDY2rL+AhL5cSgWbYVRcLmxvK
fDtszdWfBEHgfLnJ9vA4W6bq1tnmFm+5tQS+bjbTwzrhzH8/kjSFJLDn8C11EeWVfUA1mekHOPW1
iK1mIZcDkc4+0Fe+JL7ukymtBMDKLoaNEBR5lUe1PKcIy4dPUMthza44mmpeqQ+kOqpbZm1kyNo/
fQjLydDkOTOpYe7BnPaPM2LbaTIbkHHcXy7dhVcfmAkUwrdMlNZS3BhOqmhBzWFomfRmfsbYUf1i
1qvU+1YEvDbh86lle2nehZS4Pzo8nbcwQgaixOHoq3aNarIWJ1LyndwPS5ciQ+t5CBtse00Yeplv
/KAF3ikfy/oNeheaTB9B+9468Z6og9YwuFYwTaOheA8VrG8iIse8rxP3FRDDz5ndUzDku1cBzAeS
NKM5qOlQx/U4sYp43LfAON1B+bUfasfUfaFJ4rQoEsn+okKj9v9M053wcvyTdOVp3YAU3FO4jRoR
jVnW5GYq34218oQQ9iqTizWgdea/b6C/nBiholZ/UybJaiFwrdX5B4SfaMlw/+nuVcPP2qWlXq6n
VYq0WWpkFBay2rJ7beoxjiQ1gHb67XsH3d0U/iS2gcwxuF0M9/U4TaYqDaA3om9SY4KHAfBat/Lc
jwci+nXTecpAbn6Fj81UuwwnVfKvS0NWluSqAhRl9zdIeettazui/5MTsz9WK7GQpJvNJHN8Ng/u
csXUnbF4qzx8GjOaxgO6D9mwPJCpmAyFU9dlQKsHlmEzDjP2pQqAvzdZen8MpuiIN8cnh2SCoKcc
+EjlFIfJvNeIxzbTQxUw0wQi7HIx6W3GtSHopfY3ICnJpiwt6hMEXNfGfmy1mKWGknqTCgqS09Go
2G4PKD0A2fKY8El3g2sbWK4vgMon1/C0nN/Yl8yW/q8148HiISIutO9BPbwYrDHQOseqsLHTq4oB
z0S3lcEqZAx8URbj33rAmwDUqX7Gm0t34X0CIuNGHHiMyVNlm2U9dVwtWgyrUxhnrvej3FViDXho
JuRMkUaSHP0W3CyRiJhgl/Ze0n1pxf8CzrzemGFQ1OEYKZXFAKywU1QJKsFONDaE/t+QFr/E1uM9
jRz6Tnznen3BwWa5hepi3cq/EvmsUH1WP9fsCipIajxaNnHl8dQppyY/Le+z4+kEIEQt4DbRpkra
MT8AEB7jseHH9tWeCOClPL/1kF8Sicr0QqlPvaD/3GS/mCP99lkbLSMeE7GwNqK/IJjBzVso+ucK
5zjehAVieUIQVIUy/oKWmJcpnRh1T9TStN6MZssZm98tsBsz5hxBwRnjB2bwKtVqcggWIxCggYft
3yDS5FVTUxXhtRzHVWvhhAzSWJ4W2VvM2O74cSeYmGsyt8h/qLzEvn0n+ivZCJJgMRf30AoM59YP
ndorjVgDFkQI4bl9sNUYYLcfPaBGaqNAmqVJHyO+CB018okwiW1JJLZ24bV72gTfIkgXV8vts/ds
K4nPPP8Fity2OiVxNsNPtJ0HBXpQX6SBmtTkECm49z3vq/DaAkCg0RiUx53LTXbyDXgiMA/N5YX0
qp5BTvb1FvSB2qWwNQTKpZTkwA/jWlepaewfWoY8CGwX/YFOEjnopITH3hzyIMgj/kQduPhEEeig
xPC7OGKdquWeWffnZkIIissNi7xABmf4UjpNeyH2nUa27TkbsoPhMShoI3qh/nJPj6LPY2ATVQES
o4ZNBUT9FebIIQ3Fh9He5LwX9R5OuVT5jAnLuCj5D2Th2CHrFlrPnIPFR5RlEleWmy5Q7XtU0gxJ
KfEzHdrUYiCvWUTPguAM/Z7DrwLggkMxfTo0N/hH1m9ChNZI4kQ3yveJXT+LPCOF/2Q9HrESdv1Z
XBEA9NFZ9WI/0kf4l8K9A0tjnK5SISEgeGojpgNRX+FyGiQueJgS6bCDJ0c+1HQ8DZW14QN/hIpa
aPO8taoRE6iZLhiEO4AftQf9/bzvrIDN69rPOjM04uMo0jEb9YKi22xdcF4aNI1NaG6LkWDZvBMk
OBdws614AME3r0h54i3mhxwbOX8637akLNVFhJWEQ/SOnlWaq5opft9tRs86pW0oy4I9DBayFVnj
ORj3QpgZrIGNJWepnZcVRJq4dNTK4VOqfrRIkq4m6IozAH6Qt6tHFaSNk347rjwwPVV+4w7r1vmP
rH6Q7y8IT2QcSnsXrhMozy6w2I1PzmFJoALCTROgYJVTtRypSgHDbOsu0AGBGToz3wRWK3fn7U2g
tgP5SOwKQChXm6AMu5Qqbsb4q01Sb9qEau7NJgS0gjZLOuxz5KwxRZ1rr5j4q4GDUPwRf55eVq6f
OtRCH90BrAx99AsxUuFA96qRDCiVU+pMmF5REajZhKsEVSXQj4zNptMiPllMZ72edzJr5LPz4Bdj
B0+p5741dJ7BqqaSNl1nlrADp4IL7pEEWLxIz7ZsEv1SZt/DBZrNVMyaKbHM8OcWhNO62rIb7ZCt
viiP+sqgSqIkwGAwp70fUHMGX/q/DoH91YgZYQtCf0f18WYjPw+RUXoPfUsuRDZZW/cPcBcxKehR
1Vv/G/22xvGS0FoB9HWVKG4T8bU7V1z2HIDzIf2feqev1+koqumbzy7gWPemwF7qrAgKg+u1YPVJ
BLW5tfX9yrs5B2VjwRxegEnyPK9Tcxd++ZY2BvX66+EnIt7IyFqyp8vonMl/8P/F+6YYRmxr4kFS
9L5jTFY3NlRBSOlXMIEuqI1JTXbuD1IYq+4C7cZim1VDmtX3owa6FfhT46qPxRhyJKD31xPE+0GW
uHt3JX30UioVPk00qLD9AF6FOSns+P82ayswjYgrRP4ZqaxkuB2IQDGbDEi+B5WOI3ulubEJhqFy
gWRU7w/sXKsCrdwuxouVainOXgFXZVH1PZbxHawCQu/4f3UlvQVrSCe6uUDgCA3q6yFlJ0CLECub
MV7R0FFpV+t0fJDDrcudu1iMCFMCX/zOHTyuBe5jYs9qXpF/jjA1qOoh0XKPP3qtNIyjlsJG7Mcz
NtPmu50PDzl6f4h+10PRTjU22vAg5zdXA4jSGDSt3TOBqYlbPHJd6b2wuHXZ1tt4eOOxQyt0ZN61
w4MuLqdTqonBuFy+J2rEzzkkUIqq4F18tBLNkFzNVZkgGl+zs++7MO3M3Nzin23XuV0bSMqjmNDQ
P6+br/WmQCSmsmOaicuYx0CX4zNgLeHI7Ls+zHV6nFUulDaVAD/xqJBB3Q2s5bA714vTSaZkkbhY
GtirWCqIe/sszB/fX/UbiUrH9mLXc7Wu3uMf/mP8BYM9yZV15Ea/xS9Xr3WNaIiemLLkh9MYyVSB
f8C4w8g1GfEIma7Stv2gVGf+fbNEeIqkbSVNZd+Zf50PRjB5YQzqHwKOLFqcjDoiQpXT2MDW87sl
OPcoZzFcj+pkzN2/PD6UKSv6xXWtDe9DVnTOaf2O5BsyuGjs26uyYJExKJsSoMH0SvuWGbZdVVWn
vFjV3ODj4gnJwUlmUaNPs7967Or9P+IxqKFfVYUZ2KCmJkSJUDn8Sbz95SjDt0V1eqeY3n2ttfnv
Fzfw28TeK2BQIimRUbGWyQQoBHWV3AjD6voDiJIGB71kniOv79wfnBKXLLlHusUTDkLS/4qd6ovB
FOsW5/0e58DG8wbqdOSWvQiv76YrSmj4tDqLfNl2PZNEI3iBOCkmppjjt1YIiqRlQJWw/qI5LrRL
LSKBB3EN5E8jPfQODK1DvwaB+i7J0DPPIFro0tK+ZswnKVNFtZe47tYboG89HMykJ++WDeKmZGcn
WeYygVp7b2rMxrgAWj2B2C9aITfeiulrMHBMKFs/RKLPtipYO2mT106ZzJav4WgutU6MHxwYFe0N
nPM2cKyg9nRfqDaF6RxmvY54nB4xnEcujwIu7UvLijrQHTanm1XsPi9KXiejiJulxwL2iYlrNGyw
l/jDqnQtQLPm7Es91u85jUd6nApzb8Z8h/O3E3WA5XzrXYVyG0IZhlXs7O9nLTm5d4YeWgm8uzbH
Tab2fO4ndzSFk6pibkfaevIDrgwy2tH341tVZzjtPpo1bRVkbKxBgiPPmxNkvWaI+3cohQ1zsYcA
nHDULAH8bWiIApyX0H5N5aXRjVA358lxhejANiTsv7eFSHtJQ8w1weCxPvMLduNWhmMQQKiaZv6s
RKC9xsBdrZYiYcaAknccUq+nC8nFGRwlTjzOjWkZUNR+IZjQQ/kf2MXX/pvmZHNYxDtqanoaN8UP
xUjzPRWiOJNGgrBduZt5TkwvCSK6T0Vrnc1girypOc/pRWPnFCfXR2DW3X2HUUPof7tuQE8oPi7i
1v+6KAygPN7yeUgnIrWAdC5+VJr/y7MK2Z1dk+uWRhamAPzEwcGeugfTNPdkk9Bo2ph/iB4qgaw6
4o10QnBNTtPVoRfav0O6oGvFKnoB4Ef/W2zpB3b4603DVAzNw3nIoD4KccLztyH2rhd/VAttmJKH
XiilmIZhHz2f5zELFKfQ8pHtWovrglFPmw7fb9BpGy08bSjSllAu4zC4+pjmYR6D5R7XyETU4bz7
1DCVfNzZ8wftzSk0S+UEC4yzoz6biqXbCHJozcrnN6A+U4xHF6ins2BGxEUsC31auu9sIe+D2+dP
h3DlATwwlg6AxRWCxEBEeFU1zm6nkgzkDEo44ieUdkNcRuhmxtB8fZXoJz6PSEjEzeETVzZ0CVm0
daFUSLqRpwsTNfuB92d+IU/7kdvKnxgXexahQZmB1Nx8ETpCPsWHxvif/0HeRWQ5fmrpQ3w2oOcy
vxsZctFq2W0AGE6G9RanASfyAu6rb+9SzLap2pieHh6GZVOrlbCg0bnBi0uG8TJzgwdyTaN/FLv+
yM/nNYNpVpmq/mGZWDLlpsrFjtBCJ3O5raIWgFW/JIuEN7LIqui60tpJU4zykprHm6X3+JdYRyRR
EbppD/z+XAKg8lckML1c8r5KIV/ME23xC3M2vQ+36C19QYO+0+lGBCR7pINDlN2JrbOzgUsuTlH2
6y2+YlH974ua33Yzo2WkY0QS8JRO1n6cn6BIx9zEcbAVckXIE9QvZ3ADiLiiv6IySQsPESVYpbqf
pGbmo1CgIkFLur1p9weVY9Wp7Bi5NzT370QOJwcpNirBCcgq1cz1tyhP2W5VZ5i2d9wqc+D9VpIv
PSdhBABuHx/ugvnUq3eemfA9+A+C5VxfGncELWfuoXoiMFb1janPqu3Gv9EKB8RfduC0h0lsa8EE
T5f5spsgLTDydjjcLAbitZ5Hd60OKQTIFbckvmUxU1y51g02h6cGMDT9yIYEPtv3BSlmicZejv+p
UBRa9lPIfALrgSrab+uTk2eLRDtAjTCkeNO0giHav1zOcx055ZNDRLSJHnghAOCIYcUK+adrAirc
58cSjLDJm7bqWIXvjg1S9zim1PvGHg+bG1CatTm9sax4USnuGQ5115tZiaetaMvhVzyLcAMzx97C
iVUuxaVJHZ4BDAuh0JC3tQwW0iQZz4FtCjJt6hTndo6FcL+Esmz8uMzeuan5X2i3xlGxXebTIG7S
zY/ZgMc/CpsMLXzeL5YcTYovlx4bcYjGzLFa0JZayHqlyj4dQ2x9xyDni2c6DjLUawEJ1AujQ1Mr
iDcAJFuiFLEfz8uvTLrmUrIoYW6svC5kCgk2Y7C/NZBGDNIbAejVVg76r2tzlWJ00mwmTcYaxUth
owlNUpfgqnl6wgMKJrBDQ0E3iVq/Q23GrcebaVWHYntX0geVjCUrNlu1/t5oaPQwwMmg6DUafa/q
E9qW0a07M3aPgntsnMBwQZfUYUrrhtSEOdho0RCQxHWtMPsoItRGhwPAbfQV7ewSk4/p4DUNKd8c
i3J104aFJE7PRSPf2Ggj+FfTMQpkEJOno3z6AU1BHsYEEDygu9S2wnxPt4e2r8zADdFiPLpKMnNW
U/nxmI+82ftlfp93S2X7N2B2ip/xboevlmKBwr+h5B1iA/VXvcw532doz9x368M+jz05J2EeIrSW
c/KJPoV4RF/hDOMhFJYv0GVGo5oj4nEm1Q0PmndqBi3iPSuE1pNLbRo3ypCuokl36iUm8W36OTlo
F1BQINqdJDxSBCfVVsjIYIs2vjg95R1EJ9pWD/zow45AoKpbB4DIgmeDWWS30dJbfdc6PH7iU74K
hmhXKyLtwwjPQCLcwcRZr3jGqshj1auu4iAJY7BaDROKMXTvI8YfFvUFrHMF7+JmOuibgdR24mH+
eWPZzFACt+r6dV06KtlbyY6CqRCRbxb2zyBHYf9imYZkwFylngl/FeZXDXoG3dKVIEfCIuk0YCuP
nBMILeMtMN04tCeaep+6jwxQv1rOBsmepk8/CLYi5nvf6N+hK19NJsBj/o0uiZG5Pw+sR2MTWxSa
Zi/5lrMCFwQwGAGhlqbXXVRxTfdNNVZ1eMwKZzG9BwHEUHcmizJTG+t7gAdO6mD86zosEPLrJTO2
kI56Qi2VEDXGLu0hm35UNCzZ+nMtPwWqj/LS+fPhERz5BOPCo7Xk5T9G29WcjqXqVMmrDJ/EX3fu
5KFy8RbWarZ8EQoTott38HULjGSM/TyIoQeEEb5Md8j8cqwH5w23dJ/PCkO5UUnxg/qTjYRrIAUD
Qzj6ahR/ddwH5dED1kwfvHl/uXx8JGdknPULwuW5kPolYQg0nhW2E5JIKLfdrVsh1aslaemvVaAJ
dmI7iMs3qgv80adbwfYYkbbdFG7u3c6lXqJeSgKwZBLek7ZMO1Jpi8nAJaLcYR36YmTIbftD6CX2
UT1ZqziZbC+NCey5pCvUxnjRekP6dzo7QZHZ/JAqLcy05b0BeIu6EnGY1nbSF0kepNL/aT5CwQgB
UEz9W+9eRWSFv2FflPL2ennhKpGsJqE9YfZjTfYNIg+yE3JllvzPT3YGLUfEyslIiqc2wOMTxex8
qN2B2V5OqVid+HZDb8G2cYX3ePaur68fYhDDYZ0NV5zakySIhkjLIHD5uEBXcTrTZ8RIzxQ0we6H
+uBT1zBDp8TGHJQE93jw2WZYQyfDM5stJZ4RoCPSbwYiMd8+kNcU5nbx+zKfX+ZG1MgrhIPIPWA7
m6j6AHcOsRZ1UpAnLYDJz7Wf+OdhqxsYYMcTTW38neeoe+96RPLIAf8TaPVEj9Iu5adhxqYWJsfM
o1a+cVTsT6oYOEoE8qS2DSYAZJJswvg3NzaKuUf+rBQrdTfcIeV9DZNz/91+HrZgVgrpzgsnfrF6
P2ZbfueJsUKwsobBetJ2I/IH0EKYskzQwf9XMrkveGUw87/hpPnCmuZ6btCDoj22WpL/Jw3eY1Dy
Z/nCgfAr/RY5Itgj+9Q0Xlrog77BY0Od4HzGI7baZbHgagBRJ+viUY4ldonUdMNgYqq0nG0ELZ0l
dzh/OwY4PIydbLeFURNbDDQtLyRbqiFpYJ0Y8J544h0C/iShYDiCmcND0liO0WPsKXGJpWpgJCEv
OtLnO0Sh9B46tIl/qdJRMunSUPQbcI+/e7i6nmCKLSh59od/Yk7UnXjj3b2d0dVyZmg482FSGof/
SqZaBpWuZE8gMfdYL82oHoxuym8HZihPNqsAX2/tf4ZCBssDFwALTpkDen6m85VmTXNMJV+ro52k
+kxi/ethKei12bjOs7vaewp1BkD3BmU0fyqHODteh9OHY9A5xWyGSBQGIq81SOUj8VLNQ3/bMlY7
8twL4Bw4JHUhXYzSH6BK9ljZyj2RtC4sORL4uv1byTTFhNRYVOpWFwizXXZLGCrpU5BcwGMEtX0z
MHHqWzEC4G9fhg7y7mT4nfr6k+UPMVlaYQySLF26AsuOLmZL+06BRBPvQYQPabJIGOItb7u2ocXl
0E74P3H08aPxIcO9A2rRGABpW5y+5dVH++u2SeoO53aSQllsDIqKoS5rPXNtymr9lARgulO2Xl8v
+i9b9YDhNqpmr/VBN5SkRdLBxWL8X4dPzztzV6MKS/ZA8DomqXaba6lmKCfgny11PMwEAKBlZmy9
yLelzltZ3n3XjySbHf5zL88l6KA9lnY0aAUu4XtR/jSq0DvW8FDoLKGrzqf3R2zHegco2tr7mWSK
8NvaQvwbtkdVi/XQRd7LHX+XroSuTUwGDJUqvwHfsHxZPFNNSmSttga6utxAm9cBNXD77/ORH4xl
bAqNWqi+UQ/ubu/SJe/kKExcAfYHZXaKgJEgR4mWdckxjwy2lcJs86vItDRYXZaApz3h+NWg2zzv
if6QKgAFkblsS2WGtr4glrslZjiEKvIhfPqHoSJo8ZyE36viTo7mDzJk4ENRVPzBhYuM8i0yZAc3
+r+3sx0FSUx1OdsNbslmcY+ANp37aSopTix2tGtKrIs2dUIsjQ22XnSwA8bCpi66lagRM2S7lyps
IUSM+5ADNC7sL7cR5hp+lANTCgeixqG5Rl1QQSRcmGp0sqWHN2R6rNiNE/VHbtIAg4FwhOeHSncI
622gErLUNmVSkLLiVveiI2UPr/6+hSp78BCzRKs3cnXdNRfM4H/pXf2wXkqT0wsOiEnlin5wEFVN
IHgwBrhqHBc0j45c9GBYYtPFSOFuBuo9g7P5ejEEoQTnRF9j1ts7HImJm7bUDhEY9Iyif0SGJq89
pOaglFijxSQhZ8qs6zAnBdx+8tfVDOZWyCZEKOT1/fR5QmYmzqgt4EPeT6YUk2leDII7173t/Yt3
ClpHtvN03KpWCxp+cUf6WcjWcYV6pQLuHuOD66uvzx21252ytBSh3bD0HF0ELp9d+ZfZFdVUFUvh
vG9fLYDdkswX1UjmdYSOIB7t2SXYSD4LLBJI7Tn2to2n+40hAVcEkTjACSk61qCRz+k7kOAyxYZq
HPakIPAhpkT9rTF6GKKnZCaMUvc3qVWuP4w35fBDEqNT8qSZMc+ResVEVbUkZA+JIzeJs5ZhuuPW
bq42m621+kL09DzWSOJSY4y2olN+j3VcmpbSZLQT8VyWLHghhI/4XiAtq+l7h+PGJgPAT/LSBhZE
PUYUaH5+g/CKpJ3VKtKwop3xH9vaCBM/c4gszt7DOAk92tRac8973SL0XEzstjpf+wqd+qoTr0Gl
isUnS/h9HW+twAYE4HntsmrvAdHZl++jYwtAmxCvyoksiH4vpj/l9+ryW6XC0mAh8xcJJRWFufLb
SiIr8Vrq2ioReFY82FI3tZ1PH/HrfLjqMy04cSZv7+FKbabFGcuVI9zYEY6nJK44E+I/wt34JunH
QLx8boDhWnla6XrVBYGggqUClsaEqpf2Ed598Jzv5BOPI2SdKAGKThsp4Sb4yrtOnioS6yuiCgH7
BXEBIl8dJQFB8KmO9duleMyrt3bC82rpwRwEyJqGk/MUohRJt3r5YjjLRlyQFho6fD1alUOmJSgy
dGkOkoBgxJbTIpf5C2oxMFzbaKSpLSR/wTC8Ce4q2uOw5+BOzz4rVO1ea3lP3n8sxg7N4wBqgBPA
l/IoxUNH4RbgezKAnysaCNMfIaPrE65pmQe72kgdiOykV0+59yR6VFnezQzFW9N+GYz/QMl1UmeK
sXqnWn1LTVXe9FXLr009ZXklya+hNqR/sZFcx8sOEgHnYhwfh5vHSdNlX7UqQgIdQ2u0VSBtALWC
NSInxZfUGJFBDE2VcGPftnjLPufX9Q7QZypsqOhwj8WmMxuVrIH632onyPpcZuGbVlaDv9lDeZf4
fs3krGcxnXUFIknslb3elhS6w3AOAuDF1WzMdz2oB7vCv9VvSp1QZb/gLiGcC8U/dFpPMwv22ib0
q0bSWYV5uBiG4hyxgsn7Vz/IgY+IhdlqV5/9sRm9AR/DDkVrPM0PxSV1JFyHGTEpkaB8M+9NJm3U
iMtumtKoTvOZYFYCSxOaypubm50zXEZAf1bKRMll27QAv3QD3F4Rbs1h1YPTzCwmoJi9LXoY4s4q
/4Ia3BkCo0nbyO2xbFbh3ZLZNwmoQrLZcSEZFOGEQzyaT+AmxqhUF2px5y15JaVuwC5pkoJ2MOIO
316MwZxjfRmJN0ACVVRFOYye3IvDHRXwUtKmVC3s/uJouwuF9XtuVQO11TErwKK385EGo2HipDPm
Psr4am1mCHQ9lDiey8lmXx4Ft4qUmH6hmDwsePwsiwaDa8TGwek0lZtkVrZkFsRyFSfHPHXI05k4
A8RgYxDubvjxGJtvPNIa9Db+sI6f+PdRnOl5FzOd8smRMzsgUkJh4Fxj1XfMefrlLLOPAHqUqVLF
zOLdSeAwS+W+MiGNruKHJeyqXgEMPzr9Q9UEj76kSc6v77ec/ocxAcQP+QhCDDRk7M2lIERmyfzu
claGywHZmoC3xcpcDAndW09sh0+Cg/l2Vmu4UbiNJ5ikQLQEUUnRykIgBf8lHtkmfusCKf0MXTFh
Rn+UzGXMMAByxhf0inCrqszaNrcFbURf/mhOxn4cyDID2YCgmXXt70QbSRKXEk7HYbQSP+2kN5bk
l4aBjbdPFuu5YChVFdTU8RCMgN7toC/qJXgEgMFB4tCS+IhzuJhVorpHEJ5KQf31+90nLkaZoJUk
WWFVWBDsXIaqojr3PUzDpkzCe/cCfZfPVRmtAfyZgHGIj16HdIPyvctSU8q27MauF70/2FUn5px4
bSiB9sQ3/QGC3COuYJTT4VRqo/GANRuEBts70X0tdnKMAaySQ12bGwtI8BRjcI7O/AMmQxVA5AFR
oAyBnNsnySX50MlX3xW2eC2mqzigyYfpRuJj2tHhZE2lgHExnImS3GucOvV1d0iCMyacL6qWeLSW
c7FfoeYtTP52p/8o4UqKYJv43EsQHj8VIrXA6g39bowwn4/hkSmAjk5+LgSpWdD6CXG2M4IaP7Nj
qEb/OCbGkgBYh5AsOTK89hiU9xdGMhIkyA9e+ZHvYMALddgtYrmJPH+Itxt3t/xhSD+GrNeHAWQW
MelhV8178HUd94/SP//6e/7R89BHxjHrKMRFWcO5ApYkMeWMbwlRzSEY8Pkj2ih4zE+lhWSWdNwU
kEhXF89pMR4PDp3c3C+/uNuW/ik0rLDAnfFA8clsYvxaphmrXusMbmY0uj9zqHYEbnWL0DRaYAC3
93wPXlivOhKHPxVWoeATNl5mrLh4HO0qB1zGqYvlSh0hkBObc4D2j47Fd/15AY7VnoPcLzCidJg0
eK9HLNOn+DcZYaDUDhcLEsMx5iguI4X0o3nScXh5WmtUW+U6gaTNgrEInVuIyK558FwB6zLAwI3S
a9rLP6cqNyt7ySZI+/ukdDBdGE2V/MyTV/ZTxKPt+g3P2VD6FxS4W6Jse+DHX89NbQQMypMmrdZi
7jO+gu/MfMuL12N16fE6Eaxd5U72wiEOGqIjhe3UFbPRwWcmjIUubscw7D6CnmTc7ok5lkc2LZhr
wAaFNfRLh2qW7CjcQ1Avcl22L/cKkEx/T6t5KsxJmFJAyTGsRPeroG7bxxlzyWH0CAbOb/4LgYrH
2AGbmLw5rXKO/uZ0sFp2yqbgQbMhZfhFm6THVj+9z+fs6xL5Ne0WWw8V89a3TfdCu7mm7ukR+BfN
DAwHf7xunkpv4Ap0XKi7a8hbqOT1rBLhifA64zEtiNGedifB0N6iI1luaxXKGn0zAUvEjrFzq/Rg
QhwSZc8jEZAUprNKYXhB0BZ7Xec9wTEKHtJOfAgJb0o3pa6SX2SB4Sp5p/CCkbv92zQecrzuHZ1Q
rXQhofGdzGzoJlbyN6TTdeC9pXlfHONUf4i2Px8+8+FcJ7tpwMd2EY75xs8NJ7TTC33b/UP8I9JV
qVGgg7vxuD3WklIyjwyggG/czdMAahxsbDgYGX4ncBLcoj2EG3M+uXbRxaMHXmLHmqWbfNrRv9VI
NYHu5rJc1qRaBcagNmJuHnp6fSXoreDoEdJXm/0a0S+YDiORsJv2164QNcSZXn9jQhd3sUXU6KuZ
MjK1XxJC3TH7K5UC+NuacckJtv6I4dDpfh3fd73nqeVimJ+aBQW+DDngkLxFvVq2h5ArBTi2fy2P
sRKuDWNhMlQMxeg4sqLCK25rSUkDKROYfBpgoxI+BYn1kdn8Vly3IWDIaqT/HxJl3C2pAXdOvb3Y
POquNAw1e2fx2yEwJQ1F+BEdNJQoJIOOE94gebacLDaY2408zbDkpGNp1N6pyj6PxWumovfw6Qrj
kkWyNKP3S13FcbNasMyikgq2ndA7FRbkaj09/Igpzg/zHmdTPiFYU3Z0NcupM8H0X+ey7PaBanDr
vDSUw7vxi3QgxRLZwzAzMtGRHx/jNX2BzL5BIPEBkTyaATNbEsZBsiK1t8NhFHrAQdABKvYGAj2B
LYlHeuyisbPyjOfZkrm6QAvY0EWmCsjiA6R2w1rxHUecXUpjptK2q5Wjih+f1DoGiN84DGdJA+xm
KchMvNc+W5N02UXxFzBcMWqxv5RrJvQZW0PmPfw4B8l33wSVJAIdx2z3qe4IxrY2c4JyQfds8ob3
LiqT11UJvqp9AGC9H854Emenx9sLtM4L50wZ8wrKvKLqeKwK+XvkB8XfilQ+QjK19F04Uy4aDpTJ
0EASzGKaR2zvwJ9mzr7obUmdSRySke3pBFcY4z+6pITgNJEYkYG6rItjRZKXWkIkCAdU5PCDCCOo
9I8ImQPGtPnuCjlgMRjpaoou6myOJwEIRXHUBbmg95bUQZzAUDztnfMBt04aOcmF773eIXihntxT
X8XMuEhqGkdoojm4VWMzhoS0N8872ICLTuTlyI3pw4INubaObNpkPjEkGsJNMfCwVOI1QvPC4LEA
qL51agjKGl4KwdxttIkL8PDTm5tg8k4PuEBVTJ+dFq+RgAXeSEgsXUaITwXWql5PgHDlCxPWblQs
tpoqw5HHXsr2VuGUcSJA899GWqsa9bHZJybs2zwjO6Tc63OHxAIJAXwJ8+NCn2QFslJxrGcr611W
LDQKtDK/XNHOoe2me3mDv2eH9/Izzg6b0JHQ/gYXDkMwgt88276aGR8/pa8y96yOc1VEMAYnhtpm
qI/I5CI1MfKSJSnxOJvUyxuIXQz8bqiZIIUMEQuxS2TTxWC8RygyICYV1gV8dQBMx7WJ3KhOXNBj
fFAHljDb3Ri5Q4Vbl7ee7lrBh8JJBtWsF3mBsG2Cz4uxJehDoEZY6R2yVX4f7M5mKTV1gW3fniPz
J3VkTlCqiWPoMa3+3HuGSla+PMm8DasNuDFGBY82KY7BGdVjfKXzOMUtMhA8Ewx/3gx4EHw4S5eK
nwVQh0Mh/U9gL1fNEw0zHbbS4ABufm81Cl5YP/utkCCYkXS8qdReDFcLx3OGSvL6mHRh6/63LSDP
p+J4LEVlk5R4J9XQDiI2SRKTiZHhwdCVyvP4ytlGGCRakjYY4UPsVLKkwn/Wcj9uZ9ez3s6i65mr
ufejbmLPuix91fg8mmzZyLk+AWAnl6oGP6Kj8JzBH2GWNpcU2861MucjYRh2Jpa3xbq0lqy3MKN4
IftYwPvivSZs6oKyEwjq4gAOilJIsCdLHw1g0JTDFrZMpnksn5JizfN5smbVexi68m/0LE5VvIxD
z9v2HhaCpzU3jZ65M34WlitYAvzU9BBR4Di3LqdjLv6fhlf/PfGxXLMcSZoMweieeHku06s3DkAI
c8g/DoaLMSLiy/IzHMKn5bpT3ZpiEnICrImf/NYrT5F+b/hNsbmzUyZjv/0ahZLPYE25yP+fj9RE
dyMB+ubv7bh1HeDLWjLCsdEg7MN26bkylENo0Y73Yg8/hDHwev9f1rWUwjcXIejRC60e4xVJBevK
zcObTjM6h3IQk7Wbp65oMznlkA93Kr00Fh+D95M/a7Gnsl7hbIgZl3IsQCZZ+K/RE/hCLHSK7YOe
Y/SOu7BCHitxXxgeo2kBXy5AHP905LhyJ5SHwzmHUAYXgHsuiRGwJBXlU+qW4SjNR/IfCRDWMCgz
igQ7ENRptkHtnW69Gd6rmBLbEuB680vSny4NUWoSSbVrUA6h/FtLl0tOuSGgStzquAnBh1FQnuwf
Yb82P0vwFjo5dK0hTER9HVOlfaFeuX10f/pHEeuv2d3zir48H4R6KFsufju88qcFlJ7OVP4oO9yF
Oc4CUm+wXHqvGgjU6JwAmgQaF4LGzN8xcxbKZr8OZZVZC8LSbN1vAX/qMoEalnyU4wu2wSYFOxQP
qQcTuBVjjhFkxALHQ7v4j+qVQn8rs0VcUBIIMbiYWh13JObLMnWXmFyb8m1o4y2Ek9pxWw72zFAZ
2eDbYsvJkk1Z6ejOMX/z8z1LaOb3WWLska5FmFSxv6rEmCYHzEyZiOPDOanxy1C5+eVyZ12E3zvt
oMuNxfPbU/6acrTwPJrDSM119qULpVCepXU7XXAN3TJy0eHkLDNy9txhppbby9QOAKCbYnH5ufko
VttCA/cs5BFkGKX+U6utoFFdl71VVJNc/6VM/j8MDwdPPawgREFi+rbKfrmChvbmO1uVYwP0TMin
XhUn2TskYicfHhvJbHGYxYt8aV5EnUN1Hec0KNYF3svr47HFqDTK8RN4tmu38o8Nj8I3dC2nL1jD
04vYFyPyPLH/UYYb9F7Q5k3Trb0LUw/+kSuRvPUElBU7IrgKnWRf67YbkbVmgFmCNPT0CBd1b862
hcpH0k0XxOSQLWwEnDCzhBGieKG/dZ9TDvio9UlR3IP3nJut2K6FoCsB5D4g+iHYz1FyoXRMQ5qq
Pe0Mtx2bz2HMewI7qgXIBLs3XFNAq92AecArYVECDzIt4rOyiyWnqpcGM0l/o0tv+p2DpVMJtvF8
kaiHS4fX0C00CYSOdl0KEWyS/taa5QwuF3tNb/0wlDGEHrRyakCU8WOUeQQ4BXSAKc9iSp8hHRgT
M5v0L7gT/61oluggKRQwyQQx9ERWrjBnUxr+bTubZkRddl6+aBDF43lo01IGMUl5ck6YCbYzF/i1
9IWUsop4QpCmI+F3LjQsIgk0h6G83kHVzcVgCFCVK7tkYjcuo1JNG0ziwdiNlkB+4AEkybjek3j/
jvvsc/rbVh16yA5wjYLMi2ZqFjgXRv1bbffYB1/1q48AcOPdhOl5yAfLNUtw2h50k1uyhTDo+PD3
HTOWxJFRtPdLFQ6sWXCbQ32DRfUDZkcQC1D4T4S19Oh3RMV73ln8g8zpVbl/xSf2vmdjDKKcshIn
pDB6Bwy9vkldqWSI2VDqPapIsVz2F9eZKrWa+1jXOEnQvP+KtiftZORWMrZ7dhOhsNVb1m3XxnBW
I56DJ8nBrYk1mAq4motOMNYqbZl82mIYIVfxdkTWRHPPBR0EWZvgE+CDdTgq7eG2zoDWXOTR/WAw
ok4fd/Jos2T02xr0VWelredPR6bi/emjzYeHkKSdHkkFsQlR9iOlECknjBsU+cDTgBXLBUGl1JLj
L2bmIBTp0q4ECbFxV9z3S7Ux3epEl0X47SVzq56BGsTVO8QKlRuxfNd42aTPjgMpsR/eDJvMabws
gFOhf7mbPINSK+zxX/STWc2YZvlWsk1/BezwgvzmRkgVCncqV7cSUkn3HkZWj/MkdhnEYFJPPXl4
Y0BzkkMiSZY7soTl8PgSm9CMssXfR9jfKUI/QJYqE8ljLMa47YWeoqNfhjiFUZIPElgy8IeRChcJ
eTfAFRwHVrcy7D0HwYwq2IHVKPCGFftqZqKnRl+1/fguBw1u2mPayr7uE0Os9Jy/D5Sg1Dh32DHv
QUIXL2MSzEFFqxOSTsRzOeju6oo8Oo1yxJHYrBt7o5mMGgpXBhKw7PgWt09iwtPJ/3/yvpTyNyrU
+79s/rZJ3lcmYQfzk7a66A81GL4j7Da9jHlUoiFutdDavximgvOQCE1+oYIxH6PAmhvqKO7z9wtX
N9rMVsjz1/k73aIeOWXDlOxYSx5iJIjr5ivdCJHhgC4EWJLxQinbTr7zk01loVW75yOLqKrCk7tW
m4VFS1iMRJgaqv69ntuyQajKCf3AWWbaqHpRXVN54D7RcYoE+LTq/Wkg8+ipGWObYBeiCe7cATrF
mrqqStCEBAz3k965GpY/p9sW3VT9YrjFIDnT+GtcpX+v0LG1AjlpaCFNPVvpPc8Kja4yokdJKMB/
3I4xO1GI3eKkMRkQ2iH8xUCemhhSP7gMYB8JLGFAeHCkiOXZJYaXRbn++lSG/hZpaOBT6TT/C7j8
rRDpDmbVqLeeDOT4mL2zPaEGmvET3W5RhDuQ1oumH+DPsX0EcCeTSBRjZ5x3JDJgowwWb0XCKWUh
wPxWY4a5DJVL6mpn3Nmi/tjb7MGFxWzGPwgWP+FTWNkvCZGHbqN7PSQaw1bmihEpIGG1SKoglJ1m
jh2ygL8KyXV53FOYo+jhODYdhxEG35f9ZrahJURBF/Wofx7cDynu7e2GDZ+itpNsZtNZHEiaQ6uk
flhlNBL6fEk5hfMNc0/8Z6288vqWXJsFPRGO3SwohSAT/FrA5SpM8Wq6WmifyR2LJEjIKHNFWzk3
LzySeC3M5q0HBGyj7PqL6pUATjY28ntx+Eb/tnXck30EEv6L8qnbIXNqZo6kAHQIHxXryCluQ5Vz
89Sk3+op4J75lz3aS9Fd/uE3Bco8YialvSwzLLrcOXlK7p2+Ld7Ajy900C8z5gO7FWJ2cjBkXcka
09C3HLoQvvF392S9hS51ctE1Hvh5wfNLAfavaX3oDJZhTVLLTth4bU8KkT114mpRSZpKH5ld6W2I
jRlOmEHO7EVUNrAWYEz2cqQJHpeN7OrCQZuPrlZsYdh6g4S11OJ/Y32nY+UNpVr4S/5T7OnH/2bh
2r9/3TAFirlvBgVhSmzTn3EP2aeX6JELjFIsx+oP5/MXscY04shoQqgBH3acMxJpoCpk3DwL9wnr
WO2tNQu2coacMs/CgzY+hLallZzq6jjnHbIYO1OiwwfGwL77LhObmMGFDD/yBJhMq6kuzdJhcchx
CKC4SUyNybzHbSDA3ZranF5sNbfucKFO1jk0DesIcw5qxIz66uNz+g8eDPN60M2pNMWh2cRwYLN4
HmS7ODPel9VP+6SuYv6mybjdncuqFvA0IJkSHU1ngT+QALfGfXU6qkf9fE5/PgAFqqeRVr5sPsIw
gKU/GGY4vcpw45uNzq5TXq7oKcZiIRNz/14MZRBwnhPUjZINXWN9HVFhCOuHe/rh6uLRFaP27Uqc
9cArMRS/5d8N7/S75467UUFwjBnX1QC09NUuuJf46aa5+7nOdbU7ovASNYuqUKBkwnJHIyuLD3IB
/DIG/uDRbZQ+KuLULYlrQXqNLQz0qgC7Z5eSr7QxDUuFhYRbumkDkXkcKhDVVfyxJuApvqf54/2W
jv0zn3EDVhXpnJQcMQn1+1kwaE8H4nlqCLPSY47tSxCLDAhTnNikoODLpOMPVKJP39xUt9OYOYGr
5WPihYdv9BDdMsRLH0WmtnJGZK+gk0LYKo3G6RebBpBvvX0AuHKx0s3bhtadmEYEasN2+O7SogP8
JfHMp7CO6cITTb3Tvmyx8U3JZbtIDr2NVxhsK5tyl2S5TcngUOS2nPuHDJu94pSVocxOrhAbrBU6
kyYRLjyjE6J20nwo7jj3bTLnVisM3LbpmjyGMbUzrZlEOQRSJ5jBgeXnLtgj1tbiFWB5Tu+y1gcz
Q3eMZsUiJhtbBaISP5lu8bCEmyKgDSVHvBqEnqqxq1ZxfY55EzDiwBShbzLwI0QRtcIuenKotLUZ
gPpdrlJQtAmYIT1QQYXwTSHVclfOQnhazqTkPrVygsVMknPswRyCXFXjkmMpuI0ALNjj9f3btM4L
tQDARIIrq5LL+1Fs5O6Uz6cHuuDtar49gDi/Wa/eAR5dlLJxkWgYDHJS1URLMqD7b8ZviJdXOUBr
A10KKsskcUVKKS4Yvo+N9+t6BtM20h73XoSrFId1JCLJLibTe2jNhxfDjzG+3cp41rxnsHjDyLzQ
N9etnHSV4FgQHbm0obFheh8tomeZDcRh87DnbzLOrHVd+yEMM8tEQgdVQ3CLvbLLPP/F9R0Hte90
D0IH25mMBA3cFtZqz/qivsMkt56urgilmleSHfWqiXYYjmg71vO99RoYh6alfYANpPFV4uwursrK
9uts180jaofYd5qF12KFK1bk8nCZxDxyUDS5GqDnRGph0HGKbNED7lHue6c81gUTGnrxb+eVL0wQ
3T7NMacy5QDvJijkqJEeTiU+U/Z7FORR27pOqiiT2BswVbf9HTbpVBb0qMGvbdiism8geNpTOxZI
izP0IijWn2eKM+HYitoxarBXoBu/RUESJsbozg+ccSA3LsSmMjVUMRmuHx+V9R+GxbIK4nXPv4Iv
gW7RGPw8Drs18/iCCyuCbdkGkjK0IdLwpgnBRRvlgLXkeCjqIQkYCfwGAu1aqN7i9DpBN6lCWPGX
K+4AK3f1IQNXEUjpj5WHMNzOEbY4oluGI58QEuyrGU1V2XxbL4ouVt3U7HJDx/nG2REgT1dEx6nw
po17YKE+pafvgi1TlPIg4Z59rNRttxkq09p8UBa+DyvyOiz8gw0KzvXXdGKQwZGrkDy1rMmBdRQq
mKeSPdZIKnbjSankza6PSWtpkHixfxo/g71mVvs78lz+HCYPY13L/YNrRdM2ho4de5wRvCEsnda7
CqTVmt+cmvWHNgf+5K4JFKUEGT45ijqlRuP8tqMp4uUGOMagbPdXDNcJCasSK07GqpOvFspz747G
lynzN2C3VAQf9E9xwY79CyLiYCCHkrRhavk81Ijc6yPsh9SmxQOAJudMEs7stszJJSJHbaXEWUn7
2sTMYj2nZKNmKzImQ928Sf5vWcO8IBs3zGraKVsNd8PR/jtE8bgBr6hr5qdBCdL1UwD1psypn+LK
LSFIa7s4QFeKN6RagA4qB/4Vtuw58V5dqcCgjkcZyTbXfgF06WrM3aF1Dfz/XcTj5Ro4h4Sz1pXa
6Wxo8ho94mKwcWFDXBrnOqUS9dMrLY2bUmV5dBi4FxEDcgMneA75EAfjI1w8mRimJCHPF2llvy/W
c/gdH+ewW/tAUy5t88n8TUMIatVBYpyGUDy6PGOJ2FP65bVq88pJquTP5KMldJqMyk5+i5ohAGEX
Oj/h70pE0n8KHoE07vl2fuROgb5gMySwd79qpL0DBFEJQOhNr0s6zDpHBiZe2XQ74ogcNtH1sYE9
3412J281fvrmvnDlBKlcY3ZHerFOKO9g1ekwD2oThfzSj4HR1X2xG5FjCEXcmvM7BCS77LYnzWHU
eWR7uD5l8CE2jVdIdKSBbbT4Z5+LgXQzNL1bydtFwK/+CHAK3m4pG+MywrEHxOjllb/mBXzfcCn4
0AkA+vvr3Oyq4C6eMtWiEfkodTF5V826vf/sZ/d6/+IEnzB8V7LNt+bvbiH8F7+Uwer0vytoUJy3
16tgsN2C6NOzn2vCnNiAw0VfSjurtIrJ0K2BPMk1fSo0dswnmPyucI27JVJ+OSTD0sTy2Z7DW/T5
9GxpDDRNrKx8CQ48mTosKtsGNa4rW8Fv8/R0nV/HiAruAy6D40RUq50fsEVz0q+J1pVCNxz2fz+k
YuAsdLqNCyMBvZ4m+6m476LoiStbHRNCLoN4KnS4cCVUmd9DrmD1BkKZhe7XSf6Pk0wsIY+dLBIJ
rx0C2rN9+7yn27zzM+HHRwqlKPpPwa02yGNcSVx0IibDIew/60CV6HaZVWuLdH3w78+uR2Wj8b7a
fbaFqniW7X+trLlMhWLUoFOKMCmrrY8ObpA8sxGF24Z66WF0/V/7o93GpST6DK+HelYLjFHlAhPT
DzB6NaEh+Dn4BaJNdZbinOdRd5ucyQ57v9YBZYZTep4xHI6fquxUQEgWFLg7zWLoC/Wy0LNHhqL6
aXt6fZGCrMVoRtfX33KIOdLO0gdGBVvP+WFv6JgoSf/RtLrz3ovF2fP+lq+FlLprkEmLxcafDlVf
nkxLazHKiadK5mKTMgcZai35sVxMc09wnhPThJrh+t/hjV2lT8pdHE6JTOMXj49kJrWtTjjs+9Gr
zHzngm3Lct0hmaergBwBIg3UjZ7uP/WgUzK/ufx/sKXmdve0OKtcGlQ1y07G+X7LmR1bS3mDLNJI
1TmUyiE14OAuAAB2eBq9jlZ0GSeDsb7jsdFzhMvDHoYistM/fXHTxumC3kjzmrmhxCddP5Q/Atyd
NzOBzLlLer3thAxDCcS+kKqgmxdFA50ZaMC16YDO6zlPPovelJp6z88t9G1wnjvH+FfaZ3CuMvK4
DRa5U51AtJvpCmTdm+dHggdqhFfe6EPU3C4iyq8jcZsHp92/p1D2eRztxXOVdaTWW/Ioyzqa7lMz
FM8CLgEEnHigBcG1OZVxb2UGQQ5amYKTNyHKZhpEYR9CH3h6ycl1AgTLoJ/g1N37o69ptCv/ISch
NlicniJSX+d3KQJ87SIAZU4VaaWz/zsVMuoIKqyRB3fAdVv4Ai/2LYyJP/Ng9z4qeR2lvGKjXa2V
ik8cQj9xmuzAiFBbi2rESu5hLQ0Z2dgU8mvlf1jhG7DX5+hZHXYQoqLN7LjVr0AaSuBa+AXxUpnf
25bXkUHAhHznLWPhBxgQopfkI4esvImJThN+M47TPTF5nLxityHSNnbPV/nOdgVPoSmXg/JnJCVP
yyWKE0Myear5ECyb40uth9UvO1nyPME0doO45eusIKrDyH8DILO2BM/IdJTCLDQrsiSHE0+fwSBN
go9nBokk2Px9IQAmDAQlZUbM8sqTLkEf+bEghNjAvhozNP5ehpRuHK0biXaoVWUmln5qIwJ97joM
SHDcwfwJBS42ch0W7P4TcP4MsEFSBe3dq1H3LjVmpc5oHUTNEgxU2s+LSrAU69r5YGyCi/wy1+f5
uWhL3INokmiIH/IfYL/gm7cL7/D015s1JnNP3lkErZcamxbbOr5Oon2bsGoM4XbOx05U72yX9hUO
W4ZoNSj9yTbBHZ4jeJy99fe1e+TyPFGOJ7LC1h0ftiAoHj/IIPFZ4de7URoKgjXHsHzw+4quZkRu
G3afUOX4aMk8P4ZrHMW1aZqEiHJsV1X1FIOLlrxP5UmblzKSbcHc8ZVhzpE1+TW0agzm057EhfHD
irvrQEwEO+zedcf4yAZ6UCCR2lQalj9cjaO1lUEaaPf6yksWQsmkgR0b1WYPgWwsL/akQpJBmNi2
wEMC8NrNw2VjzkCDPsunCqAElH2Sw3hY9eEycTSfg680boQoZZbV2O+LyHrZR04gc+6HkUWZK6Kr
0IQveClRnTchV3/bFLZ5r6FDkL0KFEaGWUudSAlV2Ea+DvMHcNP1i27MXydVHJ8wQqfbUYCLoxmB
SmW0eTAux+YGP2GRXb7P/+wNmfB9QRK8/uXH/4Zv+Z7L37BaKhAYmCDIbk62YUXOFNyJtYI3uUbI
LyZZw83qaaEOXLN0pZz7NpvkxIkMNuF27Pxlv5atKJ5myg8iKTt4G8SRFqFhc3pjpq8Y4ti4nNWY
3rFiFuuipjnpfS2dcTUyaxf4CoOhfhj60zqbmtt6659HFMszl0gZe93LRmDN9f93wnE3KoOKRmRU
Ff9Q+qbC4NQst/dYhxzEBCJQJYdXBpjbwC8X2bDimNyFTpgHbLt9NlgI+CE/LS8r8jp/uMO6lAp/
4joHZeboSR+k+PtK2p97uh3fr4voOoEW6JdPj+uZEBoWMXO6tWFF9WdhVhsWJgO5My5bW14lsBDd
oRHtZNSEg77U6Y0NVbzf189HhcJVUxXBvsxMnoJb5UUHITrI3WIo5JME22UOIThfxJTiNMbGFp41
Wrkn0A+4HorcJEAkbHC9aDD+LhC+wTgcIkvoDjar15Im0gwy6a2K5+Dc5YllQeyMS5/vrrC0kUu3
xp9QWfEdtYiQCK9TtlB+Be4ZPpmjnjjwjFlAsQLblG9Pq3E5hUnaQ6n+h0iQptJHHSMDcR2iKnG8
vXGHtaMvODIz6CefhgdGr4PJUMN7GZ7sz9vHOT9TjkJH0IpNO34WkRHlfuQjqWM1oC7j4ZYpIvGk
8o92jntbuH6E2PXtYpuhCq5O/9AZNSonS2D4q4/vdIUHA5vaGBuN3cyckV47m/lae+n15QsoU+rf
yQaM02evRQ6cLNMm3pYx5MIOrT4logviI6uMSR2FEBrMKN8UXSd6IaCJOATR4rxfRy/Ev1xems54
6vlOjsEcVAKYEdq2W44bA0Mpil/27cqsrG2nlany2BGOc+Z3zOAN44s2LZ3lFr4DtNXIbL+1uUT6
xMl9Heg7jxOVUvQe4MaM1Jp+G2eSh9j4UbtNPW0FcFr3y5blff5XtMXquiEsKqxLa9Q84sVe63uz
4w/8/MzOP8YE7TznKWT0oCV/IYWdLdekv2KbQaPWCA/eeDzOTbSZEL06jIPKme0wpjpf93ZCw/E9
fN8u/9Ti22QXxzNOyhMox1BcbivPHpbkdPgtWlpPFMZnwfcSlmFneflL3Wnx11xhJBHNOPdx7nNU
Ft6UiZ8u8qrNhpcV91gVfjQwcyK+xfQvi6ZIqE8f0zS4BO65ogMALSBNyBNxcJUvG8JR3H7huiYn
6JtUGrBC1vE0CR+/2xGAgzGn7yV5F6kuGVjB+lZsV/qogf90qaRs79Ljr2h029r5eiTV+k/D5xBj
LLCWhyZC2P4Xv5b/cU64kuG8ti7SNXKUq1QnwZM9ANNdlF2LAeXDIQH/3+UMG6l4m2an8LqJWJgX
lOlTOZg1nCoTfp8nMqGfDp1svSqzscc3wAfD6W9nEsEj+7UR+/gJ+9pMqZ9QiNgNGGYjj8fRe+Jx
3wXU87oAy4hCEw1gkKh1GOpHq822uVXznlwfq05WLE3L3fs8tLHyroj2mN7+4eAjgyS4GxpHcFvb
CSbe31ZT3+Pi683n6jnitKg0PaKMq8G/EyQnmUG67Dxm92Xb0yOcXiS7NqFxJSdtJlwKE4FAUmoa
MT2EJJXsUmfp7oG1BGuxT3PP9fX2lhBfh0q2PtDoLPQi8ZHGeIysZJss3YTKxjZjrNRdY112JEbT
BmP26PuwOaApbCZOCYRcdCFAChnYCV5566FqSKCPM9WjkGK8QmWl/Fx4qUa7bi+WVzuIboj6IHtq
BTtd074tccHbKG3u+B0cYOk7hMyYRtWj4PW0Qz7cg6Aq+GmfMya7XloI+lSyKfbOh03NmiAkYK4p
wpZTC+eNwa/D4hwUIMRNwJgFLmPkns/079eGXyDDDprF+lcMaO/OgTkse9PcLxaXRPN6j+9R4S+R
CHslRhzMRKHGITi+3PTmB9wbRu98qcMFdw+C1TpG2gIKlipjZo4a2NJU6OnQFT2NLw7Wvd8P8ZZG
46v1xYhE/0r8HJJ33CafEwPXgEUhGrvFvJaiEkN0HYhHCIRotag9x+g4xuzRYBABpIikeCeWZWbx
5VUEDK8TRn5m8yHNpcrUNpzaGWYlkO0HGuc9dQEfjD4fo60L8JW0kkf6iyyZx6BJ9TCTPFMXYq5D
xZ+5QD8szChYucQVQw1U7v5A97Y7H2QGvqNUqqj0+t31WSIbI4tYEhB48NGAXghuH3/ns6ZoM8mp
3pnW9/8Zw9pKCX9j7DC/0NUPlYBZWMnQv5ejXHcncoWTJ1+9entk6VM23LIyy1l6aAbs/HRn7Rzx
NVsTa3AOA0hMGMsFC+DixgK3Qj9SYXMN6x7etRIkqoQj5iW76ogLDPBkhObYJW/VjNUlEeaW9tm2
EfI3Vb7B4814i+3RuKyQn4DmSEZn2cgjX5MDvxen2JHJAH1PiO+zTGXhzA09eQcjI5DaD1rea1JR
oBF+Q/2RgBYilSO9W3U5HKIwYOtyW2rFYsb0/0yEV+aF+WpFxaxmMbEMBXBFQFonNIzKi4+hHmNj
nhhs5N+VjPQRpKEMyXfGb8BhTAznD14HKAkWlDdmukE0I4Qg9ngE9b6HuIOL/U/uz0UhNCPSj94K
MLiHHHp43S06CBzT8M8G/18N50UNIXvSFQmFPzYOvmXsg+SVZS39GUyl9VU7SorP+06IxL7ZLKFI
Jv9x+EwaJFlLZr3NfAiAkuUIsZ++6uafLLo+FVXEnNF3ovNO45O5EOjogtio5skUc8B+PcnqhSR1
VvncX6R2RTelam+5k4fb/mb7RZz3Lftclop69r6QpfJe6XCB+xomSX974nN59JoKIvGs3BkPzBsY
aWhq49oQBNBVFcuPE3/bEIkzyb5kpQAMPZtdg5pqiDYixXHbp+ZSxHxpj8MVw444RJGxSkA3QryE
BU4QbbJ6ySBvEIomYmf4ihbavT0rv4GTfv8yWY1+zkbn5ufgxaWx5AX1FtFqRFZdHF1lN74F0dpV
Z/4RgE0b0kegHUqeuf9dz7R0fnb26niEAYfVW6kYY6TWtlSepCUS6OkQ290ZRxT8gbcsbPxyIHTB
D7lBKJ01cYjriq3gSt/RyOkVSD8+kofRrVijAkxy0r/ke265yErppl8y629d8EBVdIRFFhTRy+D7
7xZ0gsh1eSQB7W847BNLxGIbLelgUeoqWliPJKaAJ9TeH8uT6F9Nzkz/Hgoy1fWms10xuDVZ0/pd
qH3YVU9MT6PfTq+YGXogwgh73onZeI0VeS/yAoGElFVa26YsugwLSDiJcsPZzPWPdHXpu7pxIljb
bAXbvU21qRfZuIl1Efl7983ZyGqIBjd6HvNN8ycS2PlXsM9qIAyIc/51CjHZudNI6igmUwrtWzS+
XNf9h6IY8OM7tqKALzssWGil7lXEtleTrZWcXfmsHzFfub1UeCETNpfFoJRQVWz1+78E0g1JkEgJ
USxDLw8rzoUjCHqQZfGVAHfAkX5pVCGJhzkik7Egq8FfNY94CQ1A0QnGOE/LeOVFDhVWhx49iSGy
AN2Hn0YlndSYbr850Qii5h6M9+IEGD5IsHlOQQ1ta6PRd0sQvJeoquxZWe4oBPyprKVzKCJ6wIgS
00QT4eHmv2yXCwqpuMlNeAvFV1ZcvKbgEVO0FzV8SHZy6CuKxbGGknwrxr8KfT6nORABc8SpUtfe
WYBXih4eC5m+ftPnxp/S5G9K1Am6iDamxel+u3CS0lqRkOZy7bDArR4Z6K3PMuTTa3LzewIjPEme
JK+BCCCUVG6GcdDFILQUTEFL4uOMz8ihf78PZy2e/1dmQ6F/RCLkjLo4lIHxcFI/6BiSzIk9F5oO
lTtJfU2aOhUs+zpxUxcbLyzwP/FhIbzTq0YI6dIalwzIqunb7HSTkc4K6Nt4TmakaxCqtq8DdIQv
Qfnvpy/+QF/pwjUmc78NOKjn7cfYvXAbRUkhte5BdLXgnLlw5OWnVt/kGpk9zS1d4f79CT2hoxK7
iw0+xgLo62/T3P3KOXr8ugBqlsVUbDd9Fqe47ih4hUXCkK9ipUvrInliKQK0jFf3k9SMYbUwyIx1
n9X8ugcayptgYjI09pIrGuqquA6TixS37Dv93kVf4rAPDalp6lzrTq4YBaPq0mAccEkJfxo0xnLC
mnyqiAdACKDargB7tegGDpiErXfpwWFTMCoG9FCnCprnNhHX7cHQOJe0/Y0fJBEWCj2YBAx6iXeu
h/PcUreQ2X2Nckoi2ednC8XiFwmyFIImxjsFZnRZOIqMaczwMtTxUPHEOaDshZDZP6iYeANNNIFe
WQmi8XsIkdyjbKso4AXFmfDsyNdFO/kuG689ngUq2b3jRqY/UmKVPSCV5bUD3YdWmZFLsoEqJTxA
aGV/gGr1vSFb9vWa0fCNPJVtNWdAIZygS02IQdIBpyo3vjuzJQ6pFM5YsM6XkMNHyGdUjSuM2guJ
GW262g/E5PmBCWNJobFLzKt47FZw4fmE2uJKa357R+8336w39qdsz+AK2IVnH2B/GUMYQJL35ndO
yQYsYOJUku4ZdJByqlpcOnoDM9FPyuTWUZwC4MHRhbHUTrdswPQ+wddiTKRU0SMhEk6Tn2Db01n+
S7WJak2hRc1zqPbdV+9Pk5VnFDpo1NXORfuqSIJzLUdGjnbM5Zco3YvqUXQ8E8ulZix3SeevAHEx
roh+9aDizwgU1M5l4dq0Wv8TBvF21NcMkl6g03gBQbHvQ7WRuQWGd8KbHHkCnn2QcTofADIcWJqy
6MSI5Rl1E8auk1xrxh7hWbhYiEaewNlbmoFA84bC6ZHWwbDoKthdl6Kx+ZP0fSh4JKyyltFyeLKh
mkffOO+aMHfr6b121OWObUL091riZLU9Gpht3IM92lFx/TTX+K7inE66n10+l2meaoza2Wfdtz6S
N2e6TnhGZ0wy3J+IZBq3RXeTE02zhr992QvPmHdKvYgPOEeI0OZD7CEHoZ3ylqzdeBY5ZVwxt4Nq
OzHg4JR3PuSb+bwHOpJLWjKE8wfqQWDhNsEEzM9zIjqHciq/Q94mX5yvZt451l2uEDRZewLllH6h
nVJKK+PLmUQStzg3StjgACbNFpMhC/aBYWVBlxRF2mvbHRb5aLvvlKFKAfzMxZ3Wpn1nVnBu1F9F
aw5nOgidy5+i/n/45/gAwlJ/NYas7AMnJCDlxUKHyWLuOTOgQSg4FnobtWniZAzJtmQcfO0EC3/8
rB3iiBL7TwPUFA44U3sneGv8bJogb4I7RUU9uDrXFk20iB1yMsJSbPYMPgAxSfXWflnCj4yZXoKq
1ILJB8CZJBY5W6lB33kgqHwxR+NgtxUT7njm77odUQeUBGK1e+EXZy5CcB7LDkN4i1vX4SCosqMF
0Kbpm3SXax9wzjNPl40Bxpq3Nws9fsaX7d+UR9G6IUylhFhov0THpP6G0vyZpF+y+K9qc1UO7lWz
OwQTHmBiczGTLOGYm18Opxj3ZlgEom/UpmXuMDQsoG84dePMibPkyT1TtHTjnlXRa7k66ozRLEJy
NjKexvQtdXs6QNXHPSzBnhTV5RBsODe7Lfc7hKy3CG80638F2fRethwG137xk1xd7e7gx7U0/j/A
8OipbTDKNACmFSFbV7wQ8ZTEPT7rZhPi4U2PUwAhulcdwryWkQhYeZjrkzF+jBjX0s4NlifU0/Sw
TJSxJMgq2lj05g+phr+PR+m3sfgLYtyZwlTuZI71RlIo3AB3lfajMIm7cKiFt6ZXaec6Q0qqvvBm
dSVFwGvZX/18GwGGHz6/COhpaj4Z7ObKVv8/PTSG2+7MpVLcoQ3EU0Ffl6Wb4flpxMmf3kpvRGxC
XeSw1h6pI8j3PvSppfEGrIP6eOOzLENBG+DHpAXsmqtJrlpZ4k1ohOu+0TEhLlFEz+8/Af0TKWdo
N8FKQjR6yh3Qa9y0F0nuq7V+f2pZOAt2l1NKWiDg818IQGN4AgJ1xNKyFsUI2822aa+lPfK/860H
0qwCXZcVb/6/5k16ENv3mso/IjsYJsbE1DF/x2x3QPYXftK6QAMtrloIGoTYCje3MbEoft60xphp
qW3x38d2uE0eqVOvP6rDPvGOX8drpqg0Lzwkmj+/kc/fW0GE19UzVnwNh1xZvanCpXsXNOgOjKas
3fjVFEYVqmpO2YOY2CZ/qy6KUAfDsTUA8IJwRI5oa3Joq457mnvw6lDI49ni1UKWD8/S0WfkLrAH
JCGOGvo5BN9WUM3WjdU3OnxQpdMc3eX2/KHofNjgzI5V2CbxBHbU2B6v+LYstZwbgVBGJsYu6j8+
dqWJvVGl5ILHdzGoT8VYRQ4m8wsvTefKXvpdbk/RZxBkHT+BF1sXda0HZUVKxxjCdK5mxRbfacSq
rOnZs8lgF3rpGDrOm4dGb+ZOxlU8dptGPPppuQqyVA5FLv5cBJHBHcWpDPh3vi2hbM/lkcYc6v+V
fL4vlnfGqodfjkA/r5MzG5sxeQYmyBNohhpCTkqzNjLBMmP5CvNAbaK2stdxCLCSF4G2GGuwUzLy
uTVnKImVM+wjEF/nIPGFkRUzDeo6xv09wCZrrD/kdJclyb2UH90OAKXpEFq2r1dkdLgi9xfBz/aU
nhv+szFjvZMtUiwMV17oxE1Zj3XIVvsvxttnNND7ivRJQioHhkGqNac2RYy0hwzpGEWKuX6hpUFN
9TvAcGoAzfMA9GB4CfonlUCNOr7uyHlEih6iXy8pjCm+fOJKfZOoGh3xQQIQZk1+hhZRmgMzRoi/
btp/j01na2qzwY/GR7ig7YlBwkDKhv89KlFO8+vBrPNhtctVW7ga4Xq42PLuK3iyXkEuZSDeOtSE
Z+zt/jrme8yghxP93fJS9tQgFjpp6Jkvbif/P7gKu57RbvmNXDZh4KrbeLwgkPlBvC0GzqFgBUeO
+BiwiNM2ntsK3bx1El1sMFC4jHcL2RdUdn3TvGI2gr3A8z2VGyDl6hgUuylZs7qHEhgIPue/d/Tv
b4RpcxBnpj3Mbj8NNP9tRj3hqN0AgTuT65AsPrSVowpccxf9+nX4h4oAhb2+20ml/m8iYs/AL+FB
cxb4GW3oGx5m8lM15K1Wy9L7ytZPmp+LPZUqZr5HyhycS7XHPY4x3IpFoj2Z+IugawfREB3hDIvO
14pdLcLlrMCM/EfscFsC4kLGqFBA3LB9wPsJM5vnG8XBizs5r0mdYhH0xMxmR7AoPocKXLIYxeUe
MR50BnNKfSB/Fp2cpSR8OZfCJli+VOU0t+76JYWsisLn9c5Bqy5vTMdjdX2X9/tCza99lVrFQLZA
c0WgNl4oTFnNIxyXNIhzymQFYNuAZQQuaWCNp+/rLGVyGTrkNDA7zfUvZmKnjeTrXYRLt5a1Zqbt
aE/QCqLTC84uhuYu/aF6H3X9s1qw8eSWJjLXP3rmxwkKiC8uyJ+BXe5CROkAJLSTeICK80BwzCe+
vNyHbvyk/TlPmjnecv1vVXt5U9e9DjX2AB2ym0ylBYN8zYUAOWQ9VxK3l8Jb8x+EWoErca7LSJH9
imYAoz+VN7W6g67KHnUSMrk8ExUtBEagp2aNFISFJ9WxTnB66oWQM+fDjwczq2eTlCBMKteywRq9
KgShEWsKHRjIUhbApwm9ewmgfoPlvUEjsN2gfBDNbpvjGxDC8Ih6kYJIPGlvzgNl6k3ISBGEXuU5
Uw+7wbrOy/kbXuGkWoGVPv6TKSqUEpe2CSJv/KdY2hGpCulLr0Gm8GvipAEaqjWeYki1UbScXM8E
D3sDk9XUqE4oxDmNwL85VIk4IGISxCoqNOXihA0jNyS+tvkvoIPFoY8Sl1epvkZpCHjyX41p/SAC
SAONhIfSvW3uJAoFnnmSdbs2oRI2X+oZpzhuFkxOBYjq0dpApoi8MwTbbtCnrlcHSGR6oNGaTYWw
W3Ir329Pn4m6BXFkltnGPdXHqhuPiY4tTWkFaigPrbT6lgvxxWDE0x0M3grmEZfGS5N95RSELr2V
mkB/q/AMaV0XfSm6QUarAGr/M+dSqZIuABWCN3jlkuxF2flXWbLirXJm37sW1vugowya6ozn5gkM
ulZNzfZHbweh65zzoovK+VkFGKgbVBw78XWIrygSMbApCq1MS89vNH9A4CXxGvcqcSzhXWFCDVaU
yzHTS7U7XPqNNacHi1XUocV2gmrUrktV3lz5/KdP7+bzi1FySl3Npq9yJAfNXlvSHI076Gm5NJbU
Gp/iuxpPRkVfQQeOmW7ijVd1873FHlHff6YpriGDS0mWsW2uQ7yzGMpJ/TmSmbX+ZUCTBW1lc+Pv
fpIutJ06HWWDnyjYMUcS/gkarD6xb0dzp3lnYvRoZ7WlOdCV/nlcB80pZC+s36UTJlxYzAar13VI
eMaBzO2wo0O2z6EYGNGiB3pJihXSU5ScqzqDODpFiDHrAKK09w+qnC61kbtkSEjh3ZNc1m3Unxfe
VW23BS8aOjsfVQeJE8M/puLG6Rfve81tKiOE2cqWGyT/BnTZUkT6VCiHtxOaLV3Fd7SEzfiqpANY
isyZyv+7krsGdVb3J/jpoifPjUFpv8Wkx+j1/7ed4ytTV9TjqQelop2hjRqLN1t+Vs4Sma8cxIQh
8Y5r2fov/bu99gljSbaOQbnBnfMvy7wGbDsN4nHvwGUgSxSAPFm3zEvR6dLJ8o+84JiQWs9lADxJ
NULmDm1tpl2klyqn3F79njJHbKe4hPqEFrJNi6LdnMTdQHe2RgNm1EENHTlCTV8HXNr5cIMBlrwq
9GwjWA66fUSRs5PAI2OOZSGOqp6tWvcoMWxj/OzEWzMCIynfS9Dx0LFaC4BxbXr51Uxk26iJmKAo
IK7WAxCV8co+T0Ey8B8GMF0GYUaPO1AihooMlbq+LNwOQ46SzUMDrlWYfiHleWkh10c4ElO/rKLH
bsPPCjUksW845ira5+Qpafh0TXcgKGIErckTpjaMtV4m7OrgArHIedITTa9sKXiH5I4dQCHY17mU
wlIlXVjCqjJnQ+xKpTC8Cu/wqFyc7aBEJD4y0Ri3Lk9kvyxxAJ72XZCy2lH8arF80owEANURSI7m
gdbJ/0nCRMnPSRTBUJQm7qSiGrxI9gWDQK7IPizUVFZEF3C0gzsIIDgKFhFd3JsC/cob4Ct/+cEl
MGrAvuqYxcf69oNCDkkYuBhy12HpUW268kFRM7ts1qH4cORWeSL7OmcUTDxnd9ZnGDiEjaCyRtse
ioNM8vmEa6yqDM9DjV/OrfAePvAJtJC/X09O9VV4fq2UkPR+/mYRUeaXm6pfXSmanGK6xsWUb4+5
jNXHKOMaNoVKG95nvG+HvfRa2sHJhO62feej+9yPcrTPwbYsjPOJztbfPxoKcI50q7bBjdN78Rbm
VH0XLTv5ugwHJ3OEkyNK0rcwTmUNEl8K2ciNqWcdOJeVMgBYvshOI4rr3r/2ExF9WRuImUgm/7gt
eSKHRrwSRoNvCsjZ2PgILaxlhGT/MNND/5s+T1bdYi4Ysff2kGO/AoQGYYHdyFyH1VtKl88F31yn
a5gr+uf37aSPTymkSqa3MY6DynoGD/d7QgyE4rN8dXjUPgdlwU+MkY31VAh7Gk1uykVPnXnJfOed
/WSgTyEcsLj85U9MBFmoyCAVtn6eEdd+GR2dKNRuIl0nlppvXxT3Bdj3EA/WhTVu+jpEY95gU2CI
trdEnUIOh8zKV8gI5feJdwLyqxgWi8PyHvdAbg62hHfh2fCmn142+/inS+rmYw7mwn8VLcc2rgMv
y4al7AtYuqCCcJcLvKoZm9kUxuCeyJQz9tNT3QTdd3Jbx0fEn6OwXMO0reuxwTYUQ9t+qO6kXCzb
xzAoNy26pgyXHk14ZxCsV6hdZIKrziMkGQklR2KIuOEgTmDpb17f1iS6dfBv2cOHHLtKDLOcIkJV
axEXsvlWZGmaEXlcCARYPrUjT0ZZMcvtZ87Fm8OlPQOMxNvsU8Bh+4+jyTt3o7HesAjtFdlHdMj7
jQLQENm/DucQs2vQWWD7JK4gqIT8+WW21dSOTOcy3bDaAp2TnK2RrerNwdlDZ5BctkExcj88TLAF
hSBzfZblkt4VDHYXBC0C+ESPBAWS22nDhw+T9Yv2fXL9jVXRzwyRMT8fWs2uOQq6XuoiKJGld5Ke
zjWBuGigFp9aZMoD826fcyrDAKI5iPZePrn6BBNyuBqDwk1YF7uczDnyia8XDOAqdT2O1z42crIE
wniulvUXuMYUfOJX4NYc9Xk5YnJKLgCQCSDBpl2nF/Za3a6uTHMRNZnks08YYAtJZv2mslBBq3aH
bcim2gkLsNqlsnYsK7Tw+TTTagQlCwdFUxkMoo/JD9ChGQpO2MACRmqFajn/WF3APlvyCOrxftg5
NEFgtLT7HGpUWBTiBNZGOlvf9si/+8+WCALoBI2naAvtcqgS4nkBESm/NnV/Pka9lG0iI95350DT
ASa3xc3+uQZyllCx5fWfPabU6797M7f9Lp7Me+9wgqvilLqxLBq9epTDZgQel1ix3zyI7jt1yYEy
ERGCSCC9ziC9hTDQrY1zkQerd7mvIOUeRrTcd8xGSYH62On0QL1KIQIerW74zIE4B/E1YNVE9XnU
vrBNNh4MoicWpOhg1WFhs0fIaghjNU6C/i/1z0EKNCJlKdGFkiMy9jybYlBz34TRVx09NFhvC7P9
KhAmbk8x/WIrvayALt/mUw3UG7ssly5KG3Js7LXHWtBSeB3pUW5MDOHAPEGO+EYc9FJ4HKXpXKMJ
Oo7Fr+p7cFYYzquNBm0Fj8VVQQ2NoWvPXpQWHdd7WJs62+/OudnIPNBiaKcyvzMd/Uzl9J3gEO3U
skTiWbIu6VTTEfYpj2H0aSXz4pXMzRfd7gim4CHMJodlG/y3O+XPlNsBuO6rKoN9Jwyj871wSy6v
kKwfFc4cXRYU3XdipUOOQkFNQIFyZ+mSsLlVP2PoIN+UyGPzfGTWrHWNK9lhvvPCIE9rJoFrWDzm
t5YkXnbHKqVNxJp8FYZpihsvgpGdEJNK0EAOIkiDpG2xxv6P2yPKBnLIt/AnYAhP7JHddjF4/zzY
y88uhkHBOeQmacQVhaNS6n8/xiEiP/WMAV/CumPOIAaOdh1FHIeQ8MvAOLrR2X3lQsBkOva9Azn+
O86xrmkakY6HnQnbWFN0MzO4eCTYrsebdqccJ0CFe8xPS91YDnLdQhBCL3Vb9CDWLyF6lo/mmoKb
PumB33lrxaOdsi/2vvceQ990qUla0P6TGEojNTVldBU4bAI9w7uC94JU9JDQno5iVclICXKHwSCq
2WgXsc3RBPna476l2vxdd6DOsBi2nywCm7Cvn6JiQ7iU5/CH2o7PkyHU2D3IntWFcViGRpGWcZ+N
HK7C3KryG861CuXnAR8ymM002bBDG7kB0d2PCFubZg9LsdU4OQzel5GlAgAQ9vFBl2IO9szPmF6m
bcAunoN/BvAWi1A24ei4dVil37KEUfdlm/S2RRBczCXgfCwz0BdjdqN+W8YjIxUnZQDO+GIR/Q1+
Zkutg1IsrvCk5LMe8EX5/IjIUJ/kfBDGboADkmLNksHcIm9rM8idYf/djuZRwIOSrmEUG1g4OkoH
RMnh9SzUWsMNzqYmpds9dnsH1Ge9b/VA3Wd1i3Rj+JE+fGD5nVWSavGw0BZzj/znHveyL6djAanc
qnTd8XjosGFeaco5pdKOKetugQGzoqkxoglHX/hpaQTwMk4pPtQSzTao7S94SAFE2If9XgjiYjLm
2LUpA/O6sZ2OOp8nZrDJQ92cueF88tT18Z7s53JEHPxDjgviwCaeSUrzUDDapIYIIp/Wwm0Q8qsH
rwTrLUAq9ZW0qc+9/2mXY8zKpb9pNQkr8ZJ1l5LKsCmsE/y7CpTAwS4aORcshlIOHbfVKWD/LKnT
erJwrCYZvIENmN05EhcqeyLYExWQ07WKH1Gtw3fY2JW5Ga6reRjcy3oyC7F+Q2ztZipScgDXOEhg
P3o454Fe7KZ4Au4QkOFH5oBeTdgy2nlcUJI3XNEHG5Fu5Isywb5NpLzAt+5FvEZGaHiBBwsY6/hT
bRT/p2JPE6K9mH2J9wmEdxwJfxUZm9oyqL9xdOIOohF9md7f9Iojrb18m/XTQKs329yiUOgnh8tf
EsiQBvMs0gwc2wjtmZdFiywQvYAoL+aVyIxkG3vTLg/5PCx5e1lXEFJnGpPg8+sPlfY/ZwNvvuD+
rWxTrgwpsaITmbXSH+feqf8Yb0JxILkJTNXFwTkGhzX7Rw5PlBaC/rIyq8vyRnbhKUVHPJzHtpdn
KZEWK6/oQKH8MPBUTdYTmONMpU/CF2f+d4Udqb/BBhg2QAgm159KQavvXwchAAtHx3nODIIcxu3F
Tpv4S4ODucXBy9X/yimKEQcytAyOyW2SWj3UjX+hoYOlQduCGM15LsRHY9vnTcVmaKdFeBM0YQhF
m8RykZzT/f0vWolLLcVQ/qz/Pnyw5MNuGH+XOIx4qQLHf7ndatjkwZnhmTMxrYvdXhqg/9WRkuDU
HEkwep9AAK55ZTyYPUseSR+7r+pVRU3L5+JjP61UwyDsYINx+PWuxRHMiMt0u7K47TEtZ2aJEuRc
wYfCYQwnyRWcnQOlVpxKISd9/t67NPkTcveautj1x9MisxyUFb2DkP3ewj5D7ZPGydh9u55tUC43
pXVA4UX1pz00dOF8Nzhjuk3ueQmUcvsQTzMHIA3UeSiqKPKpZVivOktHQWQ7AT0xbHC5BE4SlG+b
92FheARA29vzKux4Dp67zFQQVuc4ylTKYXjEdLW0JNET8YyUXPfxVARnpBHE41gkiUvr/YJHVeos
H/Xf+eEdxB6eDpO2APxJ1aAmnSLm/RBbETLsQafPkuE8Cg69sv3bmFlrjUEAB5sk47GdHD8/Xz5Y
GOxeb8nx+bfxC13PM5v2Z62maZc3WayU0F5AyXSnrBf84Q4hqA5tUG00XioJfkf9WpHcY8vsNwIz
Eepg46EguohKJlOmGl5KjANHXuBoMkC/HoOo4R3a1rIjYcuMfAFKrME0DvDHvEaVv1vSV2fC3dJt
cWDwn+PONSkPRiyOQ/f7nacVrfdIhTULnWcZEytkDi6KhUkzPLTdsXug/9JouLb6LlPf2gN0s7k2
5L9dfoDiXdKvjIDNV/9kVzH3IrH1fGeVo+mOx1DbVTYJDS3dBc/uJZlwrwBrmuXMZTmcmn60R+Bs
5chLaqi+amxFI9rzKXAeECQCDX87zrHlXXKRAqEXODopC2xcCHkIiSdSu/1Qjb9Falo7TYez1I9y
TMkdkW137WWh4MLA+HXhwcnN3bhCYkmQGS7yHFrXnTFBOTI6FO2g9lRKLXH7rYyaRJorM7ZtZse5
Z36CF/BO1u+vuXZ8iVSrSTwWgefnYbGPN2zZvXTCRjUbjw3jEhQMdBWKEVb7cgTCuRWdWQUF+mWf
mwYgp6ls0WgeDkRMxiENuxfL1Naz1VMGQ8oi8NDIitxwT5jLpunntk9bVi8Uc0lU43rqLsPPoY8m
X24ITLw5LXS7EpOAnSOq6UdtVziX63W2mMTJVpEQSuoDyEw372fQKQry1JGAMGGNPB6OoKJX6CGk
3JDTglwmljsm7BLu6Btl5wsqsgVluFcNm7coCkRWsWRzguOOyqqJa7pxkJBhYmA29QxJvJcbTucm
i2mQ7+quYUUZWrK5Lt4rVvb4klfBpNyz4r2XVkInOAvqTDHC2FhOmASluPqRvXDy5a31TFhy6A6H
yS7ADNIVJ3as34uFpuWBC/13lNAh4R5bXvdXd+AkY9iD8Hq7HB4Dh9Mr0ovuKdnlsCyxvMKsoU65
PvmzY0cJjqT3O2RfILDyhn8QOnvdJd5REbOoP/kZeHHYy4xNdH3uvw9MPChn0ywfhDi3hm+wYzTB
Y99ZLdRyFF3hb4jE+xjH8FE7qfJyAvmodx3Jkmus+P/46jHn1NbS33z6kiGaMDbn6VQFGih3Gk0f
BWg9UUWO+O6mTquIultbCVdLNQthL9rHZbfuArkKoWFme+P7vUAqz28vj4lMr3yLwT+DmOSBKMjH
vQuG3C5ifJA8fXeJSwYAbNPMs7u7KfaWELAXJEW6gq96kSTCHXgADYc+ekd5JKDAfYupOoptY2l+
ezN/k/Q5ksyXmbfgK44u4fbijbgKnnjR0yqi233JXkyuQA1KY8J4kFRrPzHUiZ2zaVe/ujqcMWmh
Lqf/OaooI/Cz2oHxReysxZAjhkyO13t5dS1vhObpCyOKkEE6sHwsHPbYwhi9RIvVVQSj0efclSUv
CsqmyRuc48sLQ2hrDIXrVPnuCqWRvBINj/q0il2o4ZPk38e0D9l46ML4i6hxS5+9VRmxzso2oxXi
knCUpdJtoxuQIZ2S/YZmCGd0S3RTMaeWhu53Xh1+xuAtns7GPYB0RUrd6ZV3L5IeFX2d3qLOWARe
LGt/HB9gPIYGOqKzwVsvsLHyTz9s0dqkQYIsOG74vxnt3K5ZdjoK+ugmtz7HIqCmCjbpug6vEb4v
hyGjui3adacFKuCAfiS7t3WejLLfXyDy5iwWcFlkQB/wa4YCg9l7j0C/HXO1SDRK6H38xLil5sGt
N7HhHY+l4SYN4I+MdQZ7cyAo0A9SrmFg2/OPiX5Dk2nARAl13SmyX04WZwBs1jEDDQAIthp/5eoE
gyMyzioVd3moRvCK1EYSKiN+O2CrTk+9I2TkZ1BaAgTlnsRl4Ii+ondW+CYInI4ybaZ2g3wPENDf
LIIKLkDe8f0cbgiSa9muE8WsBPHDeKrLSjnmfeBZYUDp+iqNGzFcTj9JReVMVjZlTTWL3HE19u+a
Zf7RtCLA5ekoPmes0xBbKJBVeOLUVkjGwB245jZh34z2+FzRR1RJnp7terW2zETV1HZNl4Pys1A1
dgGxyOYQZ7e1yUoZIav+sCDuLsKFcVuWiL3hr4R3+WI23GUwBqe/frZks1R7LYbI3ZhHMKesuGgG
XbH1eRfNp6pOevqupGbBdUdkjO01fJV6GV1mIl7FwAI4P3xWb4jniO+2MzlxpUdibZZdhS8xkmLN
UD30K+1joDeWnssFks0OYOakqxFQCKrr8th81qLKasIn8Lh/OnMVvUzATFUXdeYUqG1vN0uIAJMG
g9H6e1wphI15PF4sy7WK+0/Dy1LreepU6RrrF5VtPWvvEFRPmUFPxcRR0fTSjxknX2w1+lFFREbO
LtvTJ7qqu5SSx6kbIJWvX7Wvlc+/WAIc/m2T7Diqw80rZVXYRm/FkFbLDr29dygBFQqdQIjHTYck
bsdojrgPD5/Xd2Ta4h0rBUGXkM5shYiILPHOFRuKNPU8ap8o6+yZnm3wtIkDuW9CMgVO3NokiLGA
sNckyJ9cf79WGESi0qYVghnZ+mGazAis4xcWzDBcKZv+Z4C4YheGhrAXZ8m06dCtlfrmpBDZ1tak
Rcad6vtAdSuxhXYeU1LpqTJU1dIfcBMWXxS+ZTFX0A4O7klO9N3EJdRly3VRWt+/1dqjnhvdMdR6
L+gLgge9zj15T95v4gh0ptbxJIJ10tzVTHFpN6YTImjymw2H9UAxZ78I2X/hRLKyzE2Gb7S+DT1m
GRMpWqg4z5YeY0TAD+SF7DXh6oWVxZ3PS8iLFjayQ+sYU4oaIlJuqOoVtk0toTPHXFFN3Li3MUaL
a89oGQh0WRTHpuK/htNYzEjFRQQZudgGT6lVy0kFPpkqFkaLL2yhWUEsQJkWiUucl5tzLJcD4sQh
KfSRSc8OAAoZRUTh7mpC2bJ0jD0mPKt6A5LG9K8C04davJCN881G41milBbVpkHz2kq7UZ8by0dj
QcBEYVYNmGPW4qCOUgOIqIFFzevJLneXWFT+mFxYCCwzMxsMjKba1t9VxozCfQZ/Xi12pPBTa0uG
eBBMLLVp/4YEOlfBx8WZwrruf8CeVKFMcwQNPGK4CmD3RyZKJYvRizp1xdvVeuc7UcSsEPI6TLzW
pXTjKvjswLgTXEhmii0BzwZbAoQ7+qEY2vZL+St7usPlHB+IUGFZRX36yKBHaP3b0cidpn3fh01i
REaVLgmP1sywHlVhzZZhTKyOkObfBte4bqlq8+OeAWpm5Ujnnxs5WNvHZCzXP10FkhcvfG3rIu7d
Wa4V79ttiYnV75BDHINFoe7RIJCxiGChnJhJ+6oi1IKlhqHnEq5usHjCVBO1koN49YMoF0tMjb5U
izRO86iRkO4iGDx2tUXPPcQoqUgB5uEN7G/MxtMXLcbh7qRWd9zvW0grSNYGbHXfEpKw4dUcfYn0
UPCZ+vz4f11fwUlpazRMib3MrUGZeNPSG8y25AENk24090yFNv0LRPlfvqRnz2161M7w28CN+RIE
RSwIEAIWQ+JI/4kFg78Ig7e2gaEj4YM6ws28HVSKN4jxUoV3g0PB1PGP+izvHveAABUcmaiB+1+q
6cD+zix2aJlzwexiULQuYqzrFPN2hwGzikqT8cgwbZ1Yd8e+vbhAVnYjpSsUSZfjaL/7WWEwUBvB
EkQ1C+kKkwaKQ0DavPN3M5ueBcBtBSJ7YeMe3/La0XpuQiAH2cDtEjECitAFnYcWo5uMhA0RjQSe
LV00SzPlzlszhJoJmvFO9P/PC8tdgHrhHtjT4TC8wvrkGxDwIPpTxmdX+dTMeXjnCAxFeTp2fiii
U9uGHgbwxioHToON2x/biGf1a+d5W3W46m0vG+2OpvIHFPCCXReQgfcCT9//oRFeV6mhnqNZWatw
k3irmHloCDISS2LqurN9q1Ixey4/qZW79Gda2dUr06qbED4mYTnlNpqz6V3LzHVm/yhyFy6XRXcs
oxU95+m/QN3bo/t/sN8pc4/OCwopxSklH9jcamap4KPQ8UhSQq51vPD1N3Q/9883jrD63bdsTfcW
3BHWm4pY66qzV/27BuDnVxhRGBhfRsDhmDwkRCMx4lffG2+8EMnRBjot4/zxWYG4k3sSsWOtdz01
3OpqlkNg3yN/JC44YjKRjsbXhj8ay3W9iOdQtrhEr0OG7N/WqA8LQ7AhSZlfd5WTAtg+OD2bMJ0z
Y7HlFk3g8ErQrOi8mXLovrKbI9nGlVSZOKqM0Z8gG3ZYDHLmwPhZ+eA3VKZ7ifJph2zouSTJGvA8
IAtZmovJKcUpxwv3mZtRJdgo4kEc0oTITCvUIjxThmoYm+Okj+a07iTAMsM2HIEE333el5FFdw2X
C6ie1Gcl7QmP+cLgWX/lVVEn+LhSH9HqM1cTXrnI7kJG9mEwF5y7NX65sJaXy8xB8VQBeK4bBPSf
D/+6OITFloQTlhzThxIukqRN+AzdUJ+r3j3xX0rPoj32meriw6PEuLOuKjWj6GS8AB3F930gbL1i
bmBY3qIpWn6/OG0dethZCn/kakARkfiGAO8yMVXViZ+T4Ekbs5duSAEcPUXO3lmZ1+7t3YGVrooW
yjY/ilVX7FHyCMvtnBvSjuTimFXdeY1z06CB0K4MpaeBHFhMf9vd7Sfv1hJ0KtFykhGBK9c/jPag
KfK4chNmd2N7+zV8+lsYZR+1jRsL2eZnuorxncKpVfMOmdPyTHZ/xdQh3i4aP0GqQ9TsfTBf/AjC
U2crd5VqCEx26Z0tW0/ox38dtVDwkIa2Wlr5DSRjqzFfhABIfzSRCDzSaYBhn8BBWmnLvjJHyU88
M9ERvqstvxAUWGGUROGtoIZXKTdp0eNVfppviYyecq06jK9Su9bbtfgMiCrCUbYUT27LqrNmC9Jw
b/o4zZFsM07Pxr++pdGaJhjkmNfafVQVwmxJEcvyrQnejG3yXwySFLQbIciYLyQE9ST4ANYzji07
aKnVxYcHiI5TVFMz1JVbNvv2+JfFqnNnFgFPNi+g/7L8f/y83uezCtKPrwMcgsLFdFtyNTB3UTk5
hHYmyN/kra+Qzj8716d9zYI9BUT4QxgA2uKHfT9naYAzmclBalOigeipk0r75wwatGthZuV7hDob
Ynstt0et1j/BaFqrcxo2iXFoxdiO0B0R73jam774avl6thGIiI0O8SLFO+Z7AtF9bZFb9Ob9mbLS
cgfqYZ+1njBTsDP++VyZyoZvjKDF87M2/jenT2Cpqc6Id69dcJIGJQO5xPXccVO5dnTWc+6e7dIQ
fTJ5K/u6fSq9PxjqLzSdlFcRoR+9KoLPy6p9x0EDE5QFK0OwPdHnrXE/Y3YFy3qfRRCV7g7ESpEy
KJibKJzNuH3uPA8f7KAfrlVrWfu4hrKaMU5FGE1ONb7VAcElM4UZf4e7Vw9o0MIa3TBfSkqukjr1
coLt2rde5N1Vm29k6M7jn4XynZ2LjRX9GsH8EH93FWNBw6BYKOHYk2AwXo8T5eKS83QJvw34KsDo
xCaxqVGXvV64Q+umWNavZfA6RAkifdDdeO0FD9BB3TM0wg8sDFhNaNXVx1M4vzFUUsJs9ImhPumx
asrzFFjuKODJ56Tp96E/qnQ+ZsnbbwC2UIq9Rv1yy11JPjZ2NhyjA+MnRF8Al3rJkAalJ4XqYRg8
TbsWzf+txX+s0FqrVEBN6s1e7k1XMutk8lYX4l4Or+IlX8JXIG4ssoE/4iTIfc8UW7M7l3DsIoMQ
hS7Fy8XcPsVmgPaTk5k+iY8bY3V3d3Ehw4w6O645HjLaPEklQV1UJuHjs6W6FeCyO+RfaAPgOxRA
Rr34AHyhSw8jU31ASsX6R6gn2ym46rhsxkVp8CrWIBXLMhCwCvYV/pLr9Vyo7RLLwdACZ/86fo+a
5bkFu+em2sD314XLf62j01EXKCBPFrRfBAAfpZGGzrxM08sTfGyNJKEl4IrAPe4hWs4CtPrFQ29s
yDiGFbwvu+uL3d0rJSf6HdRDodYJaO5F73qdsL/nvwEwHLk3z3qgTw0gerI4wai29fhIAyet//+E
zDb3soSk9gKKUPwS9IH01NktZduVYFVyW1RrVqMGwZ/ByaUDBTvf/1y74APhddiU5wT36/+ftVyH
fUTV1o7rg+LSiS0wa4xsmB5dCo11KXJMT1aBnmZ94Izzw4VkhjI4j816/Yk5KgdYtU7IR8A+YakG
s7wFbYf8j/vMAkP+aFQ+PyHwxVDWoEF1wu96TlYvbRcdgqiurK6zAnnzELqyCWxBO3UzBf1fZIIJ
u/8Sfp3/i0hmF3excCvNYjmyxKjsT7ayKdI8pxlCwOZmBjCo8oONrXbLTKNXvuYPluxQThTZAY9G
2k9kTsv0pMrsvfTe9preE7AzDJEBI7vqdgKPY5nztWM8SrzOCNj891X/eeIQZ6tAPDcn8RCURayf
1g+tkipzvumWr6hWCQXvLJ4ZM7OPm2mZWuYjm/SItH6cSPS73G+kGgvQaST/cKBykMNZ7V87Qpqk
+EZ8w6Hnh5SQpnBBiUOYOzXa5Jk5Ioxi8bi1BlP/Mo6C6XRm0f14X1SSIdyHg98Lu/is4XxSvtTY
nbXsGG5JqsPu1NA2AxSRFO+/crFdBLOlR4mx/vOCnGb7GmwTQPKrqNUWeaOmW9j4AS2Qtci9BTg2
GRcZe9e701iPUmCxxwEDkUZaDt/DytLVnIf0eiIdTMy+5FmU9k5lZJS9GCNAk0/TmVRGWei75Zdq
nfFG4iIfU4+icun3PhErg7M5rzdThDKTKApMSTlWSmlFbOSZ+2YxVkMw8COszd7rkX3agFneUxFo
ydlLcLIsUDgPPCHQzdkZvPO9Jg+tFScif/tS42bKmMr2UjD1TuPwvkiMxGWRjBZ6lAieJbjOL7OP
YX2V5xnQQh5raZrbYeFnOuBg/TIxqgTBTVUmAGAVrgotDsQE1MqKqY2hyljtD8nAEbSNADoAQCBo
gJiTwxFL/rZ+xOn4xptZFDLiJnQYuI1H0tolKjuEI6/M3aE0/g3oBPXTA6Rpnm4a4tCCGmtPbKrx
f0WEV8kx8ZNPmRAhC3+4x4caJAK5d7Fp+/lAvg/WFxctSO290kajlr7LwMiraYJcBo5C0CbMpS0D
FOHLm4yUJmWlM+XHxaU7KO1E0M3JAzTq4aapeGMJz65Hms0dMlwb3Pak/uK+dsHFGaBJWoAB8Lfn
8mMOfT6kWDuZDU8AKfId+mbhfI7FVFjtSQj/eYb64mTpKRZbhf+K8n5fnx7itU8lLvrNRgzBlrsa
Bf3b95CIHBPw4Kh3ILbFA6cCYzVurEZz7dXV1kNDuiGWnlImoIPviLn5fWSWDSenYtcfcJWxivMD
58KOzhaOQuA9YNVIfYLSPTBC7WypL/mb4NvYO4zEUWf3AxoA7KVzgpGV/YkFzmnsCO0xiQMXQsQ3
NtnsUhlRWDwGhYTIFrNucpjiXXQ9ObpXsamGkIfkE6BEYfEZKtH0uZh7C2SXKbVtz+owCI18t+cL
L7DSpLaSsXqxiZEMYvZ06j8yvdAchPLpRogqMVcRKBtbd7wOmuGpDvpZVnW9lQiMC/Kvp+yy/fh2
x5ahBI0QaFIWT0jR0tz0gL1yoP1WOHfDkkpUQGZGb1NEGJ98mYF98YYdnaDoVpGZwf7+4eOBFspu
BiuCQ2QjoTJJPZZYwuKoUriEoGqEUaf3o049g4otL93n7YyVHM3WxombXHFnJVkbzyErLKTnAgse
aT5G3tqGsQF4If7YULirSueAKQFkJpIJrhQXmQeRNYQQckAayaG6O6WhPF5BGY3qCYmaQKWvraS/
GbsL3hmZgdklNXNkvP6Vbxo+m8GeEncTAju8aq1Iv1dls/mziquWuYwnrqFnI0H8/nDnOTIXpAIR
Aen/b+sK/CxWWwQyw2Tql0jhupGmf09qYJQ0i30LBwQ5hbXGzwIOdWQZnfHhly4qvd0cEpwfZwin
ESVYIGpEt8P39818Y0s1vD7JrJgMNhazP/tkUDxPakCX6Vv0U3pBBLH4nzcbrllvuKspQruQVQHY
I3AfDJuesKb5lxNBIxlsc2ekqH2Qitr7sOkR0RRLftS9tqIDmZDagHcj8/VTggFthj7BJS4B2aNt
uQW/fLl6kpIulkv4QwQICF4nRfqhTAD6DEOaazBOLf1xzokcYfglxMjukbxw799hdwerfXdZ4mcD
cfAedHMbM13AIo0NZQaLhrCJk8YJHVjs0T4R6OaqnFSfjhFp3ZV2ZXmOv6+skRPU7Bs89Y6o4jdr
xF4Fi3Ss7St1NxLxduhGGKjmvZudW3XcQk5sjRbuZzx+XUsuNoF8p64oMPCSz7ZCr9W/GDRVyNSu
ABWQ5zqgDdKQEKAypr/q1wVRIERx1gq1nrVOjTdpChfHjkyg91akYn0ki4f92l8RGEGwQS2idjuQ
VfdfBGON8LpxOhXOh02SbMb+4Dq5qrcdiBWf8xt6Mucs/AmJQE8QqVnJbb0YPz3A0LEQsZPXLBjx
Qg/R9KmXDPBiyIB1CUcSSmeUniZgjY4dZCDsFZw6TclhbSNsrG3r9T62iLarSXeHZpz+f/UKc306
TN/ipZXKXzTlq9yys2ShWUYb2fQVNHX+GLcb8aPgm7WKSchv595bBkOFw6ukKSmAOCDIAZxwauQ5
a6Xujzf4HrVMv/UAkviX84bBgqINooMssJSEvGRTeVZ14Y3txnQjIBNdzlNsJ2OaD/SSjHK52Ipa
Lp2JYC6c5H7AuUa3aPbZ9SPIzIRSXbi8K8jzKG87ieEHqnwvg7h689XWZa3H7v5G6IdGTnyl7Wdd
aIhM7uJEaR77hwwksfMTjZy+PrWEmSBTxYUw7T7/yoVV3TQqX0b3bJ7ed+TXh3USopItMAYAPsMv
+aFeXWJasKSiMrlxcV71wT2Fv/37lYzV9e7W2abDtEYoe1309chc+B7oQC7zE+svW2wFmwQqquU6
lYafX3/Y68P1PDq6mymLn5fQWfcR5DInQhsPoRkpt1fCeBPf8NvKIVA32UX19CCOpmXlEck4AvRR
4kfGjGPCrisGHkCKAwRS1FP0eaxReUaHrX1gBIJ7XKJ3uKzhhJ1m+P5tCuCQvjpHde3UQyokrweW
nqF8x8N2eF5bwpV+YMH+tGzNGafxfk2ZkUOtIe4XYy9bjZkVBjiW1M6GqyGKDfNP+qKZDKQOZBWB
oXYEp5+AZXCBXb+RByolRd5HiqtM4DZ25KHO53QbBOnItk7B24oE1+aE6ibQMehqWxmfZbfOUGV7
pcrRZbHfKeX0THNyF9s25lDz3BapGhh9cy6zhSWtbIACE9SSem+P87g1D92AaPUTNq6pAmJ6j2kR
Mk72SIpqhGgMCKafdu/vIcw6uDCkjyn44MHL36hrpCfs0IhDRsgduI2Q0Va67SmTmWd3UIVZ5sin
2o7XmljmZ/cjnHTcVHeqihJfnc87YkOcp19Oc7FFn/NacZDymJHUiO55KKdkflch4XetxNuKtNqk
KxXsOTCxotQHngb6iTffim+fMbl2qic6P+cUrZ6Ecl8Wob1SSGWNpf/2kiV+ocdBGVt9QtK1j/9W
J601NxbPhJOsOpWfsAByh3c5Fjb5beR5rLVrJK4RD5LJ/B1uA1FuHVbT5W8MrYqfAd8QlgcI0s1H
XXr+hQIIroCvGxnB0QqsgPTFRaws3gmZS1pm4nKQVLkZUTOvothl0H81lMlrHPWCGmrDZoLuwS96
wegkd6hK1LGr0f8VoqkEPetWOmKDMuf5SR9GpBCjrLaXG40yQUbSR63gq24bLlPM4gcoe/qVWSob
+ShMEmKn7ZYubsxE5lUi5Sf59ObUak3BuMT7mnjnXQiEY37W9sBHoGMks/gW+L9P5tApHVvBuH2t
cyqLIFtjSigBnLhO4CyFMfskqyENJlYtGNl3i63S86dKlfWlGRXqm6syqUcdGTtkUKjCLss5roOs
bc2eFYJB0/lPKXyF1QnJGAdfcwf5vo0UiDylHf+mCYM9rujuqK0uJ51RzUHhcAIXRbFoyGCutty0
1bMH46vhlwmkuT61ufX5u1boOscFjEQ7of3atFEv7XNJL9E5nPwyjPqTgVGDXUza3F8WUhR6QZcq
e8oasrfXnCeLm4cbqpaRB8VpEfHscrskKyBmtb+2FFFq5/Y5ZuiWMlsxchMznFsDmrLYuPwQbUm8
DEXSNYjXgx/mLqBq5IzfKR9TfEWh1rTBLbUCkmfCy6UhBlw30i6a+XOundcEQDXpZpJuc2Nhocv3
3eYi2yvgm1ghXVroiq5mJ24ZsAzeFA0m6nbiYM/eu3vzrjQ01iS+ZAhqwT6GCD/Fh1sVcbS8BFB8
wbdFCm76+2B8cE3mSBS6crziaBHaUMgxJgnuO6u2EUy/KzS5SH7EmK6hJ9aa8FCAolYTOYRhzDp+
Laxk9/gRPZ+WcN2ewPhLJHabr2cFyRs9O8WOeqYdkLjPHdMTLHTMw0y1yyIKjHRRxnR4TgzaPNAf
kurG4H1ZijM5YfLHqX3t8oFXV1+yQI69TEYj0X7RnS4yjRfOYf6PawRpZ27cpS2RX2HIRlfRSVUM
65OoHrLx0xNW6653mkY8JnNEqw9ZYEcYDVnoblZWlMtLO7RBVtxBeY8Z7GCJMrFO0V4iTuFNsAuG
/1ApWdF2jqOnUhWO+OovjTR+E2CphjH4dm+bafs2FHNDtfkAFI14F+bt5MC5Gl9B759nZg31GdJo
ybZ3HRojGYYPNzs/H73mELAA+4RxsfcJlsEXTY/0VcaHCOpH83GoYnxAgmMSQ/16SMaXYVv3BjpQ
32oAADthvDmmGseuM2JjWdmrqtZsXvmOchmYLxctjJOOLe4cSXJw8iM7VnzAzy5idxrwBqFzH811
SEdgdAglinGJfnF2yCNqPWXb6/LXlYEC0KjRlNR2Ga1ILHum4lx6taOx0fqMlke8EKWKnkFOEQn3
buB2tXhWBM4imI79LgWzj8qrmCrIIKEMQnlhk1iUXCMZb5/3Xi9HVu+RF/WkwQCxgr10HDSlaUyN
U7KT0iWTreGge+JDZOjuqZeXvZ+cNVQE46o3sXoGpIty+HH4knv21t5eAxzxQzJMf1l3ZCy2ZnA1
NgnCDvW2cPi0E6fnw95UkOCrWJtj/N+KJy5yH9/2v2dqcgiYfdPKEoQFGiFS39db6Cyk8AvxyvPB
Qm8Q+8IAyiYUmLrmL8AvbOcH7nbmga8mVWyy9Jl+5bAK5oDikI4jteNsUKaBZkVStJIabbKmGHJf
PwMRT8v6jSvaPz1GFcmWJVhEBKdC4pIYS+K+QY/khIInXBYXNSAmBYj+w9E1IcrwB+q6HUvfuXxt
qiBDk85Vz+aYXMcFEqCEttE7DAYpHfOds56qdQVz3mrJaC4Z+QkAnoNnWh079EE4kReWKvkTwhnP
vaSzrwfPV2ZJVZPFELMbUDu+8kzDxv6AvNCRYcTPGuGhoqnQyS28lJ57v+vOljfBkd9hIWZe1Dy8
QPCdarNZ+1hdmSK3/pJvx+yqstjFHSCqbfWmLYHLhn9mSemAUCppX/+Z1FHxnj+2zTucV1syAhQn
D0lYb/+1SyEw6IAhEdkngpLPZg5m0QC3fLkZb4cSYqxhfU6G2a3scAtZIYdi1KzpLgMfbTmHKJ5A
CnsA22zVV2x4vdIbW44bjZuF3ueOY89n51yF+tWRwupVxrU/DFrLBWXJNiynSAhJIC4JtUgxx9hL
q2FetmWMj04RJzeQF990gE7+MRiI3PIv/b0izltHLHaC1xnb1MVMkeCNzLMxULAf4jnbk8ILDutc
AG8wMeUHoZJ344GJjXYoIHKeIc0spP4E6mgbQJ6zcird2YttU4/NLCPh0EC8QHgpzKVB2RWlsDXH
aKaSdRpSaEDDyfFHkbU/U34RBdyunCcx9NnIGF/Y3l1X2Ef9aE2516RBbV6RHZMH8Wep9aUY+gNG
qVn8soIcRPVqoRD0RA/77+t7B7HT+YdgQlb9k8VlkOu3dpocBH+WJtrY+8WE3YBzZS/91P0Yvdh2
igPE/EPu5UXmh9N3NyYbTcKDr2iuadOrCXWBJySF9pIb8r8+oWguOeCpRHmaJW+IwlVtuhaWBtZy
gEo95rozSJ7X7dj+KCN5Ka9mWqC2w7BKqCFO62/f2Y7Yw/kc8uMX5Xg9FEHd0Vwcr1Guv1YTscqr
E+TfINq6F6ZXNhnxyqRkjRIWVs5fGyIkkED9FGQUHpu5ryT75tsedlCPxliI1o/Ykmqq4ookGAtM
k3v5tqr0eWw9O/BbHaUtmnYni3hTQF10DyW4SiZmn3EHBNVUa/YbwKYCpkFp6YZvw9ECJEPajtb2
mEhjuR/lwxPepw9CxsrvBXxclpof+vxDbDrVgGCeGH9HJ88dOCSw5cZ9c913XpMWlXfHWHY7Ge9u
RpAYCNiZ79/VWBoYU4+7rL7O78T5BEu+MeJ13XOoWgYzt9om/tAQ9Kd8d2c5++Q3aHRTtW/6Y230
QvWI7jofc1uV7cQnIx5gzmndBVIJNTmFfwwQlAJFxqPvL8IPSBQvQ04XMOBMYPRyyWcqg72Z3BGk
T4o+nfsTm3zlEDJM+SvUipGjSfGNMmujcwiywgtJPvrAH0Co5QK/c6xANxn9RRDG4m8ilHLDLZ15
M1gn94HM6VEYyt4NMIgNoqsdM0z85q0U3jJaQ4u9Uww1QYbsnpz5ODHR4Tihv2/ej98E6FaQZvD0
gYQdTSv0mMrhdrqJ4QOVI/mmFR8elPzqa4j+Bg4m/1LuOcPPqWTprt9EoP0IuwCrvhhiKuNWXLCH
WxCX6NTPycI5vofwnYD0X57rHKwCxtnnGGXS/Jf5QNZkueHLOlsy8KYBtMDwadmFi4aBMpeRii5p
IeBIi4BI5QBprqeVJ6bf26Jc8CTIki9wRPRTh6d5f1A65H3ErtZtWmhDju1t7l2mzp7HVBG0cp5u
LKXk9zeLWoHXdGYkkUXOxcw5wV2npVTpf4DqnYCkOKHijP8nPOorhCBsj78e7kKsiXmZ/G7gvrwa
J99S0uyGjjA2r7YGdsmjD18t7UM2TZVvNBuH5hkf3X6qjD9TGVMZx5s8swoqCC02jdqN861EUtgA
64XAl1WomvL0NiYrKg8FLzGmPwtdj8DSt35hX7qkWgwO0wN7Upn5brfyCNGdHYDuCx2A7IC2zoGl
X+Du22Dw1twId/FBkYmQRW/ppYTOKoQ9zhRyjmuhRF/CCDhBaWDT06AHuhpevVphmf2fQOo/FbFC
u7TN0x23/IL7Lt7Rfsf65OBHuyce7PmmQmza4+FP1hdwEby7HA01JWCGY7Iji53JxCIrWF620uoB
yJlV0r5w+9bkWO/EQKUteXS0cTdvPFGtkZ8E0nUNDOLXuuExaaI8Tx2B+8+qqSvQVnswCAIwnS4i
uDwikUHyOFI0jPYKEKcgxODrNrkr/Pd2GhD33Qm/i73NUFrBjJRr/PyhthEwaQMsE7hWV2/jWgAM
ZodmSRWO+WI/8JWj8nSvkFTnBZ15u7Q9yzo/56UdLLkRA7gtAYmbB4Fvl8E9sDKAlQJOyQn2OWfl
f8yoTDJtmvzsQwWJUL/CLmQzL/pBvuKf62BQHOswsqDPX/yY6gNGGNDyuQ5IQxiI7xZZRrVRDpSx
s/OY3AYUtVwsjRF0qsxqHmi8qU4B4PoTo6qzkqT24fQUK/pastsoWLw4AEXM9EQtsyHC9S7oM1fr
R58Raz+yy54Q/g2hl8wGpI9caFeGB4KcIgZALDAQltMowzk416svbPveFe/kB/kzKsZw+VszNnG6
ZobgODs1GtxjnedFybGByVgvtt7jUgYnAkrijJCUwzcinXs0mI47No7FmijAFIr3H2p58sUfl4Nf
tENzOmAsx0Q1o00nAgsEWoMXUhQqwzzYggbQCrOtUuNis58t+axUTRwFatHZqvpT4YuZAPfCUxI9
pPvOJGbiQ5H1qIRpRaNjV9KlIYdo9LqxsStuAKiPGbaowJLk90Uq5L7NIh45720m1RdmPGOOivpF
o3lfks/zHWcZ/EnN80MvUuBrDV8Ux7h0ng4OVHDBVV4A33WtKi+E9D79AVkKK8TIYugMsNGe1hfz
JXFLWiKMbn3XqevCiOl/agQEgX680uqjzfc8kPL/3xvVXGviR1vF92MMK4E2+yE6TsjnnZsQKL13
X6CVGaoPFY11eU63R4qNn+BY/LVqeTN0k0D+NiAsr1ucvXwz92PxYA4ucsjn3Mx802cM6HzKHUz7
sN8exE/6FNNLY3HoseKWqQpFIU79LfssOZ0iutu3uY+0vF7y5k23UdTPokkzofS643B+CH8lwAKG
Urai66NoHEvruMa3qg9fBSteR4Uu6Z9uCYgubhatT8DxmDnOHGlyk+NydB4mZzlt7rPe2SZczBKD
ifUSzZLjp94ZZ4qW2oAR/+vwp9T/30m9wySjP9cGfqnqqKRRV02h6sn/pmH5OjccPrltZGYFGYtP
h0SpfzEaguLv38KdF5kes2DOjH+6x3zQ0/y9yQ+aRggb5MDy98ZN88KDTSdeFTlG0L3bYn0v6Y+5
glnIog3dhbRGSzAtiaWWsXPqp81UroTy9yh8PDifkHDeym2zdgonINNjMsqae6mA6ncqjyqokMSA
j3/l68g7zfiklq6SkRpxpcep/KdYfulUuN1OX57W2HyPt+dwyZ1wVGtqTf+3D+70CWWvk5OlyU/J
ck5z0w2QfPXyy9aY0ZC/pXoumdd/vSNH5ASOrB9kytPYLFFDp3Lo8+tTj468uba40xz+2kwaoL7w
sbTHPAJ6Se/rxgGHJPnckl9+Po2mKmbds78D0p+WT1Pg7febBjs61tpQxBgtz3C2ObIq3qTM0Eel
ImC7rpz8vO1BTJO+FKGLCWyIwnxPb1y+sKHKAOezvKta9xZzHyooCGzidWnYtUAjjOHUU3tMJUSj
Jrs0W4fYrYeMsyq+w/cFuEYF1Tbi8ZwloUTOW/fzqW8cxL2rXj+pWWv8dHqN2cd/rl11zJmBuRLw
Xv9IVV4Z0iYyJtLwMnUsnHxMSuSkyB80QlHiZLZmcnqEanRpqVOD4E/0T9vQTJKJdiStcPEG+3Ie
ZEPSSL4Fr16JzL6mo0nDtI/s7m2ext2Vd9tNPuKlxWhyzo24d+TVCoL3cGTkDKNS0+yL9RCdjo+0
S68XyTn4vRNtFYhOxNR9sMdB9mG5WsyRSNstZ+pJEWpVImL5imE6ilqm6s02/CNuvRBqi5wN3s2K
WRgir15wIcNAyem90jcb4tP3th5EeXZRo1ND9l1TfbIMLZclCFM7do+Zm28N5T9Fup0yj88deSQx
Inv83ayTcwLh+N82JAV70UhMIR80TWvBsuDIDjLYZxamOQDcD9AH0hGDanNHqwW/+vDTWxVzMtRo
mZfu4IqocqZXRDaLa1ApDmrhVnkg1Ln5stuRcAK1bUhyXNHXMgURak7Rrw1rTBRqngX5P7WGV9oc
TIsCIjBJ3WtVmEGceLoPdJUlBAzH9ckmIrnxE7kO1TfBu2lEW2sZzkRNc4fK9CjBlU/GZrlglf1m
3hjLzvIUg0Qhz9dmY3WROM8CSRDgclQvBKc7sOiXfKHUQgzjMF++pc3AFeJd5hm8r10WmWr+q1ui
eZH8lXIp9/mnnGnw80OGmp2aPnv8JJZ1jvfQrNu5ymFp7/7j0heuBEXaJ3ngoLsb/kZtiM3EOsHc
0q1ZmCHWSwLcf2hb1kglCY/5+DVxagtV9BJgLMNp9DCO954j/1REis3uYeGQ8hEJXZniDSklEElh
oA24bbG6fCnCBfMLkInApCzSywtFjAcQ70y+866Mp4ux/brs0nvRu+BOmova0Y+Y2VEFQKG8dP7K
pMUTVkSJp4mi92MdaOS4CqTA4kZfjFOEgj2V5g/oBzmqOJOzqdbuSqBd5d6pIuHMrHhSmo7zjceh
vRSMOt3w1unHvAst/oKLLyQywGDGRHZAiQoHr92txFgiNQpsiPRqs+R5qipdI6ObZxtSwaREHGXf
cEpEuT76FXGPvYwqColwIWudZWg1VjLGN6VTO7MxT7A+62qPeuTgpOdAB6CpTiXeXWu7TeOZWHQy
LomGldGOZNgyCqxibsuo2SX7PutdcL1EKT6sge4lKA3vxTp9Bcweh+Y1QnCWt9HzBKxs4OMftxZk
lHIPbk9ZuCZTuHG5XTkyo0I+zE1BiXWgRxqIqrd1LEA/BertrDXizm9yIFntT0eZMgXW7XKGicU8
aaQ6+BKy2C8+f2ypLnH8keJdUMPQd9GrU87F4HsA+OrFTN/+lVKrE4HDOi3jRm5eMSCHM6tUao4k
yTSySuV49tWbU+cYWpEL18mZGGJ+dhOFx+VBOkFNm0tlezHajuvsUTEB2krxFGMVa3gLShbRRJ4u
9Gkg2woL0nAZ2yfwQ/GuqbBNoXUkWusnDZ0B9OqZc88lRWkjOE3ZoU+HttfRu2FmAzQozcqDRBmU
cDsH69/c8P2rkPOJLVB2IvQ5xGA5/BSwJq6kONku0lQIghTstTyTJY4rDBD8Z5m7niwFLP+21Fxv
aiT0LQ5E/ACIaB/dm02rNMnxDX9GzZ0enl615QJ3AnatN7J2XbYiY3UJTMfVYaXbsMVEWwi8ibLF
UKb29+/t9ylcOvqHCww7pwkMbEFdn5Xke6c+id62eYvaIHkdW5KYY0DcWFEbUuYqvd/JOCccW2So
QaxiTzLnIqFw1aK1nlZhagl7QdSjMPgdDjzMNdLAPkRy1qAytvXdc1xpikgrWmpPh252bxXD6djS
wNj65YaHdiyDwvbIFsjlWTRhDgS2tC10b0eIqh5NtDDyVqI3hGJoekumH7z+y1khDqZTYgddeDb6
AD8S4N7Mdn+l91qLxX5z+4G/QjB3uEktjztIpy8Ms2GG0lhTJBAqWX1ZSgx0q4LiJ7wYJHGUQZe+
THynQhv8D794lSF0iRmuupl3P7pBeaN1dOvFSVibXS4laHLlCwqprnv+N89aJ0I5l8p1no5oiRek
MqiTgZNa3hhj3ZwOZfXQ0KazCOkgWQkCr7qFfbjURErzP3VxL8ifslkmiP+kSwUb27EYjlpjC9ji
1QEeNeUiSGjtNVYjY91fUe1xq8sTr0O3OnF3ojuZjkXzvfYfNfYSeHWezcA420qlrJYFGwNJtlvO
VcSiY5/lCbvI5QNH26MJIjbbFvZ91cucGnMdIFy2bDx5R1e1+CKQGMQBRcWDR4ZkfrWklO0eioOC
kGY4IAGdP3XXP/u+o/PxWcIyyO4E46g7d4uJhNGh7OQ3XS/rHU8Apm2zjyBPmUuQVEHqO7DOMEpu
2H1nSd85UwboYhNxFgEwJ6pfl7Mw3J1kIljTARLKooPvmDJpgsCdCS6Soj0FkvVvucFxy5Ar7Twj
iDelvpmLhlCR1Y+l13MMHnIS2Epf4ReEyMG2szLsv0LdPvpSuH7T1zcDqOL8KoNqB/NhI7z1DzBI
DP8u40V3gBlNhqPNwpLFR48W1YG9uJ4NGIMov+Dy1jRNA2R0NYBYpzzMbWkYdv6n+BYwQ62mXTp7
o3jEKprVt3iKLNipko+bQBCdlemzVZOi04n2fiwg+sre85AWGXsiOJ1h6H0BJTB8P4zhz1v9ZSgA
0YFNrIIfFVwK2SoFvcSs2/2XMXuBQlzCvuwDAGW/mFot4494BqjHEl/iLgvwk6ebHCdj6MmGyR0u
BD+5GO3tr9epz8LdhQAG7qo/xxof77PXoC+CDvPGR20wM2JnM+KBHoFEyqO5mDkNq5HJ0PuYH19X
wzR3A+N8Mrlb70cLfP6+cqbi98LlZei9s164UJw68470De/ZHRiIymT4iv48HvgDRGoYBjZab0yH
lJuUGbsXclQYCw/e/iFymsdUZvdocyke1B0aeE3kDW8ELLoS7XCTcJmm3qD9/vr8M5OCT2YZMpht
tqOJtbJIXscwc0/xXWgnUgiNOVzNDGBdE9XeholiZPqSuQJ4XIdGeMLb7iQm/SSs2UgfoZ0KRnCL
hDecQ/OIlMzY+PNyxzAc7PJMSrBNEep93X9246P58R3qH83Memykfa70vo4bDAy0MmPiEq9Coxma
gDUSGgd8Rk5mcr6YikQBtjkF6InOL6WTuAyJM0j3QOYYp56Dn0l6ikH/l18SjI4P+Z9QvfRMetir
YUdEeE5fDNHmg546uxr0yd+g1iFopLOvZy88NSAYzJ60+83yyRcAkvhAxj5kUOVFxzrKPVA07wTb
Aacx6pRJWmOyzv9jAas/DXLBIB6MWW67VDV0S3oBavWVapzYc0kcI0jZdDh78iiyKg9mHaDsYbw3
ukU/oeeG6e0PfSD94prMB8YyUlcu/uIMNXvo8U0yjp9Ieaf/av1gMfv5ZpBXQXIBOGLOTMnzYw80
fF86Kp4/wy2xZZx402Dgro5BVDZZi1YkWUdQ65mvaOIUFS+dPXH4c3WyxmumZ+OIETblXcGAnsjW
1ugpXzzxYp9nhAKvvcJbWIgTO+b2iykHmjONISIHJoqz3RNzzMFVZtBVsZcakezH1oeUwcYj4/GD
HYwQhiYo2M9u5zBOpOpO9rA+yvFId6eQl+y5EyKUDBnBvOZ6dLcc8wMSXajmnZa1WM29tO0650FR
S5UkT7DKaUVflWYB52SatK5vxqsC29I1eL9Ir8mHLvXcw6eY+RKDHvT4OO4eqt6Wg2kGxpWD85ML
RNKv0I6rvqvy8ctyFnJF9WF3+5VOv/lEqY3CvOWzHpvbsC+fHoO3bySqLKngRxUIzBfCO/k5f9+J
ZiUd2j1DTLl8vySmZ8UYMjrBTqKBK271gaOy3fq8jpGmJoWOcYnIHLZrmPLz10Gn2sVsXar3PyEf
9vZTWPxlVzftDFDMJs1+QV2veI/Uf57+xBfm851DVn5PM+woO3niEhwVetUJIBQIXU59W8hiJLZ7
4a5AZQpvdAzUDBWWa9Tkf+a0Bv4Uv8QGJZ3Cdh7Zg1m3qN64xyh5CIm0xMesRwPSG/nyjdtAbSr/
6qZwVNkd0t9D/zDZ2KYv/XGVSIkLE87AZdWy7L8Fa/lFEDGZEwesxCoINCW+c+3CwMq3+6kgJHsd
SWmGA8C3wQuomAeKR2E/tuTOeJBqSxFSdod2w2fRNzDf0GVXL6Wk1lKaUmsgRv7US+16qG6pMmIZ
YkxM7QAdxKONsdNa1BuB4Igbe3/FDiwuqXP/YF0vNHtVBmCjpYQynLJee40sXSHSJ/kX/gQztmVI
nO/NckYP+fU2L2Z5u1bhC7hSve602dDMqrqu3htLNOVFwsNu2f2mVB/9lRmHjLuR5UUQ1DzmZXLZ
28qaGZpJj9THnxQ4mW+MOrWEcojzUm68IWjdqk29NsvU4zadHGgarHTYqVgewS8sp70AgAywvato
xlK4ecjorEJrozHHlfzJMw5kC0TsZmsCAiBcUknafSLqxIyquVZkID9fwYgIYlF6fPj2j3PRYveQ
hV+cRjsGbZd81oubMXfJykfVWxN+KBKWSyKjcGcYn3MU7mvmxxBYgvIaHWFGfNmVTqIAVD4GHtTL
8UT4Vt4MAlg6bI6jowJpQ9RSsQYrpRJ0GxhwPgFfWYziTvx8Hz43EKaIfOx+ThMn0rfdoL573gdx
Hn3x9Rq+TM+iTyOoIeYrxBWaM0jlQJdXX85KgeCK+iT69txK1Zq7LdA6DB+364BHUDfYCBTr1KkC
Oh4DcWGO98U01QtV/jXVLWJDcMIryPAzffQIQVwH7sZmTko/zdzhIWuniPrH9et3v5uF1kKzu49A
MtiJKMqo0/3nOtepHQJxkeabYIK8IEDGbnDflnAx6PlFjp8oyDVlmbDy8ZaMm7AgN20HH1aqYdd6
XzaCp+InVfa8dWdxnEdFOa5sr+fJ8NI//ff9dP2XzYH7bJp/pISv6gjNwFoavyJ18LvICkCAlbeH
2PJOv+sHHBEMc99wfoGb1jVdiL6MwYc8y6BRs0OrDhhGci9eiNh1r5r6UTrlJKctoyUQ3N2n8790
UD3F2kYlL/rhxNQkWSgDb8q8qV6AsFt3CQqy011a43xxnf+bpHF8NIhLeo5A5Et0OFABkgAtcH2r
zjzb4WlpYlDdEvcDAOkWOjvDEzN0+zFFUcB6MnokwigaU0PiweH4feTlKel/6hP3BqkFbguXhrpz
6PgEQxXuU+hr9CEyXxqwNL0vnhjYcvkEco5OQIuzvt1GKa+Wvh0G23mn8Qz3esQd8SkIqWcf3Fgu
+XnWcoCmuzavF7JCETYRxUbBQWtXCWvSvNjx2Z6P7TtVtsYzleuQEnkFRhNTMe1x0yO/mgH1Du66
rSImOyWqmtFykYeCZQMv+Za7idsHorpkR8M8jXRd25EyUTvlQLKIZ93DKrH+ugizPMB8eSbzhELf
P51PtOaKQrKoTfqGFImG85+flqHkivwlixlHgUk+YFVjWGjq4oCuljWlXBKILmCtzFh/XUbp9W4n
N0D4XyGX+olMno7DHn/vhi0Q5YvLgXo/PsHHrszHdiSaFRWL5ax85EJkyqdaaK3Td1Ek3/Kxw/w7
OUjKzGYKfSmqBGrYciqyALqI/IsWjdnxgqSoz8TU48hWQDAYwn/e+e4MVIdHOs68Ly/nHuryODaT
kRGKCAu2CLnbjU7n5PuAWL2Ky7+EdluipBmni7IGRV7EOlJJf+fHG/v9Ik06TQ6sJ7hSAWtMJCAm
M7FsQdADG6u8V7gIOpGNLngjL8YwMTND+sN0eKvATjfF3DZeJ9C1lKwRfoYZ0Y76RkfqtH3MgdNC
G1rnlG/zKIuOUfqKp5ox/P99V4Zl/EDW2dlgA3qZ7so5Gs7s/29NHfFwmFHRFsefPlifjvr2xZOk
wcLBgDn6zvldHI5TuwehgpYDP9yVKdipDY6BZP1m3h75M+OI+cwThiFEQdo8bqwQk39ulKYHBWGg
nM4MO+XsZgqFdMqiyiU9C2gRi3wOQpasoQtO3BRPG7BMCpV3j7ZAgrR64c+qHaxVMGf7AXiu6OY1
k9fS8+jNemy3erd3XrVUMXDrla7XfzLjTEw16rPp9SQV/CwCg+NdL9AryBLwk5aSxjgtxQXYlSHP
gjRvNzvI3eg1KBMEFI+XTKi/KHRXZAZsnHiURo5hyPHKGkkuCKSw5yZ0vqbYnnLcHnp9qO69aV1O
cdOr8sEOCUE0TsZqVozpoR798qEWKYXL3n9WYEghVmiXC84IxtFvV1SG4C7DXnj6Bnx9t71y74WJ
Ed/8B8rg+ClXnSXg+torka4Z2dBxws2hgUrDGtODOx+ojGiPyAbCc3aAy3hZhFgaCe7P898lIK9v
PLempph+lAeer5QgdxcPOvGpN8G99XGmaW6QPv0rcr4alpLKoGjBiEJFroUhltsCV+XVjBEcAJQQ
+bVOgKXZsUP+KcUaHPBP1TRoZvPs08lCOqvn/BSIXRWK273lhDYd9mtWd2hSfZO9K6ukXg7qoC8N
TXbwyjtt7hPOi3mTGWngEJCmCfLkB5wydLWNGjtJCI29Qe4Ow95M7FkSxaubG4ECkb8SAfkCK6Er
/ZnwraqTDqTjRaais1+cVD5y16SA2o8P56T7qpXKBL6m4ew9LZbHK5b4G/lfYU4Co2kEcs2UcFIN
lnutk8hi3M8L4h1frZVI7uvAUU3kT7O7HFD9fFM47Ygl/ggX5GkqlcNe/eTG/w2+Cv3ib87P1kTz
S0w90O7885qMIFT2lGnv7DVtXvz2KrM9qot6grITV54P2Yfr5N3oQyyYXldsAjcvmDf7+fwsWr8e
edE69Tp9vnsN076U3Nmsjk1XKHulO+o8pV64cBIQ/ym6lAgFCdWjfOPUR/j68Xy6PFdNzZ/KzFQH
M8YOV3mfCEm99KPena9sWM4r3fPwbdCpacnz6oZ+y3SQbPWBH6GE940sjJ2OEuhC33JZhAEmyRso
CRxBWZ6NxKXBP7oTkiuc9TUGMNEDzJi5aMa919ZNbl2DqqwYPltocVH81mp8OOPLOApaflYRSxHo
vAwcSdSVV34K/QZpKNbkcHJPC5dyyoxohgxGwBKN2DecK/oUsxfJz7iAb27bYkgClTO0R9u19iyT
ouMn7br7mrZOgxjZzU75gJNIEwU/I2BH867wvaPZ4GAATZgRX1PX8UcR7XOSMv0jyh3Eo5j10ZYm
J2GQNQ5Le5LFaLamh4O8hnQ08Pu5k8uTHyTSAncUc7Cezha919nhWpVWfywByf2nc6Dm0ElLc4yp
WCO1OnHMw9M0UNd3Y/PhV32B6G9NSPwvYk77GzOcIjBXSxqI/wzTcLAWf4rSUm/C12UeMP92SDUA
xVVjX2rlUEx0zwHM5jTD8HJdqUAfz+1E1ZoOaEOEqG8rkE2negLHzTz/CTRSr/OTZ0pA0rnXkCOg
Lm6lPa51ucJDi+w+xIUjz3Mep1VJAWjxYPB6rXYDkExmKVW96Sc7Zfa+eznuTGsLJZLVmJuNjeXF
FsPXPRdseta+1Zb9z5waspe5akj9QMXCneknsJbClhbhGJpOIYP7qbxeHhjPcIo6CJW56U5koDfp
dfAAnEp6diDG4mCGEZGqyWypb5b6wR3b7DHnDXUQlUhSPwkfkGogVc0oz86dMt7i0dOHTGPT+xkd
c0R3i9i8wCL9emR0rjeGT+ZiDPeEeI6V9RUXbltc8fSRo6Z+9g73u0YHucWOWidIatXgSPobTdfg
vcRyZNaGmqKhDyk2kKuP/O6I4WwQVsnGevAfKE87ZECvxi0ADCMh1RIGu1cn7QhGMWB0HUjJGDMZ
h6Z/6Vn8w6KopkU/ny/c+uUazBdTBp2MXN04y2Tn/JS6g7oMsOpFfuB7YdCr/fA+LYM65F95gou5
1CaLFYxDLWkej3Wo/jixpJ/Dp56HTmzovN3r1j03Hy11A9qyvj2dNhanYwZ/upInT+4u+IaVzKg0
AiaHwlnyjfwq1E0xqWMnvCWrFE/Yj0PU2X/AfB1o3i9P3mRp39XGYuKVNCqXVLcr8KnyOXAOMb8z
bOaW0RMqeSkCUfDMmbSfVDK+NCu6NLtXJA0kzpJdb+gf7Nh7Hq1//a30t3WGbf66Ur6Jbz0rAzE4
RzHN9jFNw1FHRzFcZoyHi+wx9ucQf8OnhCVRwQVoy8C7o2E93ErEZqgGCx1kk+WCP2W326z6KF1I
9v36hNroQi46ItobhaAXz9NMFssxyizNqcS52kzw0zRuZ4i8gLtzmTZeHcpKr2oi3rqOj+ppLsk/
uKabLp6z5hjcYqVrmkHnF+UFpVdUoDqQRWBBQricSeSAdHpfLenda5TTttm2Yv0H34vXf/W85QhV
uBlS8m51gtMksvk3Tq600Ggq6J09v9SHW6G7B0+0deZJMd4xj2Um+T2l7/DCiTeifhiSN8PBmaG6
P34dfKVWwbVc5RXyYKmuIM+MYox1Z3y9ywQeyEKa8wtx5YFOl4Od6AJVu7bZCCphiIf9Z2lK5ud7
sxUXu3+h8Gx5UbtZg6zAlAMHCmPRlFrSC4eqebx3j2R2tMeYAk/QuSEGiisxmvsY9hgoNv+lldcQ
TvYvBBXu+dVX3BMbzkyn6h4ccErBiDzP4mCAb65VMxeaI7Q8rRmAy1UWokOo8qUnZ5012pigPGXj
YVc7LHDt4h6kBTuChq/P+gSTb1z2IcH+Ux0kEyZWUKa1ERHoyeytKxarI0Yur+rx3EJIZ7nzhJpp
J2eopF3br8dCBK+vTOScl+xJdDGPxbaQG7K7M8F4uR13iLDKYZqKocOITM3PecuJdHS2O37+X8o3
TIYc9Wvl8VXWALmraptOncQLdScXozbNvKOOiY2zRMqlCp0zHrKnOSqcVCestMqWEFA1oTFBn1G9
v15I85HuC6Qf5uvMVQHpZd9uWqjPwpL7lvPsakjVJrMGxi+/mczdyJg9yM20qr30ockvR5qcIkfi
6tsoA2oDmry6gmtdXpJEoyVmv4f/O8WfT0xwjgLsNdZ/ixy4VGafaa/bRUnHAMjFF9x64K+LnBSe
QpL7KSvsfmFaq8C/V6iN4a2iUlwSsgpo4qd9tyMu46IrJB+CEuiYd9Hma+Evak0EumtYyqmqba3n
1RT5EsSS7SSTTPnKCK4T6/3hg+e0o7P0mvjyNFHs9+TiQPH61WVjA5gz8bbZUCIBdoA33GJ3HaJ2
hnQJrP/pBIoYS2/1toVEG8+c9wzqrGbc12alpPdVsBtO137LKkq/Q18O4W0A20nm1eEm6sF43K7f
RnAgqMlwTTusMJcgjvxZ0gLG8XQNRHN9quNsiLBY7/pdYXXMY1g/nQPg5/3ap6hbDPRYEkH8GovB
uOSgQUBHRLFkRd3OyOL91piilG4rXKgNSzaN5ygEkzhR4wlJvGzNZjQOfatU/apMsYvKLjFLjOD5
ZOK5uSkWsEpjX7nMLihpsPmrj4laQFsEnvn8dQHdyySdZKLmlgPVfqrGjkySd4rQMOIre3OkbwKz
e4SNG8/ZVveINVyvQiFKfTsOKKY1L3TKzFfV17lhey1C8/HiQ3SLaYngTclEiwWegSq5I9oIgfzP
UU1MEgwPwcoUfav/fpZhuTmw0g/zqzrr+SbgVqHYHZQIzqhY62KTf93IUqUdXFjLEz5y20W60Dj9
JH1sjg8/uzQX7QDMqXQxSmK4GI+ljresiTBOIEgmrb5936/qHAseXJmW8G31t4+qyF76hcRPgR9l
d63CgG54zO1indYDLsTTxo+0OZZtDioybf/iPWO66Bb7YjslLqqBUZ+wX4UR/y23jPByjXyiQ1G7
bhxSTUEYFWn3a5gjcsQ6s4vJljqTW6+U8GoOFh1kTGDhGVaq/3BWLFCRQs+LL/rddYfR/9DI8roP
tgqsanpTvIsVhDsnLnmOEZtZAhqQldrGRDT3t9JwZvWBO2HqnbSuY0oI/+LVJlPRGh6YobxDqe8r
Ah4W9BdbdP39DPHTrgaHqqeOnatlnDiWYO3HajRx5VdeZHyg2h4Ltkq3R8yNiiBw2HWbFMl/yBBQ
9CL5mVbeji+rVkj69Xh0vjTJz6r37pAWeAD4mJZvNoHWn99h0iEpdWwg9kgSSeeBlP+j+1Kk4ehu
LAfFUnrZAMoeRG1oc3OwCzfc1jUnW6b8QLT5yBIGNJvnX3chqXvqp3qU9XZ3Gi1secxo9xxWrlBC
55fWB7KJZltAmq3up4O308w2KamB5D9zrxwR3aSoIuPaGKidxJQzJUjV6wRpJnXvaxGEZNGL+sQY
RD1pgQrMmsQqdopEXPdS1G6lw/QOof/gJaoup6eI5xGV9qV5B0EA6xdoFZMaCIvRv2pvKBLnx/EI
M9MOO5DpLb0YkxQGWSDW/9K5EGxF/Aqp9dGJMVtnFiP7GCFCdXkpyJL/jxs0WnsxBtTAAUOi5yIA
/HWU6eXOY02PDWWkN63Z7cyE87qEik8CSRElywSyPCadv4pf/717dvrPVI00CDzf/IJIlL79DMFW
E1orCRZK7wHYz07+HOTgNW67iJP+YJt9+h7VACtUDSGSgLiieuBluPfq57+FbXMc82Oy09970Pgl
joKrHbTDQPQcgiRTbTJ7U/n9pfcoHE4sYS5xXQ4EhyVeVWPcCrHhbVyjdcj0bA4fqrQvkI3TBahZ
v+E93xIr42gBBsDue5XHGdxJxuIX9aSdLD1jCTKe9arz+ZPCLuI/bQkqIKUKcDDuLnNss9wthDd+
VVVQywAjkzHaFEM7PC8rVfi0VgnNk05wSNaGdG1xziGziSq512g3GC7rDhhUbQAgiVNol8+/RNLl
qgBuJQ8K8vj5pwJu7OgE8IFnCnO8itGjTBJthNX9i924PqPYp39DUXzEEo0jeVXVbHsSewO7Vckz
xB0XN6zdW/3SEsCQ+gh1i4wvhIv3JD2VGfVyN+LIbzBoRICddtDt2T5O3r6F/I1DAIrk/RpiTuuK
2GxFn4rMvhNMmhWK1p99NkZQqUr4Bg60A4nZA6QxOLG5F6hFIq7OLVjOf2cLIWe990/rqz4Gcumt
S4YUEvMEir9nYF3snKhpZmG2216nsPnepzWeIKE5YenyeK44EJ8W3benngeICTffURD1mg83VxQS
eaqMYgXjBTWE23PSFLzNPZpBSjS9QEZKzPcQxT+W4T2Q/xJMRO8K02b/8Hd4yiHvsR11dMLfFRlI
fz97gEh/gfGvjL8NEop0WlncAE6cuuDhHXbkleL28m8y3O0VGVgJUEKVDAAKP0TkbKqRJOjqjf0u
iBanyH+wg92ZyxWTUXSsT0FYp57DNqrub1wxY4IO/awIeT1KhSbbnM3wz+0+m4BeIxpMSufZVk3G
mEfwMbUeBeK24t1FsIWLkLZBvTiH0c1uSflW/1kNta10xNO/rysP1i0zJf5VoGtTxscCVDQLB1N7
rMVQpamJaLmAgd+sIQFUp2P0qzMGp129yxPdBV2XM7JG6gg73cI5IRiVcgRbGkjYZdQnmCLlMU6n
64lBj2NHyDpmFpJW/h0xV2b0RUC1MDppMCJdtGmjHKqomG7D5F8qnn8pMUye8zinZiLftWL8S7Cu
q3WCPyUywVieGhL9i9jx9pXR46gNubjOyem91ki4pOo/Ilmnb4ZqAiN4qXDUoY3XxTS9zfao1V3P
JOtmDDtNJYBJRyQ2NLpoZ8c4Jx6TrdcBrVfLZnzi0Og5JtVq876tC5g6arjHgx/4q8fOlfATG3jc
LFQMXk5MeomF2cpDGoX7KyR1GTvkXEcH8fzuWv88eDA5svpAO5kNcnvxTQaGLsLC4UGi3U9FKtWQ
F19m9uylgumCzIS/PfrMSD4Gg5xikgALcTFovvixwGjd19pKR2VTm5NCsPHA0w8BR//+8fMUQMQg
8EYzbjqDIplLJ+tF+xiMQyi+a6rlfeHY20up6EU/bqjrMJT+iDjCHThT2wA1oLp0TYJcfOJ+dD6X
V9dJ0T92Z0ztndenrHnVrgSIuzDMCDl25Ale5ceOEtQiE7lUxXBTSyUHiDjcHgPQ76EiULdwNb7p
HwzhiCOn2b/Msp+CAPxUak/+s8YU36NI0pfkZJVkcaOY8qOjwfVlnupIVi4c//W0KhQpSD5diAiM
4PWzwcz/5lIHUIPl79VJGQ3btktr8jdWd8jXFeHKmY6eMvaMZuDthYCEGz8OfRGMoy2zwhOMQM9a
4ZnF7fhKjEeSbVjcNoDSB5pbrRmqcutPmo/98h60hG9v5Ot4ccgMDuSW0z2gcLfPFaD2HJWrQf6z
YeoJ0yG4tBA0W6gBOxMU5yUK7w1upXM6xtlat1zFz/r8tTZAJ0+r4pk/Z1gd40yt3B+yWz3kvtmU
hBdO1GFidTXzs1FoYPqJYj5zz68BeoeR0+MNenF7uyNqKaSzcREmM61QnkFxabzouleYOIVTHzoC
a/hrLcYXgdbj25crJHxdtFPJ7I+Dlq7e0TFnGXQlK6uP0bC9rLwxGScguG/1lFXqY24hXdtZ3+BD
E1VamdNdM4pW4ZZ3y61CDkZ7iDM4pipQroikYNnq/QjxJV+G8U7m9i3ArXVfmQcUmIAnuvm4rgb4
+mUlGJJdGL2CMVnMBV8o0Hr0X3X6XVJg/zes8jpamAt1yh+ttRBee6muLO+YkmXTLfxa7F8ix4qf
HEiEYIvzP1IGkWVZirdBITQphiTSvPTAopahL0JT2j4Z3usQkMFl9IlSiTrArmyU4QnjGD05g4rl
l98klLtc7UvCEGNL5xyvV8YiGYi/9jiyVKL6AduDLphgm8BBUAP/NwpvLI64OY3M0GJzsmVSXhZ6
e3553LvtIRv71Q8V9oMxONXfWIa34tOfsZQP0Zgy2HdMBvU2xcYbCpLX0eF0eksTX+Jql5+83HMv
AEHIFsgFNP1Xf1fR8UMS9VhZL/htKZZQS9AwxXvXMiT+Y4xjCFOTGkZVITZFkoXydqKn4b5+DewT
EZWeXU+qw0QetnwKV63lKA4CUg/3+f0QHosRRPkPUw7ZsIWtiHloIRPJsw51yr70p6Psmh5hYq6o
JOgnxakxXTStAQ+Jhs+RVmDb8MXYq1rbC0Y/I0oZEKferKwk44RFRvUc98IxBgAJN9t8NFwGplFd
F2bSwhneWcSgOfESU1vYSBjFuxwn6wGavVjVGq313ocNohrpBKlhvlgA3IS/IsBwdhmfHZBBHMGf
jGmTV/WMEvr5bcarWAigu/VURgfTYjyMlo4GEWn+3Rl1wh7+sV8Z6DzobRZDq70lhTwkdMy8ZQc8
w0xc/RETr6sxrUm1GPapyHq+hTNAJuoHpnQj/NRo9MeK6de1/SzcdKS9Gr+DPTZd52WksGz0H/Th
CTI6BGBXIZ7l0bcpntKitoEHmNuq/PXxrSgnm0nsJrwXJjQPaVXhcBuaWKVzh9z+BpSAMxsXLLsX
4xjxPQLll3k5i/kRfBQ/01yMwWsBoIXxal7zGThKX4RPFDDCIJzXtAdtAlmZGSavY37KGwTb+9lo
K502hJf3OC0cuYB+HEJqjZWswTMIVhqoPHSAGKxHe709NAoFI9R7jKRVrQ1x6rwjFTH1I0+jSXRa
o6o1qcHoGtnnO55+wvvfBeSiIoiXK3HjnVjLinvdqY59ICud8/K6EAoaLGUHb7LacEzI04pYFmP0
ZSwRB5CXeqnIV+TfA141U/AI8yr9TusLKgLeVlpNnbUyjsxWWsiL6fxnqyOLiVoIYIvLzXMwwgmL
P3b8BS1Zd3sUHqTjhQ87OvDkhZ6GOrGxgFPeC4eiQ5eUwnrLsOeAm7R909l5orm+B4ryIPY4zUUm
vyLnQtIBk8n2V6qUB15sMjqYe9UyxhwxPexhIoTiJs/D7m5wAgEu0wwhP65ieHv+fF1+SJmRT2yS
SIoYRV4B5sxGLl4hPOAI2K7HVbJ1o+1qrPcuSa62D+AFY451xEzqpZufQL2E41lMShONz5fgyPwF
VB2EU2BTaFWAVBOBpQo0PkO0W0rinRa2+NOQJdFIkQv/c/9HlnEjAaJSQtL95JSWrJ+0IIDwvgd3
DDLcJgjSjWXkqYvK7qDeqJAleMqa3E09ZpfJr+hOPnVmeHm9bjSNCppUQWFuYD8+IUeCiKTL5CGP
pg5HzlkmaxUrh5Ma6y01Ne598cnyM1HTSVSd9I+zx825RE4tzAI5vusKvDoOO4ELTHqZ0QrzwcKp
IlCd4IlrdqbYM++DYOZrbn+LkyULGZc78vQiWvX4+ppI+fyVDZ1nDx5DkxSLVQ1YYUmwD77Psoo4
ekAMCn8l7qOfgM3LvPZlJ1qq7iaQgtLwXttXljuWWTYqmMbqF6yYxn9YfBffCu4XmWfgA/QPiF7p
KwdfsgCK10ng104jSdb5NqBOk9ClIsr4CRc9bK+3GxaBylFo5aP0gK/iFz7m23U6PUjfeuy11kRj
XYlyE58KltnkYm9SXsn6JEhJbCqKJnEiS3yadmJuiKnkheEB/4/8FmsHzdKtjI5COf+tekNvWtkz
4+EGJMyGLeksjZX6j/wXRdMKjBr5Q8jWf0AOHb9Au04gOPBWAo1C3ke2xwUQMVJDJaK6eAw3WpZd
wL0tIjNvtZr5IPWS0M9HpZwZ5cyN5/6cYGkDeznEG0BZJk8QfckKaoNNQ5ZzjSZTZ+yVE4MYpGxi
0j+NtOvMKXOqwFAvL10EzoLQfx59GTSmX7F1dZCI1a/XzckAVlUmdbg4lZK7ERJ5Gqtjtcb36L10
V8ZBasT75+3jl9j5p9I+n50ifSM7kbqglS/WmHNOyXq98yBnKNvsOPgfgLzc4yniCITRKalytPwM
slTdVckWZa4UJF2o2gLkujVpK8tRbdPmmLIUQMFLse8bMmlne6uToYYlXwZ51NOIIGB47Ei6x8Te
s7e/98VsdWJ9YVI/M8sgIoiw6bBgl9IEFrnvV0Sy9EUXZaZFFk4mmAYuOw85nJ3mdo9NwSenMs3V
2xECDa9c/sj3r0/WkMUV6VrTBRYBYVxiR2MvZ64WK17QYgsp5AY4/4PXdExNMaEfK8KMDQ4BSUw9
HKpDIfo+GpVDvezENeGUT9lyxBPzUzggHfTv/5xjDJSZ64Z0R+ZT3G4QdLyjZr1ryMQVo/VAr/JM
aFsD652ikc/Sn74o2HTbYUjpRd+5Vjz8k5shHwfzt5lKLDqz4kp96v5xx9t7RzYqzyu/QrIIPbDh
wsDC/FR1C+Ojz9MyGz/NR+KXROKBZ6vSYItJ7zZBALEzHQxTWdUhPug0BitKI5t/cd/MehQcH4Ba
I7RghDLydJ3x+HjoyMg8qzkvRJ5sYQZK/MvUH1Ys1QWk9llD0Njw8rPlXg7XB2At0nzOwEo8WCjX
W1ilhstCcH1XSGwXifyTL2T/UMWm2mxkXdq64ujig3FngczuquRqhzDWsr71+8rrsefeiOpLfCuc
GsXlTECUKQVMdv2dbhO5ZJkEXpZTYmQORj7xZlneLaQnd8kD9FEFLj1cokzJ+Obm6Cm2aM1I5KeQ
8M/wWIAj0y++EiXL+zZLfw+ViPRT7pCT/VQH79DYJU1AJSQqFoNuFpiZRoMXFQ9VHOH7jRttPT6J
UNj0329DJsphOrkGcetsLbv0uu4ERUZV5IEp85KG9XPpxSImQHdqopDq+qOgyAIE6s3Gy9HEC3Br
/0Zk0CG5uRCIWFDQC2RXA0ViSR1ECiL13MUpiUcEC/j+sG0RA73jrd2D7zX8ZeG5VALYp5klt0rU
j1iL4wWMtCbSWUFq88x5MTF/9OT7YFs9wzQxyHtrMSZyiVNqtxUUTToDTBKeRgMnE8Fcld5PE0os
t2ffU7wmSKpC6jpieyMjkbme6On88xe1IkhG2weXYdDyStJtlIrj0wV4ayxqzMAvfF2oG3kmfAyr
1UrGlJOjUGtvcfyFoeG8zBjXn9474f85cTh/ryiuxWISP0TJSWaMaJsvRK/8qK438zO9GJ/OfK7x
RwFA/2GjuNwvfSKGwJVDhi2U3c6aSohD3p2rvvAVa5BAiqiJgY+Ln1hsrnlJpDni4lXz5tdEgUY3
I/63rAzhogXQQnnQz7ocEfYz0tobTJtjrsgnss5DyMr1wTjqsUZTwjl99DewyJBxYganBrRV263Q
AcDViGdU4wwL2h1Nki0kK5JH3u82/UbkKcT1nVuIkY5KPleoJBtC22Xi4imrovJh47iRCF7wTWqG
UNwIR36BYuBGblyfUCnvm9fzLk5TWZhG5i/ZI6Aowiw7QzloRchhBltnSWg7P+xjiR+5uteStK/s
l518KIcfFq7CVX3ZSPJyEVjvWh6wvCG6aRBYSmHXdmEcVWrwY8xqRFShpq9bGI7EjtVOopG1Pfz9
z982/GWIBOgBxd4cuWZZPiy7gjJ7WMLcr9uKmPzI6SXQ6hUaFecZODw7+ksiLnfob5ManuzVYEsE
m68ak/UkEodT74hGfYw1eb4xTARDiG+0B5wZOywimmH1rrxpIu7O/gwRsxUAS3+EyPh+sMCOdCk6
UB5+Rso0ltHtTciCKtrQbvJIA03fB0mO803awVdj7JQA5U6E5wvNev+oDmjvX21yKhehoSy+kVOr
RxPHQUGT3Q0I4J5+uTtA92piDEo0+OSANbzSM/qUGwMldjK2NQRCoqVyWq0VV8vEWdsC8fIBKb78
eLY3XZKeXPuaLY6w+kLx9fDZn4rtQldj40F1eC9CseJrO0SczQMfYeCcHGOl5u5WDq0V91xAzTS2
8Yw2q8JpGZcM23UAx7LbbU+MtpHZdamQb7oBKTtd5ymnTo7TVU0C8YNBjYGLvNfB958CAX0i1PsW
68ixwCTsG5rHdordSIln9tYg6N499P54U6KO7NpcLnAgb5tBJ2TDtHEyZygXPsgFf8KDO3elXRC1
xYCTr3jJui0TsPvq/6lRBYFXA/ShxVIgZA9gyhhLYf+yeYqmmwEzBPfxvTf+7dg7CvpeYcK5eKu8
zAsqgFpCnqZR3jt+8cXLdlIVdwuHMvehdVIzD+7KnU6usRvU+wAJPvwjgudiq9F7h9icVyuGcDIy
XcoUxYftFqMDJ63WPNmMmls5PMY0/eovFajoJQmChp+kPtTvUDwNW1PljaGqAmBvDCl+ywe3HLHK
AZltZ61YtLUBe00PN+wRtrkjaLGyCeWATbSOCbRAEIcM+y8ndcOfEM4Q+/b3Wxkhzr0MA1YlZcHz
XvFY/8cE64brOXLp2tcDdUetyXxgP6nwL1b+T3tnuXCg4HiVMJK6r2UdqzbK7rlfyQ2qRQmB4Uj6
OqZkzL3vxoyNZTkWe0TJoXXRKhTHOIeh2I1Hg8mTnMNf/YqKYjKgpLxMPK6JR3+ddqPDLN77vGed
8aL5FFBVPXPuE2r1Lcb2afjU34r8aa/OPQ6ZxfE/k5lWpHFiZ2TrdGkYaPBPeZcgFnjNtBphQLLq
tacGcThkOgHAtQcczQYZLviEH+ZmY1GhXfbkdOJuMEgXSshGavQbs8MUn3sw01smm/Yx6rq50781
wuEjOdDqo81GGxT0du/2Fqq/NUgauH1+9babXX/2okw3lo8FhPvhlj7xU10njTIO5Y8ccPnk+jZP
2TmjDSOWo+4N8D+tAaSFsIobQhGQYMxdXLL1wx7N1sTMP258+7mKtebhkwZgPK2220v1n+DrYi6K
An3dwAqGJNZk/inlTwfh5MYLCKwlEQOJENUas/bASQGsi/sCfHT5hIkW4lsXbSTO5ayXZeFeOpie
G6jodQQqC9SxF4cRnqxjRYvCDrnzqGA6lnD4Vwd0nRqAhJ+C9NvSsvf5K0zC0g5kiVQ8HNwfMev3
IAAlSmeaUkL1Hpm/0Ob/1U3nvxqC0t7ZsvbVXFwnHLIwy9KDB+mKMPWjBUq+9AfaTejHVysvxQqM
wh3dlMbPu15q1kfKa/BT/Ez1MgTsvLHYSAZ3MC9ORSMqDOKWof33bIYJni1nneDSl2QiHgj6Y/tz
yEkslCKEv0TbBmRIA6n/WVdRzNVrNuv3/Fm0ibbAwVv+qYLjhmohaTeqXic38nGCN2FlFXpnAEh/
3kEERQxqWTcRaZsD75tTmYwXFvgXIlwnUW9hoAm7lsPsbubDe46mnuT1QXmje9kpwANRuMye1Ghu
hAydJJpOh2YPvQpt5oOr/tjPspy1nYozLkI0a1LwsubRzsJxcKOKLpsLn4+gMorc6Dn8VqMmdtWB
+gZSawPdDHv9hWPQhdRwdg9RQJIgDoirg0Cs1kg5+jEMLJsuOXXem0RwFTZjKt/Qreyq7aXJDGJ9
ogGOCQBIAnJuA+TmaLkGYpfSxKNPZy/PIGQYaMrEFiyMe/thsGha7UwbbguHkEEL9f+3+6fLSuE1
fu+qjq/6ILvEA9YIZFWeSy9PdVEnNIJSdRfgkZXLtzoIjNMjP4ezr+JqUwj8cMmB42LG1iM80Spr
KmW3Vf+IfhLNFAro4agvtixaZXLKTJuplqrep4wUvM6Vh8rMH8Fm8v50gMK5Ii8XDU4MMlWmrISZ
lsUHsGJVZyYhwzZxMXMdW2+7ElunQEd3NfvE91Cx/D8j7tnb/Qqo9mBHrUhNPGKkClDBDYeMyrLp
0TCpfYkWvZOJjK6kvG7qQZ1cN8YYDK8Dux/S4S84ISZaEMhtT/6vlqOOxWLEl89ywCUV3TqCPVWq
P1Uq6b0ZpHmSDpvg0zgJcHFNb3v7K0cvS6Yj6ABnHewNIhaMBemStcgb1VUIPptXQ3oeiiTlhZ+n
/EyjUPFXZYriPPQhPdpPG4hq0qCo/NoTwi48ItsfM5ZrBTOc54X9/7/06jvCdjhs/IrVtejit+zR
/FCahDEjMM80Kq4tJZ+ryc2jtJ34Kf5rkgKbVP1zyOG2nNePYdpmBfDXpIsjJdobFBEJXlKWoMdj
oofMkOk4wq2dqUgCHYwj8r7JYqi2R6f/yBdfD8h9Ht2x+IFwpb+FwN7zcSpFkRdRPiqD+Wm8Z5kc
62gY1Tsk4w7ECt140JvRDQ6zqqHEsDsa6ZvCPxcqKIsr2kJT7W2T7/31/GX1g9io34rPZAngYP05
PIW+CCSYCrFz/7yubs3qZ3x8+8g7OLhJxbAtx//cwSvv73DrDRH0EVhEnpetnrdRicBh6FL600sC
FbactGRwHaCpORCtMi0ZCGuQwUZrQuuRQ+/mhQhIssIGyf4x3uOTxIiPhjR+bh7KBKwxb9dEeOT+
XqvawyocqEr8AV90rQXOuWcBZpOj0pM/TctHGrLIut085EFb+iOBmT6hQKqpAk7Zb16VT1xUXiL9
9LpmrDCmEg+JrQbqWdOhP3M5RuWE+ZdcFklhUMGxUki7UjQFaFOY9AIJGZfPqwcXHE51r30OANAr
vnfldbOoBZO8mkdvmc3roq/XMuJluxHs+V/nIJnS8jyYCteC1PNNPpVrJraicHu7/iUr49Cz3KKg
xazk0FxVQOrl9SOCn/XKk459rD9Axq1KNUGvkytnUJ1NUbrh0H6CItrVUfHE5vCKFpnBeMuFamhH
B80AtuJCSAQlDv2X3k1ZlmSuqme0tzVGT4P226udGZs7hW/BhPq5s2Fe6QGouc2q7T9Qv7GCPala
cm3uOYnpkVpKx46NeeSVCIqtrMu32id/JmgyQAw2Cj1JkZyzdp4zGxfeYiATTfh+HtxAEvGWWPPq
OTBZn6nRL9DNK+etzK1qzc2wU23rZGEZGP+LuxcisVymYeQL4jwZHiT95xHso6ZPwPWZvkC8hL9x
Tj8iK6xiWhQoADQjut72v6SXK3aX9m6/Cq3WseuXSPa8CL1xqIkFQpbC4V56EDYt6+9gMJOYXLnl
Uhc4j1SmTGnh5VeRZqMzsoWVZwQjtkNsAaaw/86HNkESIZ1ayzZlJTTVI3v9aqgCyNanOgPfHW9c
d3OJ1VH9+U7jrrFPMspEDCCPy0aFLyO0T+j15bc8kvkEJrZzjX+8OOmxqktQxLzOwOTTwoe/0qbC
zYjAjwrW2V2oKBcaQQzRAnmQxFNR9zeCQSMHXRFlQUioHBmswk9SrDsKeeCzX6Hyx60x2PNGcH+i
DTXfgHSjVeNJ02Tipx76Yztinko0me8YXoAifdqYbzzXefiZF8nIFYZBIyFIbONgl55cDY/tiMok
6UiAoYismEJ4CRPPA6o5KRB/4yWFBWMP3z4fC6IFGPBVKUwknwgrYEnjTkd5GUMC2FkKx3W56Xhj
622vVnmdoZ+P8JN8yoECeEJ1GlL8LH/RbzGZ/pg1MdgnnUYGBDvNOlZob+MLuTUZD0grJGGRP+DX
2sQVoc7SBXYVhyK5Cett8WmM/WfneYu9AGYb+C3NdiGf0KgPRCqqlYX5T5XqTrKvYUNkiTuJgfg0
0r6fhCM3EoFTszPqYF4TX6iWnt/MbTiX32Tc8z6/q0/CvScFKYafjOJ7riNhFtu5tWP0Bdu95b2b
lIa2gCZawByN2q++PQjJWLopygYVTDQN1RqyvqPPOfVmYbrKhlvCWg3yawmpiho6t5G/Rmsp5KAc
VlXDrhfcLfsZMEYUDRohWXLstwvC130lMz/Yp8bAcngrVUN9DTqaeTAmAktQcx3kWQIVCkgPKYWP
iYiV7yGkwzRxUrCcK4sWLdixgYlWrFnjFrRrABmPlHxcl/kNfWhVZo/cseWYW67vA/mueT+3lgai
Hw+7x8U3dz3HqNosDnNhzb6VQC9H1sqEfLaCIUiahJAU3BNUB9XowG/Eu+wtA8Hr7hFTq6tdCOsN
eMAaFHtV/PZBqR7OYj0x/J5ltcBDmYtEbMf21BlwhTha7oROUX7b1kIza2WPtbF0aeXVft+Qa7EU
RaUMJBuKZ1+8Uo/M5uZDezDrgZwe4rvu4N2dlTXK82yxnqECAtbymm8Ctfg8n0BAc40FxgWROsWA
PdDC6WhurldnoGfLlDaexUZgEMhc0cCX6r/G2cP7eZsfj5mwfEQ5LdQ30Vlf0fRJ2V3C92xxP1rV
r4JAq9rE9rVZ6xxVKZhRWVrGOiTtPfDu7EvDx7GjzN3mZBzAl0C9lSHTmrfdOfYqpFxLGqN07Mv8
/w8ce79+JLIoezQtYQfVDFYGmR2QDExoYCp+fsfO8D4CkdUIk3cXVS5uFBnN4OyKWDBX4JZvg2D4
fYUHecEqA3Tfu3KfgNN7f4gVQR0yagkpkVYAUWepY6AD7reV8RYXtHwi+Vm1vsq9PF3vYFCWA+om
5o2Ovo7x5OLJ9CIhypRWUdPLScuNyLQkhkuYn0YNjOltFN2pRNOAevO85ygw9B72u2isdJA54IBA
urS7wrcSQMWZni3GMQIo2VEmuyLafnaHU6rHKpOmFK7HNZTBs/DbvWdSU2OVXGd9RGMOUIbwpuHF
y4J3VU/qYfcFcXnR0jm57sfuxnrXWJnESn1lbwhsXMvHf/fERjaiFnnJdPMCTtCY6uUHilJNNjdt
UrVUIoj94faMqTvJHwRhoz3W2s1SYjuhF0EXkig3BtvGoK/4Pa+x/iAdEw/Gw1Jc0sRPot7i5rfY
G/nnznrr0TvyuW6UwbNuNaFSA5DUm6pDV5hEKmR+znf58QKh2tMoMmmxt1mEqWAcTgWGbhNAl9B5
1BdNb0V3TX26dmY/OqNbjRhyKxjdxzUwJ8zn5o6tCUh80C4G6hvFdK6dkXwoYScbHXQYIcAwVGtH
nZGujXqCHEdFuD5lxVUxqtu6xq8MvNm92b36/rvYSyZrpln+yrqSMbj4qkoRpl3HdEHDCRpEJGP7
NbCG4DcHDpz35YpG2QGjKyCut/7V9NyOPavYyH9jBwuebTalkV2XzLVmUw0nK2e9WmEI6bu1BHO2
tx49zKeYikZP+GvfrYnluntvs0A4R2Uleix8AmzEZSJD/GVhP4gBVT4oZwC/Rwy9NUesBZcY23r2
df+gdwCWdvXW3wnlv6bcN08oWU+mvvl6QUHi0/ZTfOY0nWW5oH8leYi3MxpmSD02ynqr318roCMO
1+KtNCciUcT9LsX66Dla44vdRL/qiZUAu5Z/L7yTqDcadHew2qpWcC1wJVRVT4LwOkXITOFec1+v
Ak9pQXw0F91hlC3j12ccSBzU5xqDYuiguGHD3SdY0irF2lq5wMTs8VgMP1TbenMSrzWOkVeGUXNQ
GVuXkxt83vT4/QDIsXSEiWNwgYYZriH++yTnY1bP4OXTXMbDj08W2+g+Q0vzMacf6aRybgGok+II
60ldnLokUSyUlJBUJc/PavSdb25AE8tsudK6EC9ZH+1yQTyhJOVTo0/a75ZBu+FFriyyz72h4Ttb
JeM+j5Bt8h2ZiX6o9JLtCkCzuioumGwzoCucd80FvXsv8c9GgoXGFY/DVzeGLuXUGgTw61OkE9FQ
l5/PEwyXHht3BfEvgZ7mXjly2JtCzstB74MMaioVKKG7IHhbMHTN9lhUfjXld6wq1N6dFdrN5LQ2
mtAqUyJXfRP9e7MwqMFjGERUHZr+Su6nZMYfggG1OR+Rz3G3WWgvaPTFjkx8pDo4n4R6FiPH4gWc
Ese4wfvaw3/IKjIGqtq10+LEpkxyN/ryuycwckV0XLkRRnbdiRI1aPB2QBDQjr1GIzX4T23D5NQ/
BS7vE+ju+3R0ljSKA7cAXliaDQswI36KdonyYUgzQlsuovtCN7lzVakKbRAhoM2gzx11FdnKIWPX
e4rvj9urPTONZnFliWq47SKlPyE3K8yNEfPo4+IEqXqxGq/oSd18BU3dkhg4xym5GgE306DEo9Ru
l3nO1MluP3+iuMcDgQrRR1J97yJlBbRLFDk8LaBmSHcz5TaSNWK6Xy9B/vM76PrFB0TcMMm+BhKq
5FV1djRTPrt2Zx1fNtyO20VgaGOLyRDOQeDJ/kji1W90634UAVFWSBtr5TsoroO52aeG+85s3UrI
8qoUiXCV+JtR36AoHDfLcaHafaEl2zfs9jF3b7503gjAJ4e7SiNmySPZ9MyClM3Ov6zFDiQGEHU+
11VgLkaYkWLGMfpVxVPgkV/wiJeXl48ZVOvb1Ya/7NDz59NqjsEfC2yZbZkHz9bSSuYzJO0nOTYp
humbyplX1siQ+FJHVZh5drUaIhyHw4Q6RSBLzBU4AKEFLWD2fG3Kqz72c2ljXE8uShZiG/AjPzEc
MjFciOEd/kQ2MuGED4rXHYBo8FQJ8FWcdlvg4ULGyrgLaUSb4/YdknrxR/PtGmMD5jv8UYHPbgmh
Smqxr32O4vtkWgF5tP+KHght9Qbp4XdGGVCJc83nYHPErpFjmScvSUAAz66KZh+KgVl5FtvRwL86
X2bdwtAZKZlIWChijAyZZWzX/yNQ0XApWK/Wk5uc5O/afb4ORFgFUKGfC2C5BrQP941xZnXlXQFd
bgsCn0tp7StPhvj0LEb8+ylsb3Ub4JUUpT6/kI2h5pJU/aNPE2MeekMW3QYN6Ur3rxu6Dfih52ES
VpMkbaHFNsupwUEEVktLl3LG6MvPXJmGN3Ves+VkInEECqmbP2FYcn6rEDl9HAj4HbfUlql78ECZ
v18T04ooXHylEEN/etXRq00RGQrseyQSqURuReTZxrEnFWnrPeuurtgiUMfPLEoTTHoMpl96XVxL
7qqzSZtef2Hr9YN8nqfjYNTJzX9h4j5Wic2SGJeQh4vSpaeF3b6A7ZBSDLjgv6XL7GbJnK3omPGx
0yfMu2ApA80gO8Ce/aYntSr/y6Ebz3h5wANlJuYbT2n4QKOm7o5hL9MWnVwKQpnryDo7fRpOBJEH
vqkTOFbNZcCF/DarBY6ErmeHS4eO88GjGLa61WzJVFd4PyXC8/oYmrHMKE9ZWL0yGkFjo2ltu95u
EzSiv/6a0vtEFf202+VWhH9+4MaMMhgLFj5S8JfVZXkvW1wRF4mkznaBhod1Wn/mRAio2ybygwTR
2GNKHRQ5kFLVMi/vbpB/3TxiF2I+/AplNOkrM+nG7zH6cj8IDzS+6zuA4Z03PRSsqjszkSk/LPmB
Wdj9Ipeqs7hCFHd57rsXGtps7lSnoKD0IOezXGReRyw5eM98OTOkPy/U4Q8t2rwvPivyWNwcPEIZ
htK32xU6lE5R/lyLAY9TzznQCiiBcZEZhpVNoC+jASTWB/NqmwSVbGtnySvtSeyYIgcB7N+86TcM
IXG0plfNMyH0aiCtWNPX0AFvJ5UEXSOGoGqJjzGheaCj3MZEWcVKUjsZz7pgEWjD8tyjsTgY5YyE
7zUP0NsZ142lTIuutWPg7nllqz4z0vEFbiBHQ5U3NYrFGa2AynDoSVrP3TgE4ZYVotODZKpBCCqY
cHLXzgMdD6feUVPr6XIfLCCTf4DZ3QNXHXzHn5FiMsswFUH1nt2+89Wm9oBRvE2F/QkIoScMEB5E
1Yh4bD/EoCgYcuj3YjzBD8Ju4ypToMXD6Zx1PqjEajw10o7WMcsmmuddq1BfL8eE/8MIbE9Pgvf4
3/jhgZnYF73njASJ/+StjTdhiexJILd8yBRyEKCj+aj+IsdS8Ok8+LCBkU2yjAhav6fifjuRigJb
08DjBkpb2l+pLg01lXGnC3JA5rA5gQxrcZgE+mAmnsBZl0xCHA8Nh2/Xh8xAmZefi25Kbu9hMMPW
2Fab1R99VyiWWWHtw8Lg+ajpne7CHYbzTizZUT74u8QeNnrvewxDOLzGeMq/9nwrHetPzgZe9R1h
oDXOuVHZtYbf+Cc++AVHVX+SLzOf2TgFf9zhYSEXb3UCHXRjiWOk5K5e0Jm0NmWEV4hT45BXSRao
yYiI8VVfD75GfpQemdvV9pp+u+pbwtSgWG20UMice/XStdwGuI05fUiCBS5HgELfImZ4bAtfcI6j
OrP+7kwz1fUaBV95MQCi0S8RfvIFApGFmXCrMEAefTkQF+9pCxFOo4xqVKkHf70aspt70OqOg4xS
AkpQPpZ2MPkCgUWyw4YMLo4DakkGAVmsUvIAWgb2YnamSJx0cRxnwN72GDNrfDeZ/Z3yiQMKksn7
JJbgPMNr0SgzmYUyS8E/GFiZv0wrqcVAYFicNlfZQt37hyyARcERFLX7LG+RP8ZFG/vNm/Jf62+y
YQ0eQD5rzi1FupQzKTDseCmXjY179ajALwuRuFUC9r/hgGRzX4KlQfVebA+iaRfrlxRbpkkZT6ZP
PjR4BTapbwyjF36olTh4SKO0Wt0g7N4F4Fbalseu+TEwK2C8C1mj9GN2fEtQmIUpwVmZrrUxVPxQ
WpMwHZ11IWU10AH3upQJE961rAYIYupm4u3LPLLnqdIuUgfYKuvtanLgDmr94Nw6Sr3w4dUC7/4K
fZ4YkYj4GtbIZewNeH3pj6AyFVLo3EOAP0sK6eMhSKyPcpmkmiY+nihOe6WBzDjzgdXcAs20RKzX
oVC86ANEW/PDJ5ti2VC+G7Ja4ef6+09m0yWsBkuZELrZ0JL4FIJnGJ1UD/NA8NXB2gUOjQdhpF4C
h+nTUO7TvvUfsmhe7k56ikOKI61SlWtz448kpCPbwAht8ZUC9pWpcLIIVWQQAKCLxP/xdHjOvCo1
Ob8q9E9PaHocYK5X0fFdiFF14gbtg5dZZyjboApoFy6rd34A4A/Ye5PFAJhQlcaMm3CMd0XxIKXm
gt76tOnelCSMBs0gSdO/4zlugi+nYpQEU0RveDYSa6l12l1U373aI6s7xShfSYDiMaPNlloSoP+f
b0s2JRM5DkBy/lr/78Bc439vVstsbTOuHtKS6lAJb72zZJSR9qbvbDw2CLMgDuAhJ3TdmO6EwH2Y
t2j4CQyuXtzzE10NVRBXwygC8BcocOS57xcKeNlQzcEnsRNSg1/T8zWBp47JC2WGZjTd4dH3MvRs
pid+asdss63XBDEjmYY2sTZu5RjxK1xGHtR75QOIRJlp1tw+c75KS1zkFxwppbOFNzVbIuW8DOwV
0RQXcennfIe4+CfFWKduSrXMQrlBWTVFcVcNzcTaIa8F5SmVvIS4xysT6/U5A1kKYyNVDjZZw+yV
XOAeEPNseaFDX2VmVvgHCPuESfs5GUvfblTZfGrCIqVFHxdeq60gBWpL+NgxBhC80oBt2empbAnj
9wkEZmpl5drF7GJsBeQOUZGQWKgtYfyPnjBlvDXHc6CCnRFFqNFBw/JQhApWpK9qN0udU6lc+W9P
CKTfBhQY8LOaNcfV6HJmwlLVhKoA4zEtFkL5ouE/bxeMG2LpAlvoea1U5IouDqX1gicdyH0s4ITk
2KxWSg7jCYh+KID1hUCwI5Eb1aW8FHyHMcOq4p2JZbltroHd7cdxO7qRgdLDbynRHwXBkNpVm8HY
nu7qOM7hAv7VWsNdTEOpVemXLRHh42432As5sUYWOArJFM6WBzuMuxC9ElVJrV19PEjJ1LymOtd0
ChAJ4D4exJ8JuvImguuHBtebkW6o2t/SyxBTXpYm1zE6l8VToVKAARueQr8q8627z+tKOrIiEO1W
Whi4kx1tq+LQyAQHKdNBU7sloDUMNfmVkxLeQ70vcMXcwRA5SiFPXsusyO4YF/9uRBYWhbBQQBHt
GXZi/8GWGQcSDqCuc52bIBgGvp/w8vzaFYAK6837mfc/+b5N9II2mE/ToJjC3fTVCgQpKC664i+F
sdPhOxflCijExORfRwTr6g832jj0k0aihSILAo3Jz3HJ38bGBrJMZBgwrCnys7G+j5mEiRN6fDzr
v7E9YhG2v8Uzj1Yr+/twMSh9h04WvayNKx2OGffC8OQLcp+snZND4dUFz4GS9IGZ+/1jAA8CZD5i
X6lSGrrHwrLtCm3fwr9eExxM0tVSGheUBCtA2CaQ1nzrFMapFfAxy1l/a5Tjv9OA3ljaPxvxQ6AR
8w0vldpHwo30ZZhdQ1rllQ51RkiWQAuiiImGT8sHx3A4tTYyHIYEnqa4Uv2HNpWNQCZHEMQz55nI
gbg5lO8+Sez8248qfRVF9FHCyGdUcLJ6txHmqO6W7qkOCWIzch+DbVDpxkf3XaHNAHDXO9xGg8Wp
XHED2L7t+5AoOB0pcukTTGQhARAOEZXI04ZN4RbW71fiQCgNFRh4x0zFQg2/ABZSpyNo0iI9qcWJ
9DPKzrHvNioGz/Ik4PgyP6kLjvbwBI10g+ZK1FdnDnlhK/LW6S9IF5eC1x2vUzLNqkBLloj0Ojqk
TVgEDqnEO41/PFENIGe3qu7NDsPBHSnxcl5UU7sj/rC9cKmdfSr3pUeujQswWIIuzGh9VAyFiVm/
BT1eaWc0HsA+Uf603ij6AUZdstJsQY2MgEjhRYbktwRzkAsGolEyABsRUgUKKz1CWdI8kJBP8a4i
/eLmXBxtdgoHe3yMGBtti09BCG+Hl8nEPP75GOtOp4U1LAEpsfol6mqeKJTauKY7nmGii9ho2loO
bECwr0D/rS7ht3TssSPoYrAz7em5EAHyoCrEpzLuzYS0nmvc2Z0GK/Ea1HxTftt0zXdiTiqABqUN
OwAPAyViPTUeSLLOQ2bm+v2YyOSWfCNRUFTaFZgDu8x9/jleQx2biazSejxymzgluj1Z8T4b1u8U
j4j8F3aJPrC8H6Y/56fA7anyw4ecMarszGsIiCxIrfHVKtAWanIVvMnH0gq1NkBgJGDHUhnJ5mCG
tYG7lftz9CEbgj4/Q5fErYDL7XwkTb6q8DHZCQ63o/7l22Aci3I8bfdsig+0f/XboJcU6VfBgIIu
Ys8hNmPwoeJTECd4m/sYyv+Y9sSPDGwXqPIHYOHm7YnnTSXc3bkHFi4jmLyBjiYm7E2Msr+hjTiH
OcrGxp2kwm9CWB2NoTEbUe7WYlxh3nhX+W4KU8HnTWNyPU/KFtUmocZ5X3fZL7ZD/PBJJexSvoIi
ZvNatm4SqsgJfY96ptNrXe8bvMDKGZCnDTAOQU6gXeAEONoJ+kHO7ETf9pzQv+qp7ygIEZs9AJ86
BECl69Y2V4R36iYRiXgzpT968l6BSDBOUomZl/Oio8tjkkSsPXHGcz4oKi6mCfteTK2bKG+eS2Ad
4m2sAImnyc6jdIIn2FF+pDd1cR/hYBdzWrpt/xQDnJqvxKIxmuiRbAqwtJ2DzIT92rW2Vv1KkLPU
bw3YsjaaNTfXZPA/C2kN983GqpfmNhuo4XdX5/L4rzkKwGow12vpSRHcKDz0apL+y8l5k2viEBN3
GWEtpQa6xKcQkk0lMSy2aC8NyPTotJa84GAk1Moh7Z5KvtpI2NMOqWBqrYi5Tr+tjclmx12NEmig
+CWbZOfbsPC0rH5qFMHJL/kT1GB8W1AMkCSZhUYWRrVgRDix6d5KEX0obGDslnpaCpzRdjBYH6li
oOWz6bFN2G+SYFrKNTKszQ8ZH1nNZfud2Xpo3moWQKsFZ7aG9pYWnSS6F1914ar6xaqpC99s8unf
L7jvVNqAS0raPFt+nmJZE4al1zn5ge7mwfJqjq2p8rEXrrpkB05HHFRgQOtXsbzmq1DCkRGu5uBB
hbTvEIGFYB/fGpFYzBt3JBXAybipLwryl2y7Nm33CVOGqbUKo/xhLO4LDK+YwzdiTaY3/H8Ci0GO
nUBch+Dw5/KsN5Ij4gEel0xWndXzrtChgbGPaZ7IjC4J/cyXDiKneJAirTfGN5lwh8zIhCFpjc8Y
PSE42klv9tn007TH0H43vlRNor86n+e4lU05ds88ILImhvJCXhhEPg+Ronp/Jx06O5+fvFI93L50
jdX/N8xDNMXqxrrol7VxAnYdKtHFueZLHarmoiZXAfFNDOLB/L3QNSsibklmCjHnAQPcFLV+UE5w
NaZieDgNtkw7Uichu7TOYb7oRWItn/DR7aF0eEe3uSDwc7EIT58q54HXoR9JiMSqWlgcwzUfCBhj
R1XS+LoX+Ef9vTdSixVK9btAXgq25PBomryFf37QE8VN9e5+3m4c7MOhgRI7GI7FS5r4u5GJHV3I
2ugcZ7vyfeelpH/XB8y2tUtTBhZTDk3n7ce87tIQQ9xrz7K0UkNvjKMpOqxMyEQ3F/nl8ypmKF2K
EnbiL/Uwa8E1fHySO1DtZivnZZeRT9ZF3v0je40ivw2K8EsvIT4kMsnhuVSu3/efN5n05EFXC5SY
El9y647rXbPNdmRpnxOGtynjL+cia/PXfiT3ovh1pxQPx4D3/YJ74PVX5IffQoaRRjBiElhw3xE4
0mAFz0m0dJaDIah8bNa4R5Uh7HMjxZboZgj6uIJ/yB6f89v12+LWYDkoUbky/GILb8iHWK4/W/Pr
Fy7N4K0S4rnllJxE+5fRoOwkcks/2xq4Is735JZGPCsANt19YNRiZeSIWCrVBYNvWle5w06ujDoX
mP/VjqlIe3NwW97VlEFuZh/F8HR7M+r0UsJtOU0y2z973/bRw0W3gnhv+oE/h3AYu4+0TvOxe/x/
GL/4Ec9zMCTB53XoWH3gUpWxqlFdEuzoMaBDHiBJY0CHIWzaENf0nfDHJ0D5sBuC4teLz88E4tpB
XfhmFwaHcAaXqL36Q8wCHW3NC9xwxKmgGBhVGxppEloWOIyjyoE8/WwDzr/f+/0OaQc4iFkASqTs
3wisjWnQ+UUbAd3KBzl/IB+syuB8SInI9+Glmf1OA4erXr3KyurB63iOv6vV4cPdfIOywpinLnRs
VC+SN+Df9B5Vmby/SYQ7/H+fyx6E907m6zSPTEQ5Hc0f0ZJr0OMw9Ko7trbLt7/Rom54FRD1Qa2/
TcrjcZqlWQMco25Roi0jWN1VlMTV2M+noy1tummzfnLyG5+G5Z3mbe/zDOhonG38sRHuptiJVAg3
75ORC3SX+jghtjbveej6eAafxKTU7EboVJsd1akVp8mjl89i5LpZLRZchlXBqJkGQ+4LNKlDLRCX
XnpUM6AMKTNmh+Ulm0KpsuOI69LDuam2MDB9uJwR3fxtRlMSRZJWocamlKKiTcfC3xzO9gYgcqM7
h1wfnbousvYFSyAXZuicWh6qrLNE7Fpn4o8zlAknkZq/+J1jv0LfaRxztmfUxTt8vnRwsrs06zfr
GZ2bTfi7Aub+m49WzjFDueCoMLV/gjhLVYoQP6fU0c2hpBuj4lr/AYAgcmaSjZLje9bGSMJD07Di
b7gCE+1rS5SF5SAtVsvJ0CsCWwUkaMjIUnIo5UkRil3ocj+u0vc8LIFXjd6qishIE4XUA7NnBRL8
bCY4etmHrr5xWHtmPCiATmXhuXsxJA1zonXdnPuq7iCCKKxyGus+aFY4RiBGZ8VuQDs6F2jgw86/
sHlVkounCFj5UrzeDx07iw3zqhsK5ZIDOhIsQ4LmYDPmo2vYA/tpVE7DHB1uU+hY4j4cjlGnr+JH
SfA8lfAvWxtrHlX5+mNWPkw+z9Z360xIFnQ6rzAhaPCydSc39jhqVrUv+BtYngNHzfRfHN+qtFUR
4wu+he2Mo2G1RfePJ+FXwkup5Ci53BII88qG5WG8ZVOgFQRUtbNFH63hkxRCHK8NGjU+k0X/Y0hQ
GT1N5OA/ewC46c6PyJEkMYlfQUp7O1va+TIGaT0794QCEPPNzXXwP7bVmM2+baerZOSjDh0WTkwK
nIYU/iZWvNQaEqSiz2PSw1yyrx8UvDAC2eNvTsvVsrICIZL3/CEDyti51q/cLHgzUnFFcokgMh37
6FP/gDa9C90IUb5fQXR2aePkDeXknZeejeyFF2zgJcMeQK1EELlzlk28jFbs3hm5/quUX+ya4vvk
pkdkDA24pZRGmNhfkw9PDTDznUOZDbpDDLqi6Q6nFaNSZ0eS0De5ht+GLgVG62C95yB+A6Q7pkMw
gnd3mU3O1T+jSnqAWidqKe0sFoLWnbay/afpF/rOZAb5BJepQQAVcVJyjSmRikF9cQ87fXtYs8en
FVE1l9/IdyukiNwjAEjGovF2W0EIqgkFLaaPfF3lV7UZimf500Mw7PC+6mlO7zT/UVPBhQVcsqTQ
eGHDWJf2kY1KydiRLJa7MsIzSH6yjFf3w0vZCTN3xSb7txc4Lmn0EsstLZ+XwBIFbGI1ct3QncMp
mezkt6r6/r6kKcZ7ekNGcAYVohiZq6wKWQPt6nbOvF8D6wA6le4wKqlmdcFkxYX6jtMGdcvGfjgn
5eyjAzLC35GgiBQ+WbVW25NgXS4uVWTX3kJkNZNaZxnMSpyijba+hFXzfkV63pncscmZbKhzJnch
YezfHpcj/0TNROHsKK02I+cMLxnKg72o2HTFa7Plk4gWpF326sHfkAv3UJOkbDkZv5fkKYGTwkKc
5qmbFAfR+XEGQZW+1pKGf4IKyBfDRMlVSdGdyN0ooCm7TRgJ8covls/7EZCjPaw8BEpHXeRVZpIM
xUCSgQkU5kFQfKqBO+uTtQ6GjHnQgRWzqW7onQP8pY1LWF6Mi7nztDA7Q/sPZ0R85WbGZ4YIzftQ
MCUi2Hl5xyvdg0npLUAhh1KEAY9rDila8hjJ/ElSY4fmYSjWb8RRnp5nsdFFP1KO7cZwd67egBQh
EL63UCQuxYsiiv45f0hwFCcpvViKOO90FBOd11Nqby9dF5Xr5+fdOJfnbvYQNztmTPCxVWUHzsrE
UCsofLshVmC7c/LfFWu5g8jG01V6DeGKbGOj9ERO6hRMN9RrElfRGG8Z2W5fYldee+hfsBXz54hi
4TL8jVEGjYzS1HEUwoB+nv5U1OVe6P3TSFrYIEONy97jE36bkHxMbe+GyC5RQC0f2qDxJinOOoU1
wbJrlq6xq9lOGIDBuy5+ArBtRoiaIjwOz7uv7+TQlrEu/McseoANcwtQVhBGKzeof4kOKy670xsl
+CkyViUghJNrG9aBA2lcW+AKEysnv+3lnwLHE4rY+udfIEgT5coiuihLLKt/UuIArejY6cXQPU0Z
JSSmfupGJuLU1zIZy+Tp03OTSz1AHr2TgNchEa+pCjWLyI81HlovSZra729TKI5LXAerbUWM3wob
s0cDG4N2LsGA0oY8r7Dy4+B17xU4jJNoCczwYt9StFzGl5xVVKQjUNmeUwLyqUhQxuGuQ9BOjy4E
jkXrakkW92VgF1xB/XRde/RS8nD2a8h4hOe7y3dxrW2xhg8CQWULNlkKT0cnZRTX+izuSIK6KCVZ
jhszFPyXFeqYvNIs2+/+oFZ5cRy7oZnxLbsIKme9jvgtjEB07Na3YgWi5GoUoZbZpVFg1Fvi3o2Q
jtuIwElwvrAdBIM7wv/Kul5/sCES7rK2jV+jkPk1ccxoVwg8o2hMk8Dqlm6KUIKkZaQ9kfd1EvRM
gjI33F1grsSSOWPb8B/c9rVlWQXa8U788EZmaUuoiTbhBXEOOKSXgwgWsLBeSXxWX/Mt5V9CVEug
WaPZ79BJJpxLmgeEmi98zgeRmzgw/65mCteJloM4NmIbN/iHTRfPnBvGoI4ii8++8VkR/uQoyj6r
djPZ4xiOoYNREGGKn5A0mCtqF/WnZUj1+QUZrLOPTIRu+rJKbuocETsrKra4mq3/+bAddfBtwf8G
gFA5ecYghT7tedlN/jjC3VHcQhbHAOUcluVgPncvTcUxKk+5A7yxnMSc65koMf5aZNgLUI6P9n8O
qXRKKVyGMFcSY4S0u7j3uBaeCy6rL6jjmAgM5K+CUK1VwwPjefWbJ/eZCo+1sopOIBJXG5uZgN4G
7fztxQmfTw6VE4c++UUs7k2uNT0b6XtLLs3YJtWkQj+EMzkefklx0AMBMpE6ZaOHxgrjowZ/vY5F
yWi2AyXwfn/k5Jk7Is+lUfpXmLKLiVdeqIq9Zgepu0AfjMbuMHqTGAzdcmcj8gzmbEURBtNYuLb8
43em4/iasavS8wN+1krpcOo+sDf6nlJ7njeKh81pUmDjN4+lohhWHyGQ7QDZkHGb6HOBw/mQVKKO
AyAitnHycYCtorqNv0yXTSwnweE9bzAJyxuSCxkz0e7DSLHXNpVFb34WZ8Yq3qHEFYQQttI948m4
C44MjKdPdSu3KNtAUxfBf6k3vIg7MLJf5MMo3WnY8FXNtHNveLqk5M0oE8M9v3r0NciGtm1dS8wS
fXQWvJfX1UuCW4RSDD6+I/h59YekHZccdzV3Qlx7xfrkYdWd2qCHRKO+kR9WhaqEyo9c8I7LImGK
3IEMFsgCIRhDCbR0wmdAdjsCypuywcwldPwaGtZqNFLntjNQA50ecUqIINzcVaiT8IcDYOrqmT0M
7yejvljlqu9a0FWENnQO/3QS3k8z3zPKVZPdR+MXwuE1JBFiUSUZy1p0UBhdtrHglbdME4Pw+TE+
G7ZqYjEVnfXb/n7aIOWc8+PCgA9qyTXFR/HY/KHxAosRaB5448Qp4nCvtBkxu0jyT4o4y7PkRF6G
Y+nRyrLPdJqxk+5iVwTvxkCj6i20vpNPDSAfwuOAOWAdn4QacfnoNYra3R5psQJIH9+QC4BZf6Qz
XGD+vJQcya+vmXD+1tMFWPUbinwGBuzSqP85stCUcvvvzzxijB7kPY7K1tmLrko4BsVtLhM9Y1Zu
bXXEj6o6NJnBUPi2X6XRmQ/K8CWyEHS0PHJ1NTkWtV2mRlDc6Q5ghif3IEGEuBDZ2m0T2QjoDiAQ
3Tqh6RoN4VdbLPD0zQjV2OIvU5jX0T+utEnSGiBtW+kr75wWCSBfTFqduZRc20hjHJoQYNViXE2C
XEEYb2eWRYBG5VFVNCZ/jMgHG/SfVbwgs3wfvAvg+FEHVDsqXSC2Qc0qLxxVrV2w9HSeBiCtl9ls
6T3kk16zTETF1v1tlqH9lJUm9Wrsz4QbmKp905djA8Y9Aut5flsCDBsv9zcHmH8bu5BMJC3727+6
VpbsnadbAa/5EqI062THmXf1iIZhVU2BX/ii1VO9GLaCTquSv6CxFRqXaNl4hAG7Dsc989NWt4Ry
eWC3janStb0TXBZXam/qnbkrwt9gshe/pfrtvIpuvOElUXn5nIIXq/LKPnVH78DL4rkMJr03irLx
dWAwVuOMkaC/cX6veEzlBVmm1e4cNBDSORmUVGpdMIQTQ6KXZ3PFS0wNNbFJsxYc3Ar+7PPqwdXD
oe9TVElCg4SqCpM1RoCOPM6kZ4i/tdbS42QWOR16dlwHdhEnMUtZq87PiCFWH0a4l7Cp3seIIffo
cB/pkHKWYa0Dgm5XWaW5S85itqjsVjk5JiCOi6OHA46xN9Hg3tGzhE36+SFoDHmAr2sDnIMWmgbn
bUHPY3qkVkN1TdMA8ImvdxiE6QyYosQM3Z6H8Iw5M2ptWy6bebtwendRj+d5eYWSeWtWZOWvbzsJ
f2PVPxo0O3ZkbLYBCIkPcInOWu16lPDhLdq+jbEXzPRy9K9vYKHUalKzDFyFljMCvvr8eR1Xz0o6
qgrPB38BpnSeMFzHXfyQGO8kFjYiyRrJayMHWWy4vPkIQORCAXzUsOmOH3F97e67wcis3bQ2ht6Q
dmjsvCNSjiGR8StZde43dZIabVg4b4Rmtvh+XOjZ1iuKRnLJdkyRpGYvokuw1tNvSl0M7PcOpHbm
IY+b9pJPtqjyy51bAMgh4jfWOSLT4M28l+QI2i0j3V8txkXqOOT6tXUXmLg0OYT9xp3MsiYBtpnN
f8FjZ8lLL1/eEvhwSxuUcDmAkni1S+SwJcoyyr62lRnlnY+OKDFOBqMHMcXYjF5jL690QZJ9fSUY
42cvcq8129rxg4kxGNlxKWUipHKbcwgJLsYsaU/HmgM+I7rFtBB+qhZiwsklS6IXWnohKReMtifv
kteo2AfYZy2dk30MJZoD7tMG8/7pftifp0k87wZ5Om4z0JJ2iHB+3x+bgUWeQACjcpjlBIQZbsSm
UtQlK7y5bq5E3u9ZPjnDq49UDxuVeuWpLrrA/lYs6+J+H0ECvFGBC6YZDs+G6z5EH70AWMZussrJ
hPDgh+wQn+rWuTmH67YTMdJN8THGTjWBsfwBB8Y0vGsTzOX28QArQka5A2Da9xxTn+7asEGV5KOX
M/VxVY10qI2jzlZJS0SJa+rMCT4fcGlkafXdqMCwZV/w8pHEgKvgWcT39ekT4G4Ezp1GwvG4J+bX
SVggNR+yzSBLz5S8gokKh3Tto2GwAZBLgX1X3Oshi++kXOXah/F7oO0NCPABo6wO3DFtq1ys0M/V
D2DZo+ECpdZRQ4DMvRWJ9tPbB+fxbeAFLAQfE2XHyw2DVPWR8eRDkqmuZgMym7TQ8ELyNlYLIH2r
7qnHCFGgTezoa2RNSYvYS0UYmQRIBUWH5MS/BbFZY8ovCvTTDVBhMM9IRvMihZ4sg7eMbdlTLQE3
4MmKZPU+mR0uU/rp92LFAVwdNQKGx5LZCdaE9djVJXhul38G0ZccFY3x4E/yJW8SG70yyApUy17n
Sb1jLZ+r+v2jP/pEF6X5ShR+vDNjBVv/UBwAhm0HgxsUhUHT7TSeUxKZBYmuMg+nFXGQOAa1a5O1
u/lOCElKKvPxckSOJkzzJ0NrRUPLpEwcZ8rYgk6Amx9mQcYRlME/YooSivn5NoDMqMdIpe4nHHNy
M0/+KOjE7M2BwOO3zijsB8/iYcc0662JbDqf5a7pbGh9gCd1kuEWU4YdUTrLYQjCbRMxSzn3XTVl
cvGmTEVdBgKfMMlqkDYSigeHOtcWXWjUm1ft0jmkhch6FSM1uGh5eI1GDhqo69ByGMgba1JkYoFP
QOTQyQioyY0FOPD4o1XkmnGtdSGVR5UaB+t6wqtefdPNJq8c/hk8R2lmsEdL4i0qcYnZnWDhb+9D
1tNqz5w2BWq9SOlnSKUtzpT3oNh5X8iU1V7BYaqWrxU7eKRz7GZK/emDayNf2CntTfXLzFGIE8Wr
o2/ROBqERLu+3I4dfHFCohtOssCUrsvJ8eiEC8mXUM1iKt/MhahFwDZKzxVM8YYxt3BtKY4MiFs4
2szNXJmLJuBe8k98Shb1oqQQci+1rjFF1OpCSbnSHDTArtOiS1g0NerU4m+PHOEG7tUZWIPfRgGS
FO+gFk8IlgYYoXnux4JddhfhWpCDn3lTF/iIgnkhoGtSRYsivhzQLzBHMGTFKvagiM00qTSNr/XQ
AivCQ1Ggae4MESchH+3HKR3vcS+Bj4NX2nNrAFFI2JQaKDOB3SVojXI0AmDVKHwrW/9mpNbYYX96
TJYnILVQl+RDSOQHGD5I+1TV5kkeP7OqD1FJlzmMPCDxavtW1CIt5PrxCx2coa/WSgfF60b4s166
tA3YzUCjxpY1g9fSM/vAYeJueVHmgZinbfq9f/rbP4Fjf6B0BxAmOnzGFZxA0J+LynyagItRQHO7
TRDjNLdE+Qn5eWZ8T+CA2L3lc3QF0tVXAhrlVdiLICCqb1kj3CxCfodfPeThfJfzvGX/Abd1uQKm
AQ0kTqSS0cagKGyyxOSG8hiOSVLHu6nX5WZUUR2Ml+b4fuf2A/Q1RHprDGt/YDv0sd4y0mZYxqaf
Tv22rkIy31YJuq0fsVTDi2lCo93kMTVGEtOO5T79kRIo0S2kbugqw0wfKcJXPjowGjH9BARKe0zC
PUczdSKPbHRG5sJuhNtZ71nGo6VG+RzPcb4NuoNxxUMAW/mI5q0DvT6jnDoxP0fk1vJfwDStXzwK
GmJuFfrAnVaaX3P+zZkVdHOPzQ1RpIM52NtBuTjtuUEQEuw/WovcsPScP4AW2SKmj0rfNR6ICajK
QZhQb/Uvrlk245yTm5x3tOEzHBeH3VFQJll3+KZAV1Eg6GCGLZcH5A76DbtBmp4owh4o6keYuqfM
yzktagai8gstBVyHJ9pcpMcjUx3R/5kyhEvdLTyspp1fycohOChtP+0PzwcS9ONHRg3X55ZHjGqd
0Uprl98PZs3yJcX5pDDTpoSeLxKoTshjAzuD7eEtAXrPWFGVI+ARQgYzX1WyYpCNUCCs8aCEQfkA
h1yJfRKbcA65N/XZeN8SirkXRiPneU8Pb4ebqli62T8Ij+jRAGVMlHpIo34qKB51ozs1OkPdqr1l
N5TU8saPJn4PEffubsv7pbu3o5WDEWrghJVjpFjIePY0mcVLvOw46PoUTXQkcbGWxXGgmkY2+GXf
W3/tJAZUoG56jJOoBQ81t4GxJ7N8ZasN8NTi1qlQGo0J7TF4v7Pei0RlxYjzxkjGtSWknHMl+Imu
a5USuqQsHmMKH5GLEMqylJr3aPfBYri1D9/XePN9QvuILSdXM4VF72HwoxDzpNNfkAGHsTaauxTA
DpELtIkKS9wEbh61+uG1OxwoZwr2ux7u4dBcRzHeUDwQq+qk5eig+cMkTMFQll6452FwCU156tFE
SJ/l2WD0Z2nT0WSNvE+be9emwO1UxeliByLtubY091JvCCrPsuRoiq95fFJ0wvTBNVR1QOp1idw2
MWBx3UHjsEq5ryxdbE05/f8uU1xB/SjIbjyxFejhbXi13kayXuAGKUTYg4NKYRk6GaDx709P2kvt
oN8oOYbOgzBgzQniInL9/Yzy+nCariL3sUDD3uX09tQAgfPx8f8SRMOD3D4jdWoPJwqqxj5IVtWP
sXBtXWrT+ByZ+0nGiu+B3h4nsFkJH6ZYr8HJ14sjdXNZAsZBtreuBi1QFh3lm6MeXLdXLru1V22Q
qz+nJY6bL0fzemYopxO/cp6BBTTJNmoOZYnkBHEbByiri8lMfpLE8V2fBHmu4sxtc28qivk/jEoz
9b35q1CG5IfR3NEoUj3RM4LZh02XtBGgSApFXQAZbxbzD83pqGB88gCqfHXFZg32GzeYCBSOpqCm
ZuMw6FYJvoRUCevmflTbBJi8Qz7GezZWBI1zqzrv4qrGdtGjcGp7ygZnz9sjfAU40Xn9nc6eBl3I
m85WUJ4w6I+ktZPFOi+fxDPZNFDjRbR4RTc0M669vSH/VCBIH7NOba4EhemfLdFNzteMf1/6h0u6
JROyNh+JTbQ0cZTqw50nJRWnCnh+Fno7eeHU8ANkS0CgmwRhU1+Kr8tCzLJVJh0sz9QYWrIIjTfL
A3kuWsNKaInu4bGae62okJOHYQ2ogYOllHNH9uO68oQJwC/LHw3qMNw10pDTFL1hbDFEVIY7i3z2
ljYEA778puuuaLs89c1j/KW7KuJZk79cfR3kbT185XlBR2DbOhmknqewr1o7/AvGDf8esOe3zvEg
NJ887w/E50d6hAwXKXIzvJEQG0o7s/PQnjHJAU0JQFiFZRMcs/8ktbPWZNiag+wssH7/2n0fxZVi
xbMryccKWsJxkLkPpTU0i7j9jAs1A5TmBNCwZV3/AcNzQlgobaQv1LWSJqvI3W5sqDrWDTq25mjT
gIDDYscRhfVnXnjCUFH2BxyGNG2pGDkGzKnXXZR9aIvPW9gutiOJJGfUSJoW6nS/Zu8lhFToPsbF
aQLAK6mD+xBf8RX07T7SXeFHlpRn3KJqp96h5LbJ/R7NKGDP9K4yUchbu27E8Bv9/PMfJRpZyD+b
W9YLzaJqG4ofTRl1PpbFI9XZ6AY+gLxHHJ0ZOrbJak5kwIxLpgKW3Of8XklBo5zx7JaDt1vY1RZ9
MeukWHvaF3eobuA/RHZ+c3EHT4WcRizaFxB4mZkBD58x/5sb7jC75X36qP2i0p6TTrY4jUv6OzIC
lGGRI8YQlNjKSv3/20hDNFWmisuf5HPbdJHAfZdb1bE/NwVTR3bnH8SMfke8cOYLaNWUZCCOcP8/
Xu28ZWLdYCFeYRI+haN5V43bMv35pcek+7qeKlRDAyBxGZMkHPVXeKGWYy4kCb2BFBhSSK+Hd7ru
BZHO0OZ/9zi1Fe+K76ZqZtYwH534527BDMbPWA34f2dLkGd1gXqZBF3I+kbby3b69rYA+b+KhBzr
QDldBs4wDDKwlEuQSz+apfjR0xb4pUPqNIpfos7vkMNaIMr0hGH0Eqd2bA6f0g9yBJrcf6hHjQLl
Nhypv9GPFT50EpKPqjEg3ORj2ewraPHZ/Cp3wNDG2zP98VxbSTZZLSVjmNXwZPClfP2BvdEmJYPs
R47w+lxj4/8DQaO6+FN9gCvDIypMHWhHV03/NY7wsW0SPi6AdI50xBxyjyynC1RGTKWj6Vi32vNL
qPoA3fBAUcjdsjbhtcXxntoUlbx8KPZFvYOdx/XPTx49QxtxFlIEtJ34IU96Kj1qdskkRO/fw1wY
Sz0KWL5KQao7ENMkzq8Zf3UuJTQkrZ0QZfhtQZQdn6MX23/XCQ9zep/Cl+qCkWkkH7s7fIi9hNuI
SLS+aMVELTbtpR8wf+KKtT5AkRqy5oA+hASyZT0iD/GtkmR2w2P1pDe8jhK8Hgczoz9IFCEpM0eN
JV0lJvmX/gaQzHMgSfChqEeGJHUfBmWLu08PwCaXPRlq/CTEOqHofOhOM+KPwtYQ63dOt2QESeLt
2OPEEr/NxpX7ZPzm0yKX6C1h7EkvnnsbXKkb/oDojYD2ETZgogcag5vslswbINGWXTGkwMHl6UPo
YSJVPH0s5Ia2B/aR6wx+STn6+nXr7o2EDWu4z+6o8MHCToRABUW0rz7DXIXfXIf34+/qiHJtvtBT
laOiznKjHuRY0gZ9Jhe3tdJob/Yk4pimS1z3V4OVjF74FCQXlJbqKrfeF6c5TMtEshwKSkZmzPK9
a6BTxsuJDuYEag44iREODlEGWYoHnrWD43bQHPgtBb9u7EXAxw3EkOZ/1a3RTRDqpX5NaoEpFe0K
7ZHohp8Y5e9Ouwy1b8weupJQ6w5fi+mfKmkWpS9AbtLp2WFnKqKIo/q7jisaOUaL/BH9QUOzmt/w
Q3o2mQUbIjLZJh7bzuFpoNd86X5bmFWVusGgus1OGBa0P7LsuIiwrR11VjmEyMeqGOvQOyuyELTF
lNr1CE8cwZzkw1PEOPDw8jgSTADphtItACFcmyHU4mv4WGkCmopAhseionfI0oBWo8ra+0AoNg3i
vFyoPYlEPoHtwMOkfknUmYbh1YDBK04sVT6KKp78OvoWObgOVSiG4faa9Nbl47JRpKasY9T9NK1Z
BEmwfp9bPqiwCtUaznvcyn+6aEMjJqfTkGOtGNdIY+p1nf53qjiLWttZvc0iAtQnMIl+Xl6Oezi3
+Q+hMpuC/hpF3VTxtY6XxjZ+LpyY6fvMpvHZcyWcrb9rvIZoO2wcQd5cW0zeMEhh6t6TfNRdDLSP
IFL8XDGj0eSbqR7UVvr5nQ6ZvPFz4Ko3qEe0+kGiO+63e2l9oXonRQeIpr+DDUlPRHK/+xhaMbv4
0JmuNQgpGH4mg234h34yYjaF1OszvCRcSQwkPbYgcCXFjMQnDQYMLyguE/qGfUnn6AblNy+a60L3
y47CP3DJDhYeND2NlvJm51J9YXp7u9XqfcGGgzaFRm5aA746wiXD+qeRR5f3mbInb2IWKooyEJdm
VRg5HDdwCSGyIDwgsieYZeEPadwQEdFyW+HH5aU9bXFq/iUCM0t7prdyiMz241cyMMTxbeAVcv8g
yPA8XeuoyDNCwdWS5w==
`protect end_protected

