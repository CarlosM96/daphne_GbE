

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nmiQPan2MutAqQaWVXpAjvZ/iBqwFNaV2udCHkg38/HGng5w1CAReMeMp4eoyWT0w5TdM+B1sAZN
lkpRh3SLrg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
rTaXdaK4pNEb4nP+UlpQ89SjuOwrWuLxXAAzWU0JBSoEksB6FcxBbpxwhcTRHQmHlmxaeMCDJWhk
n1Ib3/mmIbJiHFfZ4AlZ2LAlBG8jXBjNLN3u2YQ9Gyumfi8rQPrX0NP4pwUkWRNTBIvvq4ivTW6B
uU9S4t5h0brP2EcmVKE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HljKkcZBLE6swTXGAZwJ4XDaNVq2NbhqpgzOf7gSWWgWlgfIpmxyVdKGQKEy3HdfLWwmyu92hFZH
S7sFAV8njo9dCS4qW2Yjw/aai/QYXu9LzvtmDyPGC/qzP939HJy34eTm1vASDGbG/LQAYXFl6Ud+
4SB5nhgeoTrIau0BBfOsZJkRhz+i/xlvDFlZqY3M+Z06Aj12g2CikutrOjxPYZtlkckKKnkcYiW7
sSrag4mEU3ScaCHgk5PT5ZcEVJcfrqBUH6BDkdnH2zLNRqJ79euazX5WIqc7Vx91CgOMlTwC4pnX
sijRmJcEyihv9q2KA248X+mVz0V9hqQu+LyUQw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PHbUyqdfjPpjGv8HZmojeNoaIdqeq7WB1IoTcWcSNbELNyf8DL8XT6V021cnImlaHgXJu+oiF2Uv
bbGHBd6lWElyBL08p4SVcTZBiqgpy1RYI9ohRQCDDvavDnbA8aUKDVA7d4Wr0k26hdXy+hL7FILs
bE3F5DtouY+eK+2Ih0X0tPPvreiEJqaMse2FPvqZ/Vk9k0xNXjg5NBqm4gFjWUIMCMw8BPHzc/5z
pAYlvPGLvWRn4ezrQUJ6tpRKLHN+P5fJnh54R10IsUsK8QxXKJiqBzAA4kjsoThlI7HKVkm5pq0a
oAgRQ5HYWjmzG4FMdENRHkrBjL4T3l+B5RQnpQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sRytgESmpzr3kc2dL59zopgGUtPThp6BQ9KxdXmu4H9ammZZDt6kCeXy2Z8cgHn8J42xvBCwL0dI
b05HIHKPS814/tufbbAayzTSQK6AUUarqUFixef3+NjPE5+VdvH+oSprTn2YBrOokm4W29e8RRAf
0gklFlJl5pBTzC0daHM=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qCTR5PpA30Wsah/AuFHZx4D81ed6f9K8E3/Ax36i5NlerXDpSvWA/UslKHZIv161Bbxs1X1Z7YVW
bknbgNWkS8jJmctj643ETMaA7gbG9WaJIxGA+eQX8HKccA97e2eEXMTzGAFIseBiRliZStbI4yNa
5q5XnljoZwLP+2ws6fXtR2mSiQA7RArqplmOj6YBA65jDj730BnwV0RibzW1LpUv+Gt8xzIu50Cq
bLYU6Q0MTdQ8hPNjx0LaI4qpvgF6ll/s4p6nAUiRdrnVnN8GYDJ4aEs5og+wMUQ8DhKQ6iogWevS
nrRVV4Y2Bp7bfo54QIyDDrilSfYrRf7idQA8EA==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pz7iPBzWkPbekwJORP0wHcqakRjx+irIN6SZg2Dw5XxH/PBrhTsH+q7RrHNap7KoQWI4ZZvQRNKN
09L7TNTLDlcY3A6vZOwOM1IK8vIwrduWAV95IZT/P1SEr3CORuLLh2WJaeSwTJSt/FKl5tysaJt8
Ux6F8Tt1wweYj/S5rAD7oGckZeaEZb7mdekY+U3hihiE9nkkBybJwsj1wuaimaFMzp6QgvxAzZE5
leuFMtk7gnkHEm1UnpJEVzzUukaVZnrDQ7908Ddx6PodBMo+DffS9v2/OjqI8wTgR28AaDthU28G
tYN1ifSbywfJQdh+/453QxENkb9OAGv1Ps4lcw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_11", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QQbGSB/b6FeWAHnjf6uUJKwcgoNrUdHPdhgefM5pdVMItumzE3AkHnKjALEavW4wN8yQx13F610t
tC0uuwgKoe9mMgByi7vUHu2gyGUj6aQH89pomXvVwbZHylI/Pz5WlRI/zv+mGbF+3yE2Z/gqlGIx
x0rRAHMvM5q/tEb2TYFjEMn5G3D94Qa4gl3HBKfOL/k7C1KGbVh8DnMOrysUVoF8CpKZaMMAXtVT
4SKldZrpSRSkf2OW1PWV6PwTNbP7uyhOqOi0fLp+m81upwNZk6MNTaS3ZML1JpExfSxCu39VhfUJ
OXyzpIdRhJcwucF7uoF/gK9qRrFd6CC3BkbP3g==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Uff9H67WY6Ar2K9c/+nQruUm6iGjk6TppQf+oVVTgqexw2/5Vj8ARbZ+DeunEtPo7PVNBkWbx/0q
iOXx55yRxFTgSA2K3A9bYuLY3Z0Fgzkdm2CCArtZloxg2EvC2PQeRKkhOOKQ+Q48/RbmZy6gMZ7n
iYF987Be8Qw3Dih3PA7eiBL98Ffzc/O1aoBn+iWCOgtG7p0IbWAPoNyuxW0l5iUytBKST7sWQKmF
1Cta9Wah/mA5eGiMyPAMofmRIKW1kZuNpMJ4hBbVeMwVFTXpk9xGlZpBmJxe5FAlZINI/I8UedVa
z3FBU0dFq91E8fP4+pg0vYbSK5tWuBdZNEWJRg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 135744)
`protect data_block
PDgeNPv4/EN0s3/Oq7J9GHtFEDNAatKNL1VMLnDWteHb2tSwQvfIgZVKYznHDzfxy51YGTqwpLEu
tdlGjQ8msDW9UnsNj6xONQOS1Vk9KKn0qIS5H60wXIJULU7KhOtKg1PBqiMIEzQx5XzvU4e/x3Xo
Qwd06+qAERhqYg1Yo8Z0/X4ifuzbxlcZp0UUEgcq9od+7hw4mg+IjxaMP0HHMufAqJo/xsF4dY+b
2SSV/uVSsKu5x+UBjosGv8ZruVgEpS7Tfa7kru9PtsYUqjIZp6AUrcGmhX9YBjJLvPf39W6CYJuG
rEYRdH2vYYopjCDpBO52WecnOCxDNuvJX8yFR6iNJf2FvIKlM62+gnKwXl0pNcQa8lykDf1oT3Js
fIg0BLqkK62rb6qn8QrGhF4nOFCGYpD90QsyCCTcAXv4KEzr1kxJDlWKCPdhpZp1XuJzfTs48AXx
pK3i85HvfL1xOPFoAKL9k0SWt1PC8ZPivAb0IfoafL29mq7ygcRR3bOMuZi5iymd8045KbuRzdxu
+z7OyZNpDxcR/pjzzFJa+ZFK9RIt1LBg1cZ5AfKKwPd2YZafNlhuEjrky+awE/L0AaHemQQwvikE
4wJybvVk2YiBA/wUYcXfkWpDLRa9cE5w/eUHWlleiltKKwOgTJ7ihHcBD0hGeJ6zYesTC8bMW6oB
0cE6OKrRU8KhbgzY18kYHlS08R+nuTLye3XXOFGR6YWeL/h0f+RAnTfjedZe2ePiAN/B6/RJIE+6
ViihKAJ02osioA8XMEiKwOzSN4/RJrZpPjnB2pfeJVtz1YmuVNmk7Ko+Z8PTuL2WAndFqu/ivyiY
r44nJChfW0n1coimQV/wPvWbuhjwk6bIwCKRQc5vYH1wITDu4SZW6JSRlf/pGpIexw9bK56QbjVM
iETL/Yn4zmTg1tBYA4WjSjuQ66oLgXZuN5TpzIHnaWvnvEV0PAQeq0nlUY+l+xxXFLJzwHNJ3HQU
dZtSKWqM4YAljof1ES6x6B3NZOVI7mopy2L9kMWZCcqx7ZRYZ/oZJNf+08oKkSUXeUqIR+ByUaMZ
qnCmcH7SkcsOJjsBs1BgpWIdsP3djlBRRkP/qDKreLNs8wLLnmVLzYkwTJsLLsQdJZJ13Ll01N8D
It6FdCGHmtcO7sxJV+FxSxIorRWh65zyBNG1zMQUEqTPCScyDdASV78twro8BY4bDHuWNp9np/Pk
s1PFa7DM27Y8uX0wRJ0PCPHtIUFodMjzzJsNlN+H3Jq/3N0N9WlOZkSAHIJuLmFC0akIlxJuGGGA
GTDVzYvrmyVmQ3tlhzwY7AktGtF6DCC5I5ndzTUsYlT72AP8qye7w6u2bROJN6hHkSVFkGr6AS77
+pIw+c53Y+0OW8Q7cOVZ9sdzuc0DN+p384zdv3j9lLxwVLmxUU/RUmp2SMi/665YN5c417fw1KCb
UD2AJMJyNQ6yMSJ3AxUqOqPlkRVuL80byIcJWGd2ww+Kc5rtwRvMLVB1g8NJo66gFdtyXiEXez9R
l/LZE0/mmR4itD5b+WK0+vMGjPEuIsuOfXeCKMW4neUmaXOcqL6nd9CPw/hUugT6HWGFM059uTNe
CW4KilgBYyycMAKrPFf1pvEIyyfpeUQD9KEmyIJ4HUSNfbfFQ6dKpZOYvu0Z2vgqYj5cS64rrBRW
KGB9dqLuJIPJzXKD4v2bbegdDVsELxYA3Yo2vAMr7UreDSztSA/lkUoebi3MuRu6TfmCP9xxouY3
+P0LnFIb+QdxVPxfwrvW8Yp/UxFlSCc/9YOQBbKFu22vcCXh9OWs3umabbmP6ORX4gUHJR6DjMqc
stRtfLKxgcRgF1xFIMdsBDdDcgBP7XZx8RiOsuVGrSPpAe11j3wd0WHL/oSBHFl1rqTIjg3Gn7+F
Fi8Imv8ckMm+1cRbMnTlHVepfA0svGOtV0u5SKtLRZS+yMNrwK1ch9Uy2Sx5NPXbOe9tTJ9hw9mm
IZOr1E6+dFp3YQZrcCi0dOtGsrjWdGbxkOk2/kLndLXauRkWP5eHVHINe3h0LlX8jMRJOscZKJkC
uPRpJwOQzyUn76fPRRyr8+qtRTQbdINaNQuoLZEl4PVOJi+cdxYw2RX3yXoTn32lB+OL6FI5G01T
Q4q8xS7aparJpD9M6BVLacI/05zRVaFAiC54maVElUESGNqzybOb4ubTH3w5NrdyIBwEs/6xzdpe
2ZjYeH7qLqcnkI0qSSyP8LSRKEqdKnC8yOls7JBcBzvTmaiemCnL6TVPJeCab8nREKBEmf0Zl85Z
iBml98bpvoHlcONvgf5QJ7p7qHOLnGzLdRONrnQiL6ZxJOY8Ck5LbY7zdrYlDlkpzM5jc4SmD6Mu
FkBBDOZgjj63UeLDhpQrKOzhTOXDG+azKHLk/3gTkTaAd0S8xWdQMIhlcfB3qMd1rHyyB5TuY6RT
UQ7NSnKY+3L5Xb0zSfDgWrtVgzBPduvLpPvFpb+vf8jqRoBlezFzW4tuE/43gd4LL6l+8MbSVMUs
RDaa+TvU2Uj/mjUuJLJNzbmVZEEct/ukK+SslVOUDBzux/K+uMcKOQhU6n8toJ0Fp7ZPvMrDRNQB
Wu1UASaNwSHyabrs6v2VmcxvaNoSkcsCkPlhlkXMaBBIqLSH3y+qaqvGHaH+vmMizPhceYe5IUAG
MbsZEAjTwvM4tRvPVPt5hGtslYtrhiHKnGEppMhIOTQ5FEcn57OSFtagNQSS1YKn2mR3mz2hUWLy
fJA9QAR7Ygb0bot8kv5GsshCtPppcsNlkojrXZKhGN2PX8zu2l2gw7m1pi5VxnSCwDCry20FP10l
Q9Mqx0g1rahMw9gn72mvrBIoZqwqq1ECpSYI82jUekWFkDWigAwahLxWQXXCbIEQQz0IhPwGqrh0
xqgHR9rR33Y4zFSSMHXZwhLsiTQGWB2tbc6NYfl0DxlKs/BnaVKlo41n9GyE53Lp44r/HMIjL7Ae
6ytuL8CCgLKljSttpd50GqoEdchRf2YmEG2ImBq8p74ak4aCP8kdBgQpeAfru3SgSkocgpQFm0oT
zmpX1G8B0Fcl24GxzZWoCkn7M2NVgOsUWgf9ln4/ij0NSY6tgB6FkBPvbBwCO5ZEMYw2ZOzbdu5z
4G38shI2pMXCuiJUHtz6lGeDhCk0PR9rICylchiuhsUELi+YYB2q48madFdM32hYYtLYbxo07wiK
dB64kKRDxdDJgojHgmNb9OczonZpfclU5ZzIw6ctqDmLfneXCFDDf4DcmwYQVHmYa4rR5qTAV//P
Fk+y5oq4OiQ+ZI7lLj2Egw5/bR34KTelqOjlfCz+epG5k24nSJyfpvm34VriGV8XIYBGKwhIPShq
xIUDXMpIsWAIsZWnKZs0mN/lMFhsq/8DcW7a9bV9UyMZqUAgHttLZiIkR+3PJ3NLhNKsi8Oyrj6T
84YKsiXWARSsX4kfM8J0mGD/pMByeUeulngYBq66/OyYKWHo5+vL1+Q2b2u6UpIlOB29rtzcDo/0
aMBzRk8XglSM8emN7TdrFuPsUr9dmusGwXQ8YvQVQw0eZ5Ds13eRhCZ+Q4lmJYCmVcClSSoXb3FR
rdfOcfaKPgoPXREBVgOGpOkfmtSBgoTMAL3cesyFiXDAdXfpMWvuX6baL5vyrr4a7Eb7mbnZ3gTy
GlskSxrZQ3jR8KuyzddapEDqJhVbJEZxbW0SsiqXHoVTyaHvmSQ2wGdZizxk+mZpmYCaAu3Pv5aA
EviAzGNG83MMlkkv4/mqFwNe3Vh1/1WRHco4+tI43PH2UqwywZGFXOHR2Z7nIbrRQSRLFStDgFIK
nHwxJT/f5NosVMD3SqmuUcXeTPiIqwIzcQX7K3/eW2/Q2gb5PXMHQR5Vr1ey1xWvYKgdSn8k3MCP
UhxLQYNZ/nl/RG3e8miFmUPP3d/JLjto+rs/t2LjMW7zo9KMhrzwcWNB+n1s8l+0w7Z6QwogUoOe
Kqfw5OEoMYGMo6fjkx0tRG13qryMMUOVd02nDlgiSt12ulwguSVTEAivJzmnT+1Mh0ViD/jXro3H
3wNQVoDZWgwiX6uGRsJ5vbhsKvtTxc+Og+4EIMYo761JalmyEUeg77Ogaaot0FBOeExNrFAYINbc
PrV1RY1+tu6ibq6HwayXQiPjJpTTEOBRQnqcBuKY1eeh0mtCkPoEvWagF3rnP8grwP+f9Gxa3/WX
d5qTm/E5KNOtJemBd3zSNIyGVHK/gwabqs5Urq+n2PNg9WGRi6ouqOn0BojMalgW+QhHc6y+yd1j
PpERXu6tup1lhb/WbHZ+tnue45KtGXAM6XF+XKWOdFbcH2YVcl1Wjas8lmoItt7/6Lf0vMIOkllt
LC2vb6UOFeebHxVn9m+Lkm2l0UFHZkGDCsWBENTv5bXayrP8H/pzqbFNiSz8SOJ+Li28h7PtPN24
wi0m/1W3Dmejk/Cz2T2ztL+B2ce1J3OyIO4mN4vz7xDk0TBFGuuEuRCMLSKkvMTk+2Hv5UX2vXoV
8RqQE1fqUFwgvKJnm9Hl1x8DaXQM8r9REBRhCrGSB6mo9KfCO3fSdKcjKBsIqWRwp2Q9lh6UlRIy
oieI3mfqFWEJQRKWSbUVS3uEE/r8GF8RF2R9yqF8Oid0CC1xtgb+ZWyqlz/QszeBRcNoCJmBj/8X
/XEBeWoMSyF0MjCR+lSpm0+mv5mTKrnpLIWSDIuzA4f64/MlfTseMMMkAyAeIL2mhEsd2DC/7wG4
RdmRu/oadhzNd0iFRIPiW3xIXu5WchwXHbySvL1NG2Q8/71wLwgBl3py1JC7IBKzzdAWE1fceyQl
Kif3KdMXurdFct1lq6Xzmft+u+Eo6mRwK42TxaHDnA99+RrjxV3wnZeorstw6hNHgkXdbca/T8by
+jt8KWo97PlyOjCLRGDFqQPouQNayKYAoDjSHCg4xgy5fFONgEiVUlacfTH/i46KBHBg0Wm5AD8+
zvG5q3I5apoOPUMuuuCrm1rSaZxrHZOk5YPXZad3xx5M7ruGKC+E1ZD9ku6ykZleRqk7zf3neWp+
s8O70uTaELQh8M+SKsGksCrJREvbAKYlYZgPrVzZdjfnDOuyiJ9/6BkY3S2j6b2s0aKucMF0fsQq
izrsBNAOtGHmyM9WPChTa1c794zOGf1FKPyy3dBi6Ox6iu/8McSbEssvFZjL+uuV+af4JTbjsV7I
42Yf9a4lizTkeykCG/HtBMUYW+yzVYKFtT1LaHYu/mq+i4+Hf8YUjmYzrDcFQ3OHGdLd1qfNjYLn
3Zg0dKIJUiR0lqLbKgHugo2GqJ4oQxnB+eKCVD2lXoJyZ8P5hBwZvhfxDEVoQWyA8T3KsNHLniI+
xi7wLIaaoeWL5Naqy64w2mUHoE4mHf6Apzpf3i+cyekz3P3s5thJLwABUHn8TB4o6MqdJ5hq+WMj
30ZPFEYzsdPSRWICUk81tgYx8ScWf2GCk4A+d8Gc9R4A8VtN9ClsDQcJ1a5yxG7T/xOu6zoKr99y
wsSJJmrnnyMWG1PeVbjd6QYE/0z/Y5NTLjp7JXpQDkv3PxarkLKkV2KHJ1T6StTSRloQcf1hi+ka
0PXE3eJ0qvBCMZps+CcGKesfSWB9e/esfc4ScQ9EEe1HlsQwcKSE/coR5Cw+6MdVf7mFeYqqW6/8
MNnM2AXBkPFkawI09X8C3c213UXm9WELUKIseSn7zwYuUiIgWy8A0C/yRRZr80YjDDaGYuLDuUVV
dQHWFBUc92BVBIiNsJKuXdpw8zmIDjYT50qPTk+wZfsPGfdDqZLnk+Z1uekWjyjxLbdPyQCV5yp7
V7gzN1Z/5XMN74n0odsEWybpk5h6mpnZ0kruIm+MvuTNY6uBtPxXmZounDlMYq4po4WZ59OqYkgx
dR8zCDYeHIa3PLD0qfGXknqRr8C7Nre0JbP/xSEcIjRRU2N/AR/y8YcgPwDqgps8UYMPuTjhAe/w
pJnbFzRFDfVvwhcSD7SlnNKxVHXNGIDKZ4mPiQ5/udzsWIIZH6QlC3OLjLtQSVZBT2BGhqgDXsrl
7ogNbpjF7k9PUXZPJ8dye82ctBKBX493nrOKqaBs8X3vKCrr4npaV55K0bl8Z4flCYjPhWELuJ3U
P8yc0WRIHFDz4Ep2T2ZDCf44mnpN0IfvKjJxLcxIKDj0Al+/qTDo6u3m3aj/C9c/Fl8r6oR/QMnO
MtzAnGLeO8r4DNPirz8+ICuLy4LntidWGQJAUhNIOjuKGk4ftuuAas7WRRVNMJsj9dXAxUS9lddz
X+x6+oi9N69lltN7lMWTLmJ0dMuFrSRBg9I4u+5Gyo8jdwA3qWM/9jHwYqHU3obObBHUvrxVN41l
9LNF6foQZSb5LbUP/nBQenhvJwuVEBF8dVAfJSrVbnDrfN6cCBQ4nEZrnxZ1Ibq9X6JZCXEA7wQf
DzLzb6oWqbeytv3Z1fPS0e1hGysjY+QLQ6VXNI9p1VO2yC3zndFyAPXgp/NGSC92sZAoH9kWWDiH
HEgkfTG3L1kVYXGcyIFVYLtAOTaZqhZLLKFyi3iGDiGcGgh/5HRyGq+q/R+ASuk5QobJGBBBSXAT
W5u20BSJNulOmv+fYez41vsUyZZYdfQkkWlL9Bb/Y3YrUizbh8ZVohkW2X2XXJVXkTaheFwXlJlD
yLbcVbQEoVhb9DCS0OGD2GwO1ZFgj7pZ94211eah3ORFT00td0Q01M8gfsd0RSmga7vECoL8P9n5
1DTc5BFVYWhStWgwZ5gyeEFGo/8Uyac/To4jRipcGaZX41AIWFEviazek1nB+DzHirQ/WJNkvDIX
GR/m3XO3vER07Gl55etMxSTakk2j7wxT2thX5t9D8ekWOTrg38/Ap7A1MbXxlHDbNXb0E57/MWL4
g89eU/cU3fmYsJwGWCgtAcIdOsZ9P+Qr2tBa6yAfPXkCpci+n2yglbjjS4jAyZC6+6SJxrpQaAIS
m/uuzCIqBDCh2LKGDKiDVeafcj976gXjZOB1N/k9DnDyI+M2oz+VdS+GaSxwSSVI8YHpVgTecZLM
YjZDq46S4TJ+iuJOd9wtvYUGFo1Q/RptambfFGI4ETdOo9S6uUS13eEolr6Zko5aQmeJT+DQQCct
QAEJmH0ljt0+BzVG4cY1R3VV04jeUvJwG6/PlFx7oqZxk9rQI4f99nfszt6nWyNiA5xoy3wiN/kt
Y6D54I6sm2M/0jWp0m6iMLuox+oIG1p5F1h7xzjvYlq9QwtML+qAvI09TCZMxwjWWlwXPeqAB9Tt
igFV6bux1uaykSM1Ol0BAMCKgjqKU9Px3DeotXkLJIyLjhLPy9UV7ccbGpRgRy90uHhMrU5dE8qu
Bn/30D6qISO6wTB/j+PCOZUDD6G6a26N35oZvO+UsRXjnO2yeB3bXZQg2NpdsFKvoB8Tnd7xwmAW
ezVZXLWR+VMahCJQ/dCeQ/QIVbOdeVRDyujUdSUL5/HaqDydhTtW4zziMENz6S5D3MoEU6aQq3Qv
k6zmAOGrAggEMvMYFxBSIKDAuVBJI+Tf7Gy//joklOsTvSWEDiOqljzkDx7VvT7XhuPullLjB/pj
gfgivrnRUbbr03IH0v+8pWKJato2IK6BXEWdeR80xY+SvFtL/irnroa9mfD2UjzKYRAj4qOZFnFf
RsWA795zDLiCnLDwzk2xSBXJYZAjO7W1KqVZfqeTK/XPik5xT5EDJ2+AD7MngLzhO/9YgHry0f7m
4pKN3DjowU2AgXp88bXOseNPE9+N1Da8eWserj/v6PR8FiJgbnkN68luqIKQlK6WU21q6NWl028X
awjeNPEU7DH9xatibsQPofDGtyHF1FI59Yp3zfi0DenZumr/ODkIhNAicXa8D1xzhI6OzPdRyifh
uSyG64Jpy0axoWiS+lZtvWqTB3ymLg/SgO9KkXsil/bp2e43J1jne4oSPO5Aml9l4Gbh0Tt7TGE8
nGK3N8B9aihYrtKbDyomj2xlbE01atDP1oJEiufz78SIY1Mua5pbm2+bgKqrfpe4DHfqEnpdZAtL
MSUDOGWSAaCVWgfYI3sw7OamIZV3NkJjKpZoRz3lS4VYibttViSIa7fJrDPx+uLv9VHFB5G8RpPi
GbGzGiMwveFbhtJPjJo/wXRPOX/FhbNnpl6KiovHODUllY5k731CjfUZ1Rr86OhffmrZnIrbWC9l
toPuvESpuYnlpTeCMcmDxTEoGmcoNtWLNmyg//Hyzjiv0iYnr6XFaKODrrXcjj/VIlLabgQk5Vn1
y75YhsjlNTKPqxv4ubXSPkF66BIVCgTdyHk6it5vvuNKQlJnKjUxqnjdajA9/w9ECa1uC3nvvYnR
qYmo77Wlwzkf0wrkIw/YXnoLbSRvun4iaUmgCfrJSTbRqNua67yAbTbA9ypbKuBfjU8VN15gUJVT
GSA3erbmHz/rLM68PemYUbc+TrAgVg6yvHoWvLROf16xDEH+zvJAtQgSU8RUDaCoIvH52N9vMLKv
Ao91aDLq07eS2Zsl3ZZ3PsOQFp/1YgEtP3Ztj6/aVbqrZpumTFwolLF8bPWfT4/33TJpTYr6lHJG
+pqcLFOuorToUtIpZxXpjZUTQkNdWoFUi4cBzoe2suLhkIKX07rFdy5eW6voaqI5+6PAI4Uvb6zc
g+P3MkhyOp/qX1KK6GMiLPYRcIi2cDAVgWnMN4fBrEzmoSkAlYzO41zVS3mR+aNat0nMTvoKaiZc
UXPIZ4mGBs77FFxOsiLzlS2ESYBJ9p9nv4+AxGSRQLNkWutZRi6eI0/T3ZlQDEkFn4d3SbpyF7gc
xcNSjZjFemJJwBsHYMvE9IZUl0E6+c6Tb0aDTLCz0bYgOmTDwtmb0xc/pR+syC8QzUJ9HWZprRMi
0GGHKHZtEJoSJtmO3qwmfrlykNKsU8Oits8swzd0osgCXOBGH7vBNCUdLpZhKjYCCz/icyli399L
A6+DjAqKnFW4Ur60FUTx87OyQkolTFWDyZbBgz5byaEIWLYtLYtvpB1ljT153QBQ+3ba+oUkVfxN
iOehJ1sM3eUy/IYdzaHWgLwI8u/oAWFO5IMmopLeAYSycSQweCbzHvDIQ3Wdo5pxywViPDe4+XkG
AS/Udxa/UL85QcoIRNaKsOg0z3/rC+ZG7AoCM58vNffCmMIIQu/bSlm0ReJms494CvvjK9Pj3pnK
xcHvIRwKW3d0d0zPgwZo3kOAHdqjYIOOhNzyqrIBqvqLbqLXsAj3nvcY/q92G4YmRCxVdU2E7aV4
rRXTiACoAistTdjUXbPigHwRPVVfpxgYn9HewGxwypTCem9Flq+Dwl9Ciw/+L905dqhWJ647QGpY
vyvH7Jx+PZ4Xn4b0QO8njM1dNOFZz78r5y3C1IyYGGtFGu7AbeOYX+U5XI932tdfH/B9j56szmDD
zmBprDPPKMW8NC49MYAsiF4y2izh4yLAl798tsFNcwmBfCsBiTKTP5bhj9RwNfutDUV9mBNHlaGs
1C4DFBk5DpMoMevHhsWs+b4zM+oeO7fI1hj1XncamsGBeKqfAQwRraiNO5HbQqZTMzxOkTVKW6T2
myIVe6eUqCBZb/7UWldFvepPkgicleqTcrl1KSQ4UDFnTdCdjoRRIguMwU4ZtNZqJ+kFZiG9JAC4
UJzbHPvmWBsawapZ3aOhrHskLQisPXFTRNOk2b3P3pSan4o05XslxO2xTMkaqGwmsX+ydndEzC8o
fHUV1AL2RkLkKwk97xjFul6Sh2Lf2kfscF7zeaIKg1PXEKdBRhJkzNxvvqMDhIoO+qxw2k9tnEnn
TNAUxI+KAm3PgmkmLEQEahrSiND2GqVD5DzKXposUQBN48pNEhya1GeCVk1VR8yEwekQ+o9IdJEN
K/CgWh4Gcz9rTbv7VOrRhDHD7tMnhOqpGIqW5OhfLMnXtTmKtB830/8yhs6zNZpk5e3QIE9d/C8P
y28a3i1o3mQ+JyyDeui662dzsVasg1cZjcv27eIDvVt723PCFR1Gwiud17q9AXeIreqRt5yFuhV9
S0MmPpLkLKSJ35uPE4gJkeRnENJYHmvx0Ht0nx5U707Me+RgadEGs4ZNzDznBOg8GeJuCNGXXrs/
5hHQ7fc64YHFrq0yfLY/7CYWt54DY9wmiAdKgZ83hOXLRvRbSDgiubclcgT1/9RjFC7FpfscZDp2
QQ+4+XKwsJJOTjdc9Thza4cTuv6P/0i8xaEZyDhT66m/KMH7SW541vYPL9uzqUR9Q/x0LAB5zHfw
qWsXbJdM3NR+fqxg3xJ0aDzmr+ZAPnBam3iDGdFMYDdEbwAThaEyi7TdIZp7kZzGWh6f/JQLHB0k
6Hiti/YPKAjOfZjdXl1vH8t10Lyl6/SiITWPdif02ec3Jcun3UeK2Fh0auycCy4whd/VkjFpCKYR
43ETUaat4f7cwTMiEDxIEUc2QQSXcOtMtcDFJ50EVEfOII4QgluuN7tmjZlUSXOSHLp+DujPn93l
wXktzpoMzjvCyd4cX0NM0xKM5PacSEAgM5W1aJm307YEyg2PrpsQTPh1lcqVcCSHjRNKQ+wG2AA0
hQTdrmSe8NN/43OD7Il/cm94Z5cgNhPlw5+z3NqIytKBNwVIqEBqg8ReUvMkjc5Vfi9I4srXVtsW
SeXB3r77Ya6nM4x1zFiiN9yZ0gRGtzEVmPCneHiYXboD4KTXPGDBWouSYbqrOu5fEmKFY800V9Pt
MEgDJKsODCZ6dHfKY9AqKvFtwwvqD212Ib7+dsXlGfd5/smRdQRgMaZ4MYMXH1mqFxuYPSX2iFPG
CgQ2XOPj/0Wz52XWCiN8i/RvvyGcrqMkNeGpkreZSitE8J0LbnnKKOWRYQVvFBPr940/RiTTVGka
YbEooNUy8hFokIThl9ziPG1fzTVWmNMo/RB8G39O6BV0/i02CBewcqLDsMILVJyFVK4pQhx8rhRl
o78Qmv3R8ypmrwyaW1H5qzPktFap34Wv7zO3heueoLCdhBm9IX9R2MLUdeS/sAUcZmgizDSB2V0B
YojMviE8u/5OGcIEZi6mu0hSh9zdYo5loTMCF461fjY1BNIk12tfl/zuL+S1ITx3GBKSJ2gjHu9e
DuBYw5yJWh5HVkesLTkGvUTbbklPpNU2CoAD8Yig21rsr0t39S2sPz/xa65VH1YCFF4GIXKSgLWS
6RHrgp3iGuO8bXHNqi2UuMTrXTWJXe3KogE0duXYBLEGSJh4koGsYeYYZoBQTUqv15St6aLdCD26
cEjEp/i7IzIMdTn71aBWFyeDz0cO8H3U5NCi81Svha97iAe+Q/mq+tacROg7gDFSnkAysGTtWvpW
4/Z/ey9ttVdxdBuAcM7Rdr5kxe2Ld7ix9fI3AKDYLlqcGLy+f6BHiVIzfQT7l7bJM2NfkyHymWGo
JOxjdjsGr6o1XruXX25ZoAIyExFrOmV1+HVoqkvGmxxvBDnwLXhDWbJc8RkRbfzJhy8kKPhXFFtu
6eGf21VgDSrHj/USM8GAADaqg4VCupKwPLxTInwhhXY0q1CBsMBUkyzUdK1rs8i3JrCJZrBpDg2o
qX2MkFHGzGEWpSMkmkAQET8CouyrBoKyHMtGxf8BZLqyKOkYN7M6gD399aXDAPf/8lVYDFBZVmUb
mUn/jCCSd8rzWc1pAFCao0VJ/oPsYKby7CarrKyMaEKH1R7sNcJRSr/G8woUG0/lGBS5oPPm8fWV
2adXuwdUdpPSddYBqHfQA3trf8KrmeRgLBecYgTcGbi+WrOxTSJgpOkjnWEPNUfwC2Su/LP9jWxf
hs5HnRozICLeBsLbc2nFijPSI7Au2IZOAnXlfQuGfWQ5reM1yvhasGyaiC+phfzTqsb7q1oJ4lkn
Fok4zKZKWEs1j7QW9UvEXOnx8oeWOOQiNjEoy9gxl0qwi3+DgNtRQ6E4vN7/DvA6FDyQ4pcHZb9w
PcgSfSI4M1T2DnR52UuBGuLmZbXY/j3Yl9S8oFP+e13gWtYsQV8u+4RgwAxRnT3q6aDi8hF2fdgk
WL+cAH9cLocQj4AISDq3Nx7TmXNjIFUs+iJy3D/kDnVQCUawUE/dwpLoNU9BeyvFIxaBj8P6uZmp
nXK6PKwzOOJtjTaEdAGR8FM4ADiE5ApnwYDzq+rvJUxu0MBI+8QV0tPzrFhM8TxaGt/uf13XONUY
INeZU7i2JqTe6WvXVXMENK37fFP7CN5FupvngE/4Nvfx7+lbEQZG7C5417+/gvnRZAuyzcIeCVQ8
0h5luVmaJonrMzh2wwLuODijYO8+vKP9Q+Jg/vWparkIFtjMEv+UTqpKQx/McqmgatjsMXJcQslZ
Cx6qNA30NUcilF5Kdk9qdt/orbWnDbB+8Jq484s1J69x/vyqinEPFlbM3p0x8UlACC4a4kAa5Bgk
xSfr4ZFwOXTZVXk77/HGOBVQlNRQqzB3CLSZ+Q81nGklYC2WZAPOrr5fCAm8KAMfWS6lspyencog
DNEJl1cPiQChuwCHQLGuJLlVFNj+ktTgA91WopfHVvV7ngXh2c33AaQDoYFvoVXT9S2sCGyJox3b
ek9JDKWTBWD1dboo7DUPHEviR7qHBaCQZ9Nr1ERgSVbO8FptvN6pE+WM45TMu4CMuvZTUuvQ3kU9
5O5TemneYUntbi4J69WPnjQlXrCE5w2z4l63tjqnWhtE660olNifzxGzZZ9CMtOtsAxUOAK/+dib
I7NlQbqz2ZkOemS29CX7hZ77J8tPHw5a7P4iYLUJRUYBCPmVLwkwW4jom4Wu4Le5R4wKhuE39Y3U
6MZ7ZWfX2BbNnvc2QUkJS6jmlLGJ0N58h2QLBBQqb7sFpCXZrbXJEaDdNGDJGVD2os94mkh69pb5
hWFtFHVKXH7qYEgmNWpIaLSQWviXjfQivLqPsYgeUvJLbghg3h2k3eE1PthL109yCNJkhd/l6oFo
QBCBeYwKz33EfZudCwzGlUn2gOO9quPvTma5v3/qyElia4Qy5hPCf2O6abT+a6dEGnW/7SDoL97/
L9F4T7ziSuN4d8MQlHsleZCbq5OImaqZgSp6f9xosJdWn9fox+4QNCwO0a0te3x3y3YkdJDQ3g2V
p5g97GX2qe/pcEJhwnfMFqjgwDBTPsm4CQuJul3Oh4SgC9sbVcNelSCsU2QLnDexFytssiOH4E7I
xMJAe3xIexFxyhlYUjTyDixh8DPRqwj1NwPAwwokPjAyUzwWO6pdxGVKEIZLG+CFntjggpatmazP
obA4QiTc9IBhqN+y8cjTe21N2qA9KNCVfj4o/bw6/g8pL7Tn+772jwLe7iOoSlUVXzxS4vXJAi4q
A8V4cBE5RAcaWNvg0fgAmvOsTedk6G5Xl37GxndRDf7VEMLrkyQ0BG6zyVZPxA+T6RHe3iRT+ugb
noWmWgsBpumoYdgag4ZLNRYZU1mV60HiegAfVosJz3quVwmBZh8tZ6eIEYxv6/mfaIDpUooyDLLN
Sg7Vt0oqp4hxm1igAFGgV8cUxDKtc2CeryHz7qQlw9DQzcJUtU7zX4Pf5q6sL/lnjTYzQNYbT/10
FDLvuMl5iEJ0ibhDJWO0A84Wgbnv8g9SllGZMBKZnVRc7Ww5m1V2GVdieiWsGT3hkzgvhhCM6U5U
kxmVB3m9aILKgF3b4c+GgVQprEkijAdhnWhd838MVooR3+rnngmYD3Zz9xehaHm4nL/Hz6wZsMFc
AyoIciFlohYDHe25R1WcwNj4rHEBOvyiK7hPCXSdrTNDQKNUGTVlzNYNGu4RzfFYpSEO/rwbItKX
Wh7YXJS0tGj0cP+ksIsFKacwfDrVbRYM7NjAeB1UlgePh2bGKBwVEZsph1rFRJh9AaAAepCtQZfs
YGq60manYV1VIvX6ia9VfIPho/e1OwpVisS8MOK+t9jYrsFArhxR3dybw6Bn4MQJhOOfv6RlyzqT
3K9LoyMVb/g9YRsrwaDP0aC1qum7bxL8zgd1Cb8DejgIDumIMPaNj9VuyL1ndtfOk7mVxuTG2i5w
dW1AMIuXcoaPo3sk3Ecs7D9DpzuWNwCNolVD0kW67Ubk4s+qVQzz0i3X3RhxSlk2e3Cx1OYDh8y1
PSgpBESbBvnGa3oBuykf4dS3bAPyRRiAXf3pO9KvscsfXKiCJbb/sZU+9IXPitl2NZECvCeq/ntx
Zf08pYrAqY61yfqBb6hqGBBI1EMPZasvgO8Pbx2WAeJjm8Iv/xkU/dLXpzzG87uONea80OwjxI+n
KkVGK96BNqOJ+3RgCMNIFo+iQ+EM8yeMOyexO8NcY3bTh1ZwsFsd6FIX+Eu0V8/fqZzWaBR2BjAK
nn78ht9SzyXL8xhop9vc+6VWiBh148K+LZmGoJh6Kz/v503ESXI//QKr3RLspm9D7krr3lUUaYEN
zfoOIaKb0IWTdXHKwz8GSqKwGiFuVEKPQsDupzDAXRrz++jExbkg13GaXF+bgUBJ1aBCQViwGWOq
gpfo9HbV9u+mLmfGzozTZnnJCCifY/ba5DVZJaEKsrqH7RhfcIUqRYezoUHRFd27cddRbIBKhWew
B2pnx0uJJpdQOtRR019PD7fbMRkcaNdZeIV/PNWX+Rx7st9k174vCttOGaNHUEXHtH3hxKzQb45x
Ya+zDBj/KtrEI9XprrL0jAgxGOV2ltzLyAUQJMimNt+OkUyWNoZINW1mnJfW7W0K1Gf6paUyjxxT
19Z+qJD2civQyiiVHMbmI3lJfFuu3N6/GF7LpuYC/0XK9pAU3CU3EEIUiujk6h/iSSIyfN1Lq4q1
BqjIKI0dgOt8xdJBEjofASy13AvUDsS6vJQlc4qEmLVe8cGhkzA8ukTW+7ElBWG/dNCDz5jNwWjq
QLuva3+RuugLNI0PQ8v1M4EtAay6i0gpYzX7x33h01cEk4PLk2lok386Bqd0LTOQzHNgs39xQFlx
YwrnaIpd3PQb1D7MR35yyZwhyLPkpPOy3jQI4OTgWdlaLQczCRUoIecOzU73v7kHX2dRdJi86+ky
UoHk86m5LLIbMkouS1fC1um2exYGL5esq8cxwtHmTcttEFCySh1zuy8WfAUkGbOYdA3Og+Jx/d/K
SVwTVbIB1Com2XpCZvqOVW+xvY6yqk3tNW1sPq0tEl9FO2g28zN501ihdxgVrcsya700/0YzYU7G
LNO6vsWmbOEASyNfYgxr/qVv13Kp0oTk+cyyi8rXE7ot8maD0lYREPOk2mH+r3GcFaIcbLTHwuK3
oWML+C3X/rfLoSy7+bLLfiOD2PeazHIszuRFphiTM2yySuywOnbSU5BnrciuFVF/SuszNvOftd8x
s24VAb7SatanJC2Ax2xXGJmAZ5tEzCFOrKva/7vs9O8tnss4Wp0lgcPt/TkzOc/IVDxpdWPHeih2
wkFXrAxpaH6VP83JtLofgLOuHVG6bvYMyRNcddy2snrfTZG+hOCH7+kmQpi4vpicxwwu+7QoHF8M
9k1XYHlwx3fTXVlsLH2c1sNQyatfwmb47mH+uZgeo6hOj4zuyeWd455UbKBE7HhT1ZTKryixx0ay
qr6hiqgK3lHWqPAv0Xdi/hqPvsa2xP3kyab9JOqagRrYBN8A4nhVVTOEPTh1pJmWzQ8HJKnH7V8e
AVjUxH+be19e+rsgviv7rMXc0riWgG9oz4gAzC4GcLS5LyhQ1enj4+9clpJ5kntQOZxM9nRASOna
oe7vjxjCvLF60GyEKZmTz28ODq2r8pPkOdB1kxqYX3ZUU3BIiWIYP+BA6AwoG9F4lHYN0H90uSh7
h7I+Fwlo7rH8GXnS6jHSAf+7K6zjTB4bRyc75O72m5gbZFR07H46/olu1jIKaz0hzNW9OQhEUaEV
xdZ2FVM/622oqnKf/bDQ7JmSF7LQNGQ4+2f0Qf2hWrCyWD/2Jk0zGG7HqmuXQQsfxHpITTogPdKZ
pFGEqnFxwup3rh9i0bPCU8ThfAdp9XcZbxB+BT6VY7hzUpjSd6fW0NLm7aURYD3eOICKGWuD0i8n
R29GZJjrae9AowQzevBYGdGse0s1DbiNDSVNlMHfT03v+QI8pzdmjw51CQHR10db8HAK4pYmXcjX
jxcT5ndRQMznurPD2SjnZZwSTQA8gF3H/74SaiFFPDf8wEC8BFul9gnrTvuFwNuzxqxoRt4ugBlV
wjp0CggAqUrEV0UfzljBnYMTEas9Uij8S2jYRDO/dghmaPzndljQdKCQ7Dzx6KYquSPcnxLU26bP
cThW9bGPl48a9MDfWatxls5UdcgYk5/vyV3CN8u9MjvbprRWOmPhpkPuNdfzFx+E5nQXbR8KCIml
MvBKC9VUOX9Irsag76aJZUl3EcqHpJm+/hAS3zZMWCzGNQGhxKLxJ+tpceKFkO5r1xMatrtORl8e
7tqBa4AVZJ2vxVg+db7Aqb3QMsRN9mUVfdo2BYnJSabdxILQboHtPyqyg3di8qGKeDsrQZEPKe14
l15fIvSXazxiD+FjHGCiucecS6TgKyJpEdZyhTE/ld/45iY4OZjlgZSxoeJrgw+Aef7C8Y9mPpSv
zN5SavlEurHCaJsQljQZE2m9f5OF5R+SJylnJzPlRJdDbpEInCdH2jtSOM8b20v4DemDoOTYC9Di
UYtzEEMQe/2vGCm+fZVyJQ6WOLOS+xqibD3ARAUhCjeqmioq3Z3oFkfqPxUrYW3+MohrucAfKJJq
Tj3HkuMP1fkt4veORlQ2VtAwYWs1ZLKku0dZOErvDjGXk565T4uCLG434OmbO+jcQc738yhdOJev
CHqUNUq6YtXQoChYgFbbXCtiy9YwabU8QTtjoC/NVf8bfdmJ8vzZeqBUFqLpMaxk91F/e4qYU/1M
SiiTEfihfyMOLh+KPLjqpX0PUBpoTjS0mYoYNk2IuHMxlngieDdXODK7F1FDMLVw1JanUh63eRGB
CZhyawLyPUTNE9iGTrlB6lBF6Ta4WCPLrO9A82FvkEeoRM8NGAgZLFFajFOQOpXZBkfZp38ljkJ+
EimMwURdf5+amVR9oC1wJ0h8RiVJ3VIp7lQxcLtKI2xFZnm4FUZA+/f4yYet82BSQnw7U+tXpxiz
tBvoBglVxVZT+MRBPj9E7bgc4FjpBYEVLtx2S4EDz7YGZ3E5S1EMJyI5x4yG7TTFQ9lvk+e8s15T
yKqM/fqsnjfMk76YBloZeP/tgxYzoRVBwi/3EYyNg00ESi/qKl/RV2llAkhi2ULfi9d9MpixfbNH
ERzAv7FAQyWTuCwzlMJtbLISjDPimZpboq4dGZwIbvn1qv4lHQnDYgPWLS2M05lF0s7Uc3B/b3H5
hAlHyQK29e6oCVeXmOPGA/q98h2gTKRLQucizooHGA5JfBe/iEMaFoFC/nUGqUFJO1DDDX+qifgs
AX31siYiFRI9i/TQMuAxQBEg0xHWVACXjrM2exIJwVFQPUllEnp/cE2W2jbKSjZQMJBwFCgJSC1j
rOaeu/gIVedzs/OAv9y/cG2c6H1jyZBNMp+txff83UU2iHJdsj8fDEIkmFEStBPlsqzx+5GOAYVN
g0RC9Qzk5SmgSt7HghLFpmi7oKs+B8e6hnnmOr2iAacmL/R+5uCrKeA+tipfFZiHQXAIwrNZ6pnY
0sHc8wGnhtPnk1tc++0QlAVGgaFZuKbGNS1WyYTy5TMG6eyzykcFWm1db59lGrSIkZD91mGUdJud
0tiOBx++h+/CY7CdXlyQJN9Y5KURwmXiteiwcRoqz1HsgRgYbEZx62ii1ahy0tg+6//dN3eC0inZ
8nRwiy+PJxbFssv5luZNR5zGZ1KprZOOFWcI7AEALsN1Vbk/VFtrHZ6kyfcC57XLeDDvTdK4ia14
8j4ZkBtzjtiBjiIws574zVnADcGUDPJrFp29ejlisxp8CtSnu5WwSRqbv0cqU0uKToGHMbWKUytG
SbcHS8D6WSzRLOhQcmcPja5R8Uk3pONYLC0fGUC9DxxyhJFbANboYrZiqGkEAonYP1uL+uU9h07V
+MKBqoCG+QXlHtDyi5Ecx+wfCx/cTK8dXR3WFsNiSdE3+Dd3GsoLGW6UWo/YsxEu82HXyvqF9hef
Gvp43bLa7r75VDh/l8GTGkPRbRPD9e6qRHyywcwugbB+gxq4GcP404qcqisgu6YBa/N1wmTcgsgd
etXtLJ2Z0ce7pEQp4RfyvdJweCkeCpiHAfqLM1YT9k8jgjg6+VF3ZxUgxdNHy3AQi9FEUYB2SmuR
JN8dvYsCTr5Mixm5f25uQhUY0njI6pzw1IHG9wE0s+cvgTgQ9TFcVrg2YTfzHrjwSnh5WzAz1HtW
L/ghc2AmpdXnXUUav0pcFAquXco5HY9/Dhe3LaoMOfFiVZt5E9J4pp/7IQmU0TfQwzKC48Lyiv9Y
bcSsX0LihNjQY6kLxM0ZJCMK6iwdIlACdzOHn4mF6b3McYdjV6y7qE+bUYFBxXBK9/7gnTvrgqMD
WDS+3QocydD5JVVu9ZlYQFLxnK3uynTPnSILVgUtT81px7cMVEkaEPjfPm1WFAnJth3MJ7akAHpi
xRw0+bX4j2ma4cBWtWOOb7UwKcObwwDN2FH6W+P6fgdoebdc253bwVGIKS1iPH8EUgHBhNw5apj+
A6uNhy4V3jGqH6kXtbGb9wtgFg5/hsXuNh3Vscib4Iakzhshbr7hdNqIB5hgS/FcSnSgVXubHqjo
eA4Ukz0VPhxiN/W9oCsyfY924WlUMvAspgVBITgwsgqunIgJ4H9wbuwOW7FPwGInwSXNqEC+NU2f
/mc3ScX8KGKLolhjZOwudO20lq1OeIIUA//NFMRxkLzA0APayMLizbHTE0+rVnF7uznEYZlIxk5J
cOW8pYhknMTFS03MNctrCh+UNMmPaYBReoJ276TD73hglkhonUSgmImAYIMAcw/njJ+hCQYGi4zo
gixAyQdtQP+iel2haxc5CJPK4zhuCq0EH4/Ynz5BMj0pnlp51PQRGA+yw45mFi5F+1vc8NSKBCLB
lEaONCyv0cTDLYn7/yXzoryS/eMJbsUBlRNyTF7i+vSalT9jSIMD4iK7IhehL/eLbBl90tNnbgFD
NO5WRJXFSf88hX79MZr9XRB9b79Za5cOrGweNgkrQVK2ipfuplgvYWzeZ+mNocSgeoJ36VxiIrlM
29VYZy3/lv3e81B83obrWk887gqykp6qq17ro6QeHGRjxFhgP8iUda8g1T0mfgxMBRQZ11ZFINEj
PxTlRgWv9QSoJrSGOOBmtXSgzZfWmQEAciIPJmSUYnMJsCyXz63v/JookyP1COlTr4xYk6gwus38
IHVPmjMNEgxJlxYCLdRM2b+kNoEuT434PGCi/pJt/3w2ogbhO+3GG3uR1wmPzNDw6cQzn4AJIEWg
GIHSoGPFR6y+3Vuq2QBbuItWDVLmbsZjO5lcGjcGWLSb9ISw5Re/hZM6vcyunzWNJrSOhxoWL6BU
CS5HPRjqIq9kbALpy4O5i1G/hjcinrOOTTCAhWCOEMOgY7pFU+MbiY9VCMtcDcZ8DjTp5dOLMVF7
DMUI4dFxyflJ9g2pgEYOBfEMBL3cSpE7gDBaSxb6cPDdNEQd4icUHS6fVPlC7OGF2LTV9LiRMbVj
YCIzNn7J4dNlYI0aiITACrUhy53mkObwCStKIZj3qTGl+XAayiVUZIt7HkkcqGKKJHKJXwlIB9fp
2w02GOLznvfkx/K60eY+Ffgj5czBFjoFXWVz/+TAEfF5YTVKw9VQJN/Rl6g+LYbTleAR5nsGPY0H
bS/tlRCGe7hSZxCCqcixjJ2cHuTZk8vcefEUW29Zx4xdbEAClp+boXjLkBtPP0WLD0Wk+GXgoMSQ
9gTlhhVp6JzNa3cZR+y2L7C0eFLWa1XpnV1jFObxAKBF2qWLCCFxlcupG6lTfhTCDNzyZYEPDaDn
Y9ZXChN5Llu3MReIvirSEImhvf2hh6UhqD1OwxL5yWeEycL5XJ6tGCs4SpGEq8kvDOWruh+nBDuI
IeSuV6LgWlmq1ofYbNcfcEIP7zIa+a0TP3HT3E96OL3QyQ1VL/kOb7d5hmWo3TRW2NdTd6e5e+uE
NhAax5lD6ok8XPFx3vPe50+7VtEv8vQVEadj+EU28zGMOWBrDnikyot39M/rqwGt+S6x5USp9/G5
458n1rBTLpb6lDCBbA880jbqzE4aeldTcaoaLosYDGxP6MoMrSNTE/Em1dwaWocZjry3KvIbWyjg
xSodF54uWt/Vkopv4qAkJ3XTs1xpGG3S3MKKJ0YtfhY1yG8dzsmuQpYUcu4e7vaIQUsN9Irf4HgB
g8nnWFrb9SXjPdCAgLBrGUP6jUfG+gqKGYkDzbxZzixgKpDhluyAoVptQZH3Pb2woKm6XxyBwyLK
W3wYqbXVak5Ow3wfoYnCYsz4HFO3wxAI/0OL7yeFLlbilf3KhiXbJU4MeFmV7hiLEnw236t8n30+
K//SDZkSDNDBck3j68viGZhQWkNE6QWP9yzv8PEeiJqce9cFyoU3VbQLV3PSPaW3izzZ38ib3o21
071SjvQiy2m2eirpznUR9mhcrGHjmLvty56d9GUIXjzzNQ9sJOntti8G4MBkyIc1Y5MaMCpz8FRy
oOl58OrWZNjzZixGThqLnxxFc+KOGLMZdzwcWXe8KOFsBJAeXBQLDhLt6Q5hYjqHx1dJzuU3e9km
SUEtx52zd3gVDWZk7+z6rEQ+4kg7029BJplblA/pbPvpOrcIFkz9ijhXzzHRtAePoaiACMeyAbUV
7skUiSh+3DZPzE9vBCgyQr5UK6+zW/nwg78uD+HiTlgObstl8mKpPrmRXl4MLgbk61sRQoaDvGw/
WpdjBncynccKFq4pt9Il2379/hEtBUJQkCoNswloVWk9i+yJ3dODqcVUMz4hUffUgZF79omy6itQ
yxMDbvCMwLc3AjFx4kprXhsao4AzIXuiv1P1SzMEkgNtJHbmWt0n78nwlLTSHoFElAP2zPs5bDWr
UNyXCaCmnybzHEtzIB07Owqutso/OiA6QZq7Aemw5/S9qx/YmIeGYdQuk5pJz5L2BPdhKc4a8lpP
T+801eQuWhNgUl1PUWfErqy7myWCCpqJ9oE2QQGuA7H8JMMyI0EjYtF2z3NXMS8X9hv8WCll1twi
itZScq0+WYGXr2Tt1ixXzjz9chl1y3gJrro3hq14czH5J0FwWtz/t+x8ve0vwdjjTfR8Tl5Ky8LJ
HuOkRVaBNNI5c9MkFZYDJT5wDLS7t6cgqCFweA6AEEKKHnDCSc5zHilVX0pMwTQAP4Kve8UKCHjQ
f5J5tOGTvWg7kAuvGmK6TVNG8x5Ifh3XZ1idp2HOkBxXLc5iUdEG6zffsMm/z7W3bsmpRN7jr1yj
dOSEsWaKxcmrDoX6wxUd7e+J3iepjBqR6YPER67VNv4ULNZZrtanwnfIuj0K17OalJuwX+p1eKTV
WR4SYMASkGcNarHDJaTypXrWDfApr1GpF/s8kIF94BKxdDqNA0E+5fpIvxvJR1PVylQbJMo5mQt9
mCwU4olTd+VVuoMzaSx6v6/zCW8fnZ3nYEuBGdaNb04UIAWHHjpDfvAMncrcKpOmsBentMYzy20n
IND6RH/JltzPXzYoFR+8sXjRoNMTmFaS47nUUStOzbnebZ9jjF6rPHFBdloEr3BnNG3VQjGqVwUH
GzyHEo+jPdefORTWRUVbhRS19twgXLkPF/FfXKlpMwpZtk+w8WLkCQombXSbsjbNEokQaoO2mN/O
CQXVBIKqeYtwE4S3d9n4lCGKN75jmWZXzhGg6SEtStuZoLi/W5nChp434F/JRITsqj03eIIz4hKX
wd6sIIt5yqNw5AuXLFqTffvUUGmhVzjc9hBWXBJ/ABrA68GCv5SYODfmm691sYNkvUJUsUASpdRQ
Wfci6Ko3IRSjdUMkLco1jN+WmNBPtW5xmKpOkaM5MlPQoOvWNgHDU24HvRSmeojKHr90Sg9Xs0HW
P8IlHxmDH55jVohumQ23I1x2Q02kq6L0R31/RRiHWWOzSx4Nsyc7xY4xl1Uv75XHBR1sLmU71iYU
bnY5GNJ9qy1ToquboDOIQ0F4I/P8W99kxIOTTwP20cOvZGGp/jHRLLn2qp7Ch1f9+FaCdfH723xt
ynJ22Kh64S0B80uk18UptxFp6BoONnM6w9Kics3ytLPZN0Hig/G8vCrWMwAR40dYnBEPBXMrzF2w
YuStKA/rjerL5t7ITWl5IFO8QD3nwyt5ET2LqgixQA1FCDCu4lYW2hkDk9jHYsvpOe9dVqjV+f38
riTtnNmNc2s0N/1WmfzVGxfDCF2q5Jd36tWfm9GSCB+G0vrYySX1+xo6YsDWB6tDtUeVKRPQbV1x
pEq0r8yjDs5vbVFw8DK5WdVBmgo/HW0s6lTSZFHGAWsvtHvBWiPI2X9XB6mPMYYzLEdbZdxgvHOr
ulbJTFJb2Ia3ev5FNENEmoHJgcqS664vFeFKFhShrSH9c/ESLDsk4jI+qX42itX7Cdj83HL2Orli
6TXfaIrWOOEkzSNoFnN8vuVsEX4mV+YCj40GOeRHnJe6pjFnh2D7e6E0XZcq8Jm3otISgS1H24pi
6H1jfQ17w/0h7+HozOpMoPxyro0iZCvPloWcLworlHqRfaEZUD6XO/oxMFmzFX2lPF0IxISTpryc
j/WlZ3TZpPxcUHG1oDNLtdwTvv6HC5aoCS/ANbVw/LmJUxf3Ax7HL2bRHGgKj3jyLzp598vCXnZW
3dJLgkjDgQ4WCzchM1cA8i0b9292YRdItR+aKthGaWu65EqMnsv5guKEdMAkz4kwYKrctC6uMb2P
Craicb5ZMcKwGcb9X3s+qVZo7u7R+mqbQc+lM5T6QmLVaQ3mKpVvg+PI9H0rHL7AQBOjDAnucDg+
lgb2nCVZlLX6NQzHYNV80JhJGL+fRx0tdsrWK6qnRsOMIg+3jKJXniWAMGKycI0Ce0Noh0rpnEbC
I7VjMorrLWJDlrTXwqgAUUHPcSA2MBTBFB16FxufwtajDYTtBKfIII57mHP2ICZ795D1Iziww4Zx
0imVlanPbp0FBhMaruMNtBR24vqlfvnsHOIkviaqv3s05WQRTcKHZbRSqgXEXhOpxLwwr4dzEUYR
sfyCs2gYseM7pU8tiY+X42vlTcF8+1G4cDykpH8dof/4Ph3xq4/YfYdphpVQgB85UsjgBrKNoEgE
8GAM8tqVsU3djjbJGktiLQeBfeRasH7UVjUfWPVO+HM6PssIqDU5On745ytHPpoptAKE2FTMIVFL
8p1df3TyThI5pg/zM71Qr5TRrgp8N6uwZa0UajY5TAjOHf9hd6Yc3p/wyG7vEtRSHuAbPj2tlM8p
3/SJO9NH5khjUQqiE9HbQ/Q6YcB4//cZKfrIJljRvHGHYZj8prrAhwuHQIPSWbMBAn/1B9coAbx5
ts3R0D7bmPis7KU1cl9TlLSEjNBcOOQaO2i3QNNrjuU+7GL0tvBoSQPZzlYqMy2R36sS+pQI4HzE
890oeZoPz49+jl9I5ezEdz81Rp9mYWJXjxWgJ4y4EZgAs+m6JhWhI8IiyVsuNiSmM61qkXKx6gKK
AVp9GKE3vIMBO/ylq+9113fqXLw1MIRBGuRbxeEPRJxgLrU71A3rD3n8lc28QH8+5DgNQtaWEFh3
64gh10H1dd0yQk0EO8zc2yuK3Guc6Et6cfpXikry96Cf0TZRqQnn0lzF/tmMWPR/gOaDy6FizLhV
5qUyoaUSlWn3uw8HJWGlTn3n7w1ZSaMq/RIaZMQ/a+w+fo0dECD3ctuxS5q+CajN+RsrMwKNBXR5
R3N2JDe+LPADMGk2ngaThyOkUSFtL//yPfx6VtWgBiejjnCqr/RA8KwG+UtxhTjtvgpmRJRfHR3N
ZUmeXZLeETaT5blTi9AzMsD4zuVD6yvBXrJnFCpnYIECDQgzMF+YBzocs47uz9SoBWjO+z0HHbD0
sqEvQV46iAF1yrBO4ISPL8RrLibkPp0GRHML8DnmIDWdqjS7J/o6LKfLWzdxy9bTZBKPeJ945i3Q
OB5ZdcjGswsNa1aWrCcDI/GsOqmjuk/J006ZUftJCkDWLGXYPHl4pme33aEAua8r4YmGdxLFE5R9
d+mWGUCA6mZGA0TtiWD7Mlgd3R6As319L7BA1gS0AVdRGZVOdFsfcIBlPRs5EGBpUztDuG9qQa3W
WWieL1z7x/GYPCOFy9lMo9L4pMg4wnifjLDiV18bchC2tWih6LpbMB4MgPXyEEy4ZUsQ6r3L9ZMj
vof7Km8quEjdsi84azaNeSmwYwqbNQWe7vAg1PYDvAOq16A4Rlgn9vYShbospBhs+v3Zy9Ou9ZMY
uEYK4FmInfwSD31iZ+8c9KyrIIpYLh8WWYArscFFxBQEhXZJuQT3SMef2rFxJqTcxNsS7Citc5B7
1kBRIhyEXtr2e4tOXHBxss1xtmpvL0vpB1azcIuIi+pcpeg0cUJMfUJ/SpufHHIDDk+h3O8Jz9Wu
VcX0GsOVjyxNisITfKMFNyL/HDdT3Rmtkhyp3mV2ZBHZUnqZDR/48RPGIV/VaOTy9NTTFzZoUtg/
Jw6k6K9ZgTvc24vE0to5v9GiltEVHKi/adw2UkHNs4ISz8yfwg0fR2wAJdmI3qyK/7QXJ2YU/Duq
PacS3zmMdcVELEWRUj3qsvDwvHWvFCQ0nDAclgC3x6riqOnA3l6V00zXAaGYqOyzvT9AoQHwjeWO
/jnuQZa/vK9kBjN88kQ1nbFpwGYOKyttK2z8j43wBaYLny2rKlZEHBKVF/qG9FVmofE1roRolQ3M
NX5B+H5JJvLsVh2oZcXfjz8pvZ0iy6EpI+pk9XmKaMESjJBC7tptlfI8Tj+Ngl+UA/OgBtLUCS+D
Mow7xB1ArdKQrFyrHs020+9UvKININ152AajBNKoMlEVvMQfYhBSIfFCbo3kttzyyuNvHbM2nsys
t5rFPRWBO2HeorHV1kiS1CgX9UZ1hPCMwzGvW/XGgan/dGPIQEv5LnAPj+1x6GVHouq7daaTjHFz
5vaGnVEXj6AdC8aZ0ZGujV+KsD3ELEGa0bvEH9IlMR+iXXNghIHsQsfEdAib1BmT7ZT90z6Ol9Cz
xoTj5Pg/oQSO8LFW9ETG0r7GwItyUPr5G+3FuG7eZEj4odWigsGmGpOyMXTES0Xx22b/tcS+S/5C
fwYCjEIetAM1Oy3PqmCAWaEje0g+EEVi17Jua+bdvzzkmv/48IlkMt8VxjX8Eog0LK0i08pHDcF0
rzTJgOaZQAHzrs2Q/h1PxQVO05BfOJkgXJip+r/1kzmncfYGGaVMgi/k3+BuyQ8arANle1McmYQI
f6/4F+cEkB/0H7d7sYsV6cHl1B7Goy3Af5fwOyD0BDKWH2sVToWSjqp7sbrAzlaGTmKssrDKDr51
v2QSW8HUZFQVPNSq78hhJ1xNlhEhgQKKvstT4Z3DkH81Gm/F4LJ/2itpM3i0QFP13oVZ8dOobT6A
6XnhuiZulF2xxTdyZEBjPtvNBIz1H1gjdQomovA9TsFkeLts05wiT+yUfzkR/D8/PIB9Pzak9Oei
1zbHqzivmA2y+aDAjsQcxsinjhz4/122tkkfP/6uNtUoUn4qm6EO8dtGXw1VU5LvH8LU37COHrlJ
MtazQ2AWApLhbgEjRCuW1dbB/e6JGcOaPvWO70KxRFElHE/QSmB6ataFbhqjSmIx3/vgv3MUt+X2
SYOXhDDq3s98RdVMLRTS+WresS4b5R+91g49lXIS+QzYjC0FtaK+hsmiGVjo+6nNSaLJwnCaiIpy
AhhfHhlRTJ1nmnc+CioU8BdfxXC2yWxm+c6htdMaIPGJ+QWOYYeKfOGruNqJ0hTAGTf25EIQGr9S
1DwV81aX9pZeEc8PvQ559MB1y1SSMrxDltz3t4cwgJviUcaHvsXvW9///faOjxZ2Hl6MXINLc2QG
2ac7xEnhhigaYXWrxu82MTaX0SF1jJ5mhzgCEIjI5ya/AETvpt7plKtoo3aqxAfAP5qkIyzQooMO
pFJc+Res3WuiIiZ+KVnw8l/YfqTF6Ou9W+9gNCfHf1hqa6ie1b3mQvLLrE0m6midCM9y4vEcWed/
r8TMTTO21+RArCNhkSOjcdIjH+JEeL6qVa06S9EMjqYQs9gbeaJBBbBXQuRJqpzEcIvnHs4NW4Vt
q6kcIEPsdSAsvper73S00sKAVzcOtUinynWX/Ur30X/VI4+7lD0TR6SF/Jq6U+HFU0rkuuPWFerb
VZllEPLULA6gbI+cPA6+ZrMXxrjZmIJC9rdF73su/wQSacYfuXgNTWM2rsbdy0nA68rGzcWQ1rG4
CsJ8HehlS9TAWS6FXH8lyLAEjwzmh1wkY4QUFU9Kzt+64CvDI7WOhHRspZVVQ+DO7bvy+N/YE5Ug
Wokv3c1cE17TmGxqL32HX96sKrd7ySbDD9dfJ+vpC5biaqqqvbN9bdhgggyTYNGYaxAEa4yh3D1w
4okg1O/pMi5YHIkcvBLty48rYuDBWhlKRNzrlNE8vMzcnQ9OL/eFHWkKzbPQtAgbMCYJu+Xl0VF0
qYExTbG0FbfCHakC7b2hDzCnR8fFNrzrrU/rYQMvNWyyBTO7/CskYvqTb4CoOyce0qcWn/85gSu1
WLjkQD6QyU9ZqGbd363lDyGTtgiAbPmmy0BtMWidvOX5MWZacAFNwLsfi/kDTP52btSvx3S5G+/d
BAv/WkOX348RGr2eAoMR+6DwrPDZMHUdqcGD/BMqCQsWwSrM+YZ1mj2UFZzDLpkV4T6LBWKRZ3gx
Cc07p9VQXYJxmtDXGRNuiomsJXF0yzzUF2de0xEmOkGqhuvh8Mo/r5J94EMdLjp9dgfSgIAwsFW4
1fedFCJ9fPAR7dCQjlCG5HuRYIqkTRRm0o1tdFaWGPMzYweAY2zsehxV+TX3bnYgRhMThnMRD24H
yZSQsbHrM3Agf3Y5DJ2OKFvdUkV3OHDo6etKM3SDV/0WgNKqrLQC8CAFlIRiNZRCFRPGpXnCTl/g
+4EiD0DJazrdNQ8V35F22Lhj9puPi3beByuwGZLkxglvfC4fsEc3QbeIYBFkosojUtkDYBAJCw5M
RPJ/NhR0EgGXbd+F/STiRsCkWJB7DO2Pz+MKhbpDouNRBG5ecFzcZrjsYf+xfvTCpIXPQe/R0QgX
OtjPrQsZ4SJkIJ/SnYeab4kzVzuAr/ur0A10bSMb+WO3xBG+7rJu5j3PIF3hii0NSYWLVUsrbHMi
xYVJw+LpeDs2omT8sL9rK0jdqHX8Y+DHWBaTlEXv9KeR1XgoIZgJSToyagvuBxiCHsMvZNQcLgXB
QY/icLNh3nJumSjz9ulzgiM+0zUmjG5KscfJE8ujrIx8P4k5V68c+ol8N+s7sgnwpqMZG4KMJ5PR
FRipYkAvT5pCOQPKjbMsYdq230ODObzuvqwsa6cLnYLjtK79lEr50S4dzNl7L4WEFx0kLWkk+JLD
X0yee+34EG6sMIU7hIbJyHzZhHdmCQQ3NFTSg4TjvK2S0a8v92V6xMpRqOCyijcve/BCFKMNYQN1
gY2n/w7dcl0jWolOLtVYSmzk8FfeIhPofSbAzFNP0JTpBlsquNLBFLwF3S19D4Y1+OnYbU0Dfg5j
U1Xsr8plrgFQlBJXkalg6PwQBg1GPcKnky+GmdkeAmBCkKa9L3LDBSdvTcP58Ko2QxGs61Nzzq9H
NsOUmHrRyT1+dbpvUpt2ZEZthmgpcjgo/HZyKy0NLoq97CGuDxf4e6hE9B8/wWa9VzSHNA2jzG6L
9L1xaMm/MaFWoqBZyqBd++KfNrAKtbBgg4zWpKGiYZXthwN+FIJmJmKbDWMmRQDarCIOGXiWxr7b
DucCCbT2XDT561a+1bOKRYyugVLo4leYDoY7vWayaLUaxwhZJnTBovGmL4YOUO86XVqoWGzX8f7y
G4z5Tnq7OpVzvpZPD94VnjQgzKxobtdbg96mcvL3PbJhLEfKdJ4Mz+c+zzMUDfi8JaaGLu2uTy4p
vgqKB9gHdD0bJeikxODqhTNL41RE24ZYrinIq2djqZ7I1sn6eyblsYRrB/T/u4kaQVL79rw1R+Lz
GWHQZKzax0y+y6lNdSi/Sl9GqrynmxNbrTUrZLUw335nua2emTh3Y8AyQm5L86JPzBuNY5bH3lmh
dZrN/yVI4lU0kbbuVjPMA9FHsj/VD+O2yayoxKZnY4mF4qHOizglAlcM6oi0BEQH1xO+3fOxZ0H4
Xb7UX+ee84Uo3PCV7uwnqn5NJfJGMq6PkGtmNwdoXez++vwsosXNsPiTK5RiyQruEwekU4QbZfX8
lyeRW+s4bhR3q4gMM6h3+09bKe/8/uFofJzYlZP21nLeTgjmjO+vMwzHNhKeQx6Yth2tKhFIKm/F
SJW5+xBBzFeUxU8/g03ViJX0oc0mXl+N01D+7w/0XTjvjKzlTqBfpoge4K9pfB4FSxPVu1XNzRjv
tP1WMf4TBaVb/nr9ty0D7uwBvvU27alds6S6HYfih3uTv/O9acDazbFsqABb6AzK+xUisGB/1u/O
klTNUlRH9N55GIOBhJWqNTIIqe66r0qL7m/lgEi9vRhumHOUUQBUuZwK0LHWSncvg54SU51XB0un
XgUhmDHOpnFW1FITKnZDSpkmffxp40XlE2ZvEPanev3ploBUxUUZGdkW7DY2HV23hd6c/PZ2Wjn7
sZyK2zliDIqw3ztfF5oAZR8fWSy1Eky26ylxSp+jmSBWLzKMYuJMQch43k7HUaCpoGW++8+OnTPU
38utislku2s9EPS4sGOvMdpGHP2zb/NX7j1M8CS92pS25+uf9D8+PZSs8+60nNgq6CnnvL9sQcOw
wBgIuTkdjCB6ckQA4z92l9iHeOJLxdAzaoGYRQaa0+lwATJhuZaziaY/+GASybg1MtTmoLxhuTM/
x5R++Nw/viP29ELGRiNAH5lAZqFab91OCNfBjNVrNmwWqMovIrsPjepPNXYhRLsEAdFMgh+H4CDK
R2GVfIizl7Fyw+hwLj9j7mInnM+Yrld5an4bFLn85JNxJy2+ooeaR4DSteaQp4Bvs5G7m1NCZw/w
hSwXU26tHPvXLjqbjqQnsTeJQA03QIs1/dU/fRYldsVQ5C6zkZJe78kGZZCJGkIDwo93imzEKspj
eTH/iC6Azn7LdntDtk8rZtV1z5vfmp4i7LDH6zRLRK6nDxp83jQDRCE3Ka6RCl5j5Tgkbf1T4wi/
F6+dtbvRKeNydfTtBflDZlXNUDEBORtjBVv78TZmtJlEv6eT3uTCMyHgq3MGuHZUMJYOMZicpJ8k
yaAYxEY+FNbGz92GvAYfjmMfo0m/IHEQVfYPIBenPyp53t/rc6yXCeQ8U/6te95LZ07qaLBd0W/i
x10+gTFNO5I8On8kh2P5Jbw8IQt/QCFZPpdus/e59wcN07piQGDVE/of+NNcWtUGegxPOG4YIVL7
DaTqActoFWyqrWBD054UZl3tliGeK7RQE4U22zlJx9YCq//DZS2cmNv/1IVJboPcGtWKsIZLSs/q
0Xhz1oKvsoSS8a0O0HL34xMDJ7q3rIgzLHwQrcTCtSbv2nIakf/046ZoZdDO5fdPFEL4XL/jJk9I
SWemuPMxLm66C8BbPphK1v0bQ6nwJkFYYr4FO2g947fGindrGvNSZrOvaGfFGXQ3Oh9gw6eWZtrP
PmNX7QqHxNXqpbmt1GJsUMNcdsBq1YASBn6WTqTxdrWvaCuX8EpxK2WvKELIEN6qYh/99rz/gIxH
UzEwc+dQKSDyU//VG4qvWU2rhJ0FoFJXGYoZ0ioeLhoVPE83BPzI4jBlknyjxQrjU4yloU8hlB4X
wHbcwIuDFCTt6M1YCSRKbgd+Ej9klZ7JaAwLbboRjLtR9wYXOTnz4mVsTTSytHKwmkvG3O+OS0ST
gaVAiuNfkj3Hv/5WJX7WJXqyDn4VCQReFzXNyMWJcXj54c5oszAm8g7msU3dSa32bdluBz0TYUsE
LG4L19tK/X1XZIEE92qmX+4MMaJztodjFzINZLMV7Pf5FORzda4sXaRTgx/OlGq0UL7O/DTIdTWt
RQP8e33KbVwvNFrbFmpbqRYY8VxEwWxblu0YC23j0UoSn9vIT69BHvHCoy6hjkbqlIcXtNoNln4z
5qSMQfyN8W2isJLB4SuBBHi9bbegXCtS0LWDSZhj396oczVEdR3qGYlpvP9l8lJje5aEqR+41vuP
9o17Gggm/5z4SwiA5NtB1svk82j5MV0mq3nVZhR0ZOIMRLO3cmGl5DEvVbiDJKdS8e4jbHHzUhVM
ovfnDO/VZQa+TmGsYwlpmptGjJcM7ZzaOUdUJ3iSjlFQfrWe9AlUA7lK4JOCcJLZBQ23Acata7h0
f56wFHC+6gdveX7ue+7kQeiHdtvrn15WemV0D2rkAKfzDrbyP/6mz2ClkRDnGhXf2gGfOdN/k4/o
JBLHdrxtVi+1uAxL0xH0h6BQ1A8Z6GeMtl3YPZTIW3ql4G6Ra77XWFwMC/+K60vO4tcOtnOwBSuy
OGptdxtqVJw4IDKCdZnBHakDTuEOJQkT+4sicKW1zQy/lzQjGQaYeTiJG4rHldOfNoEz51E3kN/d
NQk3awuVTgbvllan7YvEEYLlDnoy2RZkKjnTSyQ/Fg3e+f5RWXk56LoreO0M9FmlGi4XVUEWp+0F
Y1XkyH+QKugU0hNIXwe7UCKNRjaxySRHNQ7LJOnfL3Dgwa0b+41Ni8bSpzmb/0mRqC0LQASDxXIY
tt+SEB+hizwDOgsd8IQqqCJmF48Is4/D7RNdPFcDHVJv+Ftdf63eilAXFt/WQ0fM2altm4SxJJFl
y343b0uSzOjxM2Xcy8kES52LgcEYNK7WUaU2wlaiRomjXsj3XsMTCKY9sUgjk7/02iF4vTontRvm
2atbG+eoGASBYS3XYmZfgacq/HXhRS0Q/nxKGulxv9Zy3aQYjq7wZs/qpdLV8eT57wxJOq25xhrw
YA3My9XZ0RDX4ZOMfgety7ucE/D5TNJhNxFsDCN0UXosMvnfLWyo2AxrZcavxBiHPWYZpxJ5gq11
LzzuQUjSeODwLSbg1swcA8JndcXbM/Ga09lKCt8vrv/HO+NUBhTbnj4i96FxekqjGJNiuvlzWMH1
9DD9o8cVHmDobrRT8N9N9GZH4Vq13b+m1i2DBYR8mX345vEqbxMBCEE+5jR5BoTF62djoVlgLi4l
mV2Vq7x6zaitt9MGAMk0lQT8rH8j81ip86/SYLoh2jRVZfa3r5y60KmwbsYX8b70mkVYpx8kbcdJ
o8r440rDtiTjWTdom16ueUWiniZoG/qLa3k8Ql/KeQj/BiiZWbACk3RLYiQt7O3/rwOZp57s7QP1
jX+uOv3mEe5Ki1UCTu65xfH3bP0LVYDIZd8da3qMPQngqFS+dTUZwWuyb4lSFjm3a24Rx5gq0yRT
YZAgx/ZzFqdUypXU7iartgmYlGz+uhqWiAf8wZNXeB5xxmpzxgqGx86R1zEEO/ilFF1Bv+i+9040
vtPdghD3zLP1UiLph4/Fvaqlc8BRUmWusPqc6suLsJC/lXnGX3kGlMHdO7zxAYKbjItzY76dHxPk
aNEJD7vUbNewoiS8jO6zdSBsMtTR9mHnUHMbgQ9Hpq4yR5OC9zyV7+GKVwR9bIEpnaGn8oRP9Kqz
MHb2TBGmp1dXpaGNERNHgTU3Kn/LpABueTnYjRF492972uNGUhaG+j6AzGmYmZOtoC76I/5CWhNE
ZHEs0etq4Jgi8cUeJLxfNlJE9Elmo6wazutEdJhRt08qscOfSG7m3f/NDgQeqNzJalm2PRuCwyvH
DuZp6enKuNGIcz7OPnBZUh9gd1xaTWFt1BzUeVGMflM6qmwjHwnKrgPP/h3Udq0FrYFtXlK8kXwL
JhTPGhigIQlsYn21mHX4ZRQlkcRcuMxooQeLlNPta+Qb5NKrAH0ZnuWunRSYbSq48C5owcJXbJLN
X0PdadyaPqdECl32WiTb6lXz89pQRhS/xefssL8kDm1ei770bGFqqvspNo/Daszm1v8MTe41PvvK
SN9aLkNdjSM6i7Q13UcVgL2zJbvrCch0L/s/+c9cnn3ETwcB4o28vMWu1ax6uEuSLmRCkmjhQrbW
P5CdyixlKSF5b9gbE3lsxtSvNBqHqcWf0V3nAb1N3wJrUCMw4qc/qMm45VmqXYlNwD1ykhocDw2v
YdkHrLDBMv41EC2QuzQE+pGg8KE1O0cgWMTiDq5HhzM3IvzmjFafR1obxhEw/NFFdACvcmRVha2R
soPIBbP3hXWrzwQ5LqlKxQiEcnRSwvN3K3Yvu06pGrfIgkDtZTX/bz8w13D2IHISTApa6b3J71+0
lCEDPCfmu6Bc5y4khIFqfhLWET0NPBSqerZ2nyWHNY4XM6ZEOntzBPZ3swMPwSAbfme/evFPuv2l
xxUptAMwA9SFReJEU6wn1SGNoE23zLQZQqLNpUm9k43pnF4xV9eTVPIWTLxtudob+TpD2gbqfMjB
5yHyQov5C+wh3kFjJsgwLWip/PmUaPnNCs8UrKNPVe5U0vw4ytM+JzBgk8HvOwMx1/rdCfuzf1cD
+5zZ5gOQpqEi/rPHiwiVdWc4HTDvv8kNaou0h+h8sKnsBL8FZo2qoNNMms5v68HiUgjVe374vsIV
jAxyoAi80UrvznsF1CKJCndU/fp6HaF1Als3TACbcJ9PUWH6wzwXtITj9ghMn/BoPUXrrimscm6S
TSAz6X7x64/G7QJ3vlN5VwCaCApxkxY5BAHHiIbMb/lgoAXarHi5ueLy58Rh2uu0UMvcppYWmS5w
kZoiMd2irb+7xnUGUx9vy++Rf+y7Qqb7tEIlh5OCiKewO1yqSwZwOGpBC1EWFn0xnXDZiUY7cgxM
wQ0PqeHL+tBmH13jHqy2lyeXx7xxzcWhC+/MuKI8bCGLRjwGBB4zU7iunWd1+HVPW+XLLPKhXLez
Z0uxhFOa4CoukHpbwY7HJi1YjD0/yy350cXyKh26ozl0HYPy6gcXiJF6CD/sTndsDccY87dhBPcu
95OgjYuY3xJ8XFICHPpuLCu4Yq9s+/dBxYLZ9XqtmBw1gaMSGmpklfGiH7ihaZIAV82/rC1h0EEU
Z8Jl60EatqesgFaTe23oc4mHHdCAFEzCWKBaxX6KP86uRK7c6yuwvDqvgTzu8aLrrvlqtUucZoQI
0yy+FQEz+69K379YF6Mj4ylB8lFA13uy5e6Qr33PvwV6ABle0e6hFijpOtp8pQwSy74LT8g5x7L3
2TuvKPgnXk5fjEpg86TWLPmRiRJtSosbt0OUMfEO+Pv/x/vrujqr2L0/OCR+3KAZ3lumHGHNOwhY
5sdER5RbyEBGG9Y2958XWPfpu97NkpFHy6tsihhJGtwEMyv0Jx9FMbx2p8kNK1+mE1bCCChWWjl4
5XiL0CEFETkIYK91eeQLBhqZ03EjOdZ1nkJPRLMY8w1IbWQILkATIDR+W02lbI62fbe5Lg/uRroM
7gMrp6oy/c4aw/z1Dati0PoJR4YuzyAFwaF3mB6nHVCClgtqkHRuXG3uZ2Qz3BNWzg0duY4hqbJ2
jueS91OfQN6lhQhb8JJD1b5lSnn//NGplGrDEc2nBog/JuvUtycjqKO3HW2pHL41ixY1bmyzNKlR
IoR0b1hQ6+M+fsSlo07eKEQK6YCNXwA/d9NhyySjOsr5JkczDu9z73sS7WlujrSll924gReN+gUJ
PVwaL2weFa94FmbYOZGUS5WmAvg4Cr5D6xOv93mw0llu2EQbvIyS4EqDnePOiLzMDbei2lGARhyk
GY0acLsrYNUwlmNDVkQsfAWkAk6Rrl7Rb0GnBq46lGbLCiMVGVgBboX2bl63X4ov9O1bzAUsCvjo
Q6E9yizYH8EqahsfNcHDe3EYLQgkye3JEp8luJCUgBf8pLdOtghOH5n4AgEk5416DIH2ZHEEMGHg
Y95dL0LPUdrVtcheqbirHIPDMLCYWaC4DXxxEqHA6q2TBSbsmNoDQ+TcwwgO6I6sn53jUNTfRQDS
ogbs7tJBEvDllGkeOEEVv1O5sAu0LtZ2f8CyBWW1a/lLikKY0DA5R3+uK1dxseDr8ayrLtXQ5bky
XMPZyWXL+TDa3NS74cMvjdhVP22RCV16EiY6N1cQwy17iPy3JjlTB8cdxKghTxTR6U+OkSBCiigA
mcEPnKJkzyCyX+de+O96MP2T1GvRodFTkACSRFI7b21wM9yKoOyfh/lBqsQqnbQ8nUaVq6zUCzZY
zbRSifcZShV/YfkLur9mEzgY4L2fUYZmARbmzJeZJtM6AZvUQtGN8d8ekkMzmWOL3+TRLUfcLj5I
2j7iuwiKaaO9mFEB4Xnxp3ncq4J5KGWrzXUdytMA1Wkk20mC18qa3oBFjiHvWZME8+U+bA1R1rYY
MbAd7b4/39YUzM36eOL/BPcfDfdBi1jwSfQ5SHzWCY83Yv4ejxz4iUzdrXMW6OGA0RulcAcg8AjG
7E2ag927PniCe/tGHplBV2KIGAK2CdQjP95TMyZcOAIixmZzp/fLM9VaKH2t6hH60Y03E1qNpI0R
P5wSpBvMXVItj8FJf+lkM+8MZVWjqHlFJNu7kUMqs4tl3yUxn7c8fvWCAboGs0fdlDejWOMk5VPH
tOA8YERFU42zTBFeSa9stabSAl/S22RQp/EQ3G/Bbb1txcebWZi2LvJ2bQeIaQWzJnYFhauRMpXG
WGi/5mXdF4yISJNGEtLZCczsb3qoQL97mIc3p3NapUu18vYH53uPazhOz8mrWIzapFYfa8TALn/Q
a6oLgjTqObSm6DKQLsTeYu4IutqW9udswwsiQf4xxVRcJ9/sjk6lQpg4cT3ZQhUBvjTLXHFKdd9O
d+k2kIrAf1IzaOyG4cw7+9fu4fAc8TpQewPXibc3Q8llSuZU8yEozSVK9I9yT928WAcSKf2R9eiM
JZj1FeUosSXGcF+hl7U+qRW365h9o6Zpl24KL7TReGthqDz/vlVOKkZS6zPokBla24zNmqPUK0fk
PMQO+q8nc/VRy073HOH3fj1EbWxvmZm3fDzve/KTxqP9OSQMwMwlr0Elm7yzfpmgIOPnD5RmXM60
4fhXeWd7s14kkQqamFqO/5cjqwXBAovbo0OFyGzYltPK/4s+XHU3w2Y7jLLDuD6pM0RtBWhn8i+4
pRtBrMd15t3aAFjVYpAdpLDYiJjpmCU8B+bNklu/0toP9i7/7kSC1hwQtwg1h34GfCTuU9gG03i1
BhWVX9RWhyN9VJDguk4jmLdT4Oi4tSXS5i+BkfH4lxG3iNgE6d/WUq6jG8P2ncyMiW/t3g1fmtUu
Jz2p8AuEAPTf3tROtCFISFNEqI8qpDw5iIFubQVfkE1p7OLJ6aW4TUyiqo6uhokQ1KMP9AOFw3EE
Cs+n3pLxcTe1mOkTWwI4J/4lkugLBedgUTYQ1jSCP3Jbu604iXVMjjaZAZ+zweNutEZ+VPdjOxzX
4XfwNbQFlPRqL9D9f2jkWIQDlMQRhCJwZcSQnZmqZ9Xh+88sSDj6DfGPaUTrthHJbVDKxoY8797D
GaHh467ywNGxahiOcITDkbDTcmRwE5StEIW+929JHOnhMMJvQoixjNpUHVb7/rBb3c2dJIFZKWuB
n6WdRNyULmMc0280y2mKfUQJDMV8rrlGg+8L3jVyGxHYGcYWghPiSGNsTtm9RbNzHWH3OgZEjhlV
QfrVVXTBVTUw2HYF997BhEnBiPJu5bOoOeXM3NmDCCyWS/cwJWREwivI2Vl5gGM/gTlt6SthJUUC
qXou5nG0Z56i/e6w8jl9EsvTCrsE9tJdNk3KbBIskwcVXS0wEFvimKu4d1n8xZN38iZqEartKMt2
//nvHJ3OOoaVEy1ZhUjcZ4HUdA91XHZ6WagfgzL3QIcLVVY2NdL4It2uaBmYu3qUyBt2qf5Rkj2y
H5x9EG/YktdbsisV3rchmiWMQx3u4EeVybF77uqEJZz06ZX5te7eWQe0gaZYeDCM7r6I7ITUGnaE
kFjxSW+jgjQwfWuf70GV0/0k1jewTx1GXdpXS7AQ0Nj2cR3/h+8y5Pl4q50FimKZ88YpALBuZOTI
4XNa+8dVjK1NU+V8Fx2BUneVt369sAF2okANBhaEs9LFiUqLP2R0OgC95PzS5feXyXJzR5/vE0ar
iaMi60mKD6vDiapkQS2UsA6KCzakeUNOAiMPcZQT9VKS/DlqlemiUPiRNTTp9xfsirmDvl30Cli8
FC/gfq69Urwb+f3CYKDAgsuRpnMP2anZhT+ZRCjun905EkEzRNfhuG14e65Y/UsqkIeJeF8ee4CN
hnrpfnEWpzGDSlT5hl1e8XLINlDdES+LJrd7hPLexP61CSbEzJ63TYqPLCayRjYTuqeVu4HKwW6H
iv9r6L+2vwiteSceAxxOF/tCGaSXGrZr3CEfATx3ggLjdVsxMTpPGTSzGdz4QZUUULuQcjeWBMNN
PU3Ti3tw4P96BDOjwWHsVWcdN24qoRhHBXRMjdQKz7FvYco/cJ5CipyztUm6X4P1EF4HLydInGJ+
GZOV/7FdmZ4H9971cfwg8V38LLmVzL04BAIpCRmS/sbcrJJ97PO9ema7peR0TcEZDZzmW6HtElvh
O8GmyR3Lv/fdWm/mq5Zbzoj6pJ7b11FT2L9bw5nasW8B9c/JT6+SxrSgWskiGX6OLKsH+gk9GqrC
wotAmL/ClNumcmVevagQwxeNzb9otiZjricz3jSqCGq2SRRxwoVwa9Rx3/eJweZ1pRZ3RS1wMyoU
OPXmkkIa1r8fUzvrUF/5qf3GVoIsdqMPzvYiIIVCQuZYk3i3FjEes195omp/mgco0vrbRhUX1a/3
66fSSaTotBbfTjED8VsS4w+LDSpG9LJxsga+tKTBmqDOt6QqXARmaYwFxdD7/+6DRurjfRFNdbIJ
v93JBk7l+w70WMkVXNODWliXMhdLHzHaaZh9VGpMT61H2Isdu7Q+SBFhe4PD9v8XoY4MXlHaC0Fb
TKYZ4ktGFdtxn+q3BZS9cY90ssIAtDQFSp/c+s3GrjlDk/Ko1IbbSjuE+oWihz6peVsYu7UcMN5r
jfsNaZ2xiECQCojiEEbP5cQqUXGtxUk6OHjmww4TJzIL/gejL2nMZdjGrCXeCdqpzgK4uiGx5+cf
G7kGMS/9BiKBJQ+O2dIK+rR2iZ1b7eyR5EdHS0S4lyqp5IPMmru9jlb0rRdFhAHGHT2f3WgILlgu
XduVkKPEGJVU+thKC2VQWd/2aT5esKqzLnHPQjHp02K5PT8sOyreDzz0Gthr6cnpP0dTTt3bFRvT
TKD5iXhDj3HT12/+C96nLhS8d49Uc+qYrzA+NCKTqp/xn4yNJ1ODo9RqBse5z+JBVpJ5s2rgGYOx
P0RIk2u8fnQC3dXkVNJieGOlfbLBkHdzaRdnxy7RkdqSesr2C6VI5RCIFC533ciY5xcID48E88dY
sTojwrhlHka0xQkKyIcsr0LdqKartHk17UWCu9eexUkXV+s5Lbe6b+nRYqWSMAvwAyOX6ve6aWL4
wcYPsfI1twzIo4T0GCUWC31N8nelypiKFNNRKYk466Y09sgrop1X9oGybfP43bURE0WDoVKRfiZz
sydTuK+PTGViVlR1KhWG875WaiIPbUpRQr9tZYX4OT5iF8Etvpa6uMULJYHjhWJJPTz/iXOZFEl9
3dNTUnz/MN3D1+WH3vF9rMAu2eArc6/BxrMoLG58w+STXGdGfQt0s7yWEu/64f/oSOMvy7Fmwm0H
S2O6zLXH/0Ah9c0xFGL5x2Deag7bwsRLcAoStDOUEmY+j3glm3+s5SrGvJvO6NpYjtwOA4YfDUlP
AirFn7Fft4GV6qvpenS7gh7CFrA+34vll/jW1LdJarcQbhBoFWKRKzM7AF0p2fIFeCw0+i6kZne7
W33NuOoxW5YGxU2JFmusHh4zsr4SY+d/2lYNQWeIeFzyd1rQp/DvbHlETTzOoK9n6ksjxwqgRmJS
32rbQGNdkZA4FfUqgXgYgBd/Evps1d3jcoN4Zlp/OP9aE2EpYo//0eyCYSqLkgsVO0Fa5pHZYUaj
2z1u62c9FlE9mYBgBxUYriMAt7lo4hW/zN2lE0mmIsdNQptHg4xrXSoDSFrph0JdshLAwzFuY3mR
zzwkoOcdfbrw+Vov8n6TizU01E5OuYdoX3EMMWsmO7lMOsP1iVFZIMAsycBlQ6CqFsfNbcAo6qpz
AeKKUYI8LpmIg0WF7V1wI/JohEN/IASenGRmWNbPGLUFLMNcUbQjWyrkCmP8iaBJpKbSWl57Y4XK
FI6JWjB39t2YJd8nl3zoojlHf000TmUJ7UL0QdvZYO58PmX7hpj4sUNUZrbI+QjRU5G7nwXfVl28
jVNxmckUVFPvjZMLjmHzLsgeaYQ9PPihZ6fVcAnAUZLFi9klJLM+Pd9KRGmhn+1+67ohMLgm9Jow
8T5/ZI2pSbyyH9FF3ITMuM9OEhWxZjANSICDdGzBV1n7MKE7OrgXeqGm0PkHPw8mp72V4xg44T9m
IOrstpbTBMYJ2SqIjSFCVj3EB1V1VLagVFn0sDYx69anSawq613e3GiBSN0eyQKaBbzezCWrFytA
lO+cg3z3Jm5fd0S/5BkgN57GOEzqSn3ER3XxOz5wWgSwmsbxz4H0sfVXI8gfT0ESwDV+oVYdRfAU
Fs0MXEbiFn4bPuiVKfXLOrz5Aw8b3pgdXThDM6wgH0UsQaR2vMi4Kkq3iWqjF9ZtpJ6KvCV8k1RZ
pY4js91JFdeiXOonFEoHAiF6u0cU9pyS07tFlA4CVWcw8DecBRW9x6tXZY9+MxYLni8cqXB4o4UR
csNYIfq25Ep/DgbSs4qJWOfG8keE6Wkq2+ddv5/2f4UDtawySA/G7B1CqsN2Av+bLBh2vClEkWCx
vRwrZBosJkdHuzOX2++fBWZg1L+AWq33HmiykqGKC0iXRJmaTNICA+jfrrKz+XbjX4m1TkOINXC/
yGn4lcZXHXMHQcdW8zIYcJ4Xlwb7q2l/U3xhhY8C8IDoRTReB5mf/PDAjG9YPrMbSNYQSQZdfZAD
cxD8+y4K3/YOFA19KlxOynSIg0uEe1WyOfI4N6uHNjKCmHf/qOIjN7zJYIxy0vCnKCYwEMSNZHvv
4rmWKnjBJwWJGHqwTSMsgTI6fbyoCk2VfuVkZlGTybT9GOjq7trkCRFrv4OP4G7bio8DoT5yQcnC
vzI6Q9QBPe7KMHrLVeY5K8VmDGvQNrWUNGCmwEVP8a8pKejs6JOVAVnC3Nq4aHGphSxC4z68SMTI
VP5NG14FiOv+fSO3s4aZ/RF1LIpwhvt42yXNbLt8tb5h+T7QX397fq184n7Itu3Ugz8QpsvND9DG
JMPHdiuoMTFTpX+gzIzCxzKJYWH15u1x7/lJ1U3r1IeedpzljdxBVRWG8396Z2n0vSE7h9KquAgp
D5MC4nn/RcH30NRNjvBVcQyP4BghPGJG7gQkw84icwsxzAhjSetWQBffm3VbS6mVTD+Fx4cyLJVq
xP0CeTCe6/sPqzKAvXHV3AmNKeZn29N9Mqw62D7f73y3lyDdSoB11emfxhxWFB6IeqDKao60Pr1Q
uP8+CKPevf5t8FPqLMr8pfKawpjNBKhnkNTnyNby/1cBYVZZ55aEK4k5FlovLBw/ooUFR+W4wqgt
WP5rTTWSoU1RR4hziV4/xtl3MnFvLA31rROBNFhPoFmIj7WGQ2fpfxTePHU9icPx4WZDmxizoGHh
+4k3htfvoPnoRTOGAgTAB9MUcr+hOrCPQGXYzt+bQWMlO48XHl8aIYcWhhgAcPleZBINeOUDqV5N
Y1uHt+S7fGNUxQzGDhRufFO0a27zjNFKOanaNXXCbXzWHCbFw1gt9sAJZhXMYEWNjDPJgYX+3FPR
hcmvrySjt2Zv2AQBihndA87NwMXSU0gJj1QdXLlLvFrUONjnCPiYmAIoBn2HeaQNu7NG0rLv68B1
bt0PwRI/iG00GtV/mNd6q7d9yZkCHpQxW2yZbZuAgv3A/WF5RwaQ/fZg/FhnguWEqADj5Va3B+oQ
QnyHsFMIuBSvj3wdhdKTZjBcCw6Wwz8XlxNpnvJj+C2p+wfoUksvcu/WZHC9iqETWBp7DuBny/71
slMYjVTGJ9pznYrckaspQxZczaG4Z7GGcUh/FVCxb+xga8sHeZg+QnIZq/XhPR5yLVfbAo5QHQzX
5QM+QRs9Zf67qxyqtyyvfiGzstoMlRmg1yxX0BnYvZxptC0nr2BMa+my/cdK3hGi7GexlbIJloPk
cdJYjeD36stY5HGjc52eBs9Uforji6KFj2DOUHUjQqDxSzKsCz23dPbos964dvl0YWFtivD3HS69
mTdoBwoBL2GHsHbMnD/h/C5X0JdhTcLKZwAYZMNzEAgxImXU3PUnzPZd2INW+SoAGRgdc6aWhIqF
Qjp7YEwYtaU0c2ey4wsaVMoxY9/6umhjQCt0c3xhbEnPbYoT70x3wLS6Cg9DydFVUJceyEzsDsvO
WELlivYf/zznzRtsnzt+Unm70AdqUBVqReV3RHzbUBbhq1d9EEAZ6Rj3yW424ma//If3+fVyAck3
vSikpPFJSg95+NOOD1vg1PV6QaHB5Wpr7z4gzO5nstAR2pK+bdQdRuDDyFSnpkTpO87pL7Im79Va
cxIHpttdShr6tlirNDeyA6l1FaCC1uRpU/lUGhXyNjK1wCqzinVNv7lAcPov0a+VCga6OPV7cO2X
6F4odr7umep/KUcunlQvELy7A07OZineKOT9SC39Vx8mzpyLgmVyz+JWkQyPbsPs+Q8OrhcCSfhp
5WXD7zw2lmIj3TLMG4dJRQKITQIaTR/xIDcujJD21mjbGn5V9fkt5XIJPTYo7swIWOumjwlVt38s
HP8DVRsZpe0aG81hfVUFCt7+zDOBBXakF4Otwd372BzYABjRUjkUrqU5193uqX0Mpf1aosS05fOF
lTX/7HQzG3E8ILeL5wQ605z8diwZ9BDGU6u3QGidN5iXoGWb75LADE3TVWvfnZI4A0vbG4MTopob
Ec82uWfm6xJ2An3iCwMcjsnArZR2dnXeiIhM5omo9GSusPvDRjzSkpXFs1HnLJ0V9gkeHb+H8MNW
bCyPfB3gVh+m0Qh6ijMtxyep9AjTGoLsZf2IqkJAfMWZUjC4DHfrMOM8GxdfdBbXUEFojLAvozwT
hISZslN6VJMKtXKi/sj6i5bP0m4OAkkwPHLxz8Bjmm+MwjYUa0BC3WeRrSImuZEGWFEGbOfi959C
KL45O4H9tMJ0cexPn5aqLw8Q86v//jAc0CmSJHEtOMZuSooYE2u1vLbi6z8URIDY7Tr4hD+i9GjI
xeH66dybI8x1GzUHEuabCJhpQoD7Xpu/ZFKs+Qd75/o77Th0LBdDVZFA2YUCAThW8dzk4cXtxOwi
5Cjo2PUPoGsywPvN+InapNm03+LqJbVhfqejOO7xPT/HrXYNWz/q4mGQ5x2bdy/eF4YdtjaVIlrf
I4ArcWn1I1wexYdnGYHwJTjY16EItnUqIrD0HRRookHSUXbKA97Dibe5DuX9QZMmgCQwhjCvCi7a
okAiZe5BA52B9/1ZbEDxgyj4kIQ0JAwiJBVQMq6q+Q+HOnoDc3sR1w04qgWdFMV6tvmqTQcMQjXS
rjhG6qTgiChUgm02lVh6LIQtAdG8ZPzCy8UxhnAIEaFbPbFYuRgedC7W6iSTaiMlAdU5/lfIN2ab
CQSps8Vg2Us5BcS+2+RtP08jsd/FDxYUTrxt0YimJ/USdTRhH2hUyTf4J8ffba2DS6b+X3jroiYN
G4kWENaGEPyxofKth0FYqQ5dwy7m6EA4cCLTijJSXdfaVCNwNAlyDV6j4QZkcJkEwp88jcPelovA
NFsS0fliselmoJhIfcYhPvaWB8AxdMcOCZaidheWc5g9qyvpDQU5ZYboR84SZXe8KzZqbYGsiUi3
Bf6uOJ8QTELn6R1oa3nUFlnYAflAgPhaF1iYvUlcK7+kaDZq8yWg9hVGGCByilbOfBDeoG16y/Me
N+UUn32QXkWCNyIFQCmxPX4Dzf66dI1WLHZYJEHnKJ+tWCg4I6uWOthq8Ohw2efmOhVDk2ILFyTN
1n5YQgrHB3XmdkuzmVRXcyQUfw7smjLutynlR1a46wnWzH5/gNXTr0iFS5N6niNGshWsqlM8S9aA
IusHx1kRQYEiIYMjjCO1/M/8x6q6tXhJ86tlYdxeexnqJsMefQ4CdwtXPSAa8QKVJCTCmW1T/EWE
IQQKG39j8DY9zlTXTwzK1Xve1gLBzkbt4bfqZEIVqAz8XrLluYyEWJoz2c02QWSLqADjfMK1Fk/n
Y9nonksHoBuAVWn0P6X5H35x0eBN53e9XZBa9cbdYa29wVIUtHwR8mu22cbKsGDfeTJAvi8HQxMO
IYlBUkPk1/KLwsgpkqS7+ZS/aiI+P42eN9awnpyfBltUMUhxwcBUWp8vfSqRwdrNNurguCbq9kDQ
QeWH2E30s0TfKpx1Fs5PuS5jqsO9kaGwobw4Mb01AB09Gn/L2IqALn1mAbIQRR6nNz/yFVgE72UQ
q2NiRiyth/UfeRtCcO/KMp0KIB32wXNpnhiIzfbknBMOz4zB4LrXyP2nvwEx58Ov5uzI8BV4CjS1
fC5zkpgMxvy0T0EwhMWABY4KvvuCrLvxxBhdDTr4axyQHx1y+84MGrHpymA9i6QcfJgrj9nsKkNx
mG5ZGaVb6JnhfUE2pzR0uzl0/NHc4Y5hmDuuLPR2v0gu4r9ti/9/FPfK4lXATKxQ4RmYVEhTpKpt
O0EZai27UDwDeKRWKoxlWVqCIPVQ0y7GR61F4yBSkAAG1cVfh/o73hQ14vM+vPdFTngPWxRlFlyL
K1V/6lVVUOnXMXVoQefxk6xBeMCP5bkc919iLvapNG186IVED9o7EgRvu2LwpeM0jsGA0uOpzmpw
sp6x21akdGZx7hjbjuLAcNbDn1bl7oIiQQZma/a38F1xntezfzeJm8tfGoB09HTr3voH/hgg4il/
VT1AgZC/e19e1OHupK5tcHlO570geWhEgiVmV7EsaFXjlXwWdkw/0Tk3NFo2Qz28iJGEFTVzxRVu
d7t9KwsTa8opiTcRYWl3vgxryysGDp9GrVn+t52o48+UjQM93H2hq2xRiDewHes52yQCKaHlHCC3
nYbxTATvlBlHQ7/xCeBuAlHBe2w8BcHzzqrhyCfZk2xXGOPB7xItNdGwdFFa7ioRntfZgIsP00Vk
U9hg6h7wt6sDhKcz9H2VCTU/k/TtqqGXd1ZsDqqKgIbh/W+zgvgcFc+EQBhsWB2UmA3eLIWJTAc1
7O1bST6dvZFJ1Vcs1fkNAkwD+vZyZkw2qK7UkzqtHzqmO5s28sOUG3WmlKhms9KjQoLE1+VQecjz
6oheSZdCWOt6gCEMog20K6SY3nJJ3s7GyG1EX1sITARlovCX9v2tCEl/1l0zk6xAwVCAD0ovov5b
r5Z+GHE+8V84dTj47YOR6Tq5OoO54XtNDh5foLT89ksyTx10FYvzqvxpndvjWye/Mlu63e+d/tMO
PRwHFljVbX1BO9+Fuu37fqwXFmdAJXta87iX8LSO++rXpH62jXuICT/GAaArxhsj2Dnk9SzgzX8a
BHu7+w7W9phN7uj4XFwsrpnc9rpLK+Y8fsURPej5XIiGBeX6WB3osX9K3acuoaWH3u75rBkQZvBM
G4geqGHwsxjawGhpxqHjgVE88lUgc450rzL8dX/ZLUwTOWGqZV024RJs3tyg4ye1MTJkKKb8f2qF
nl9WQE6Uhrdrjzzm2nbr0oWk8anKC72zN8CdOaX5q4KLcT7gWvk+uo8tRJFGHk44XjVCe6nk5AyL
OuhQHrAkURUmKtuvRXDZ4zk+gZvCX87B6sRuG8BkpXNNkueCCzJpvxmQUj2so3VfPCCNlJSh7ZiK
Gb7bR3VWoDyS9IXNIz4OHTK+iiSmeLKN88pPtn65OCu4habMfQOMMgow+M3C9p+GLwq22xpV7kwx
0AKUC39VgEFqwdyOFfiI+JRyBmJ1vW8lCSmyjn238RaKRb0hNtlcanW9znlILd8Ln84lkpCT94OS
3r+xPKRHdTO0KVvTe71yDO9GqdSCF1rM6DmR9GhkJGDdaTOom8BikmBDKZneWaYuFdbTHV5N8p65
hJr9UJeQr9cnsMZnPan6hIVOysHprgFzhaIY5xAIX/WZ/V4bPLL4EXB85GX2xqxKpsuqgazmYhCE
jnxxupNm9EkYE7o/cWcIw4e3dHxksV2AnbwXECogZvOY+yKYhHCuNlBBUs+RmOWKH4OOj/EOojgs
E53LxtHz4PAAwvh0beulGzvOL7MxoFGkpxyrFptXTLD9ZUmNmW6VD3EUeWT9y2HD3x6OtpL5Y7kA
1dhrb18mqBubNGvQoiQwmtmoaw5SLofJTg1/iLq7jQ40vXkr4OVJNsQKOnKuA1ZxZEn+v93BvWCh
Zs8fCL/ZztzsKC2ErkDR2hpFA4p6MP4Xh4GPTCqlJw1bV3mvd3swZxsO1NTX2VPR2Kd/JlXZZ5bp
ro4vm4UX51dmFXlUF+xqwnFr1u1XmkM6Id+fQkbcIT8zbYYLXs/bJULZOOx+n/agpKQ/QyeTRyvq
7jnkZcF43zRn7v9w/2Pz9HiawJtOysWJFu9DEx8O1bcv4lzG4IgPGq8vKKTgJgzzJlcBv+hR2don
QhSq+rw9HcJnijTwIa62Y//7uY62w4UCkQoCB6df0DWjjRwMZGRGWLa2oi3BpRk7SNTxL19rCJfE
F8dVJmFw/iJSCvgfofXaTE0l3/i/P72dLjRLugnxF7tVQBMZwfJghmR0skXZ5xjImMZFEeTC9u2K
qEkf8qfyjAmv+t0sIKe2p/dF1T4HSRK/k29AuHWxnBybFqUE2bWkeAXvb2I1RJzTHQasKUfCOcFp
XpmbxqvnvR8uC8wQA5I25TgGrzLCXhsmOn21oaKfdAz3OMmCpF/KECDHAY2DEjPmRQCw6qgdCRYw
PcAMgT+yA2AsBQO6IS0BroxAq3mBd1l7KNoXH0KymRjcQHb2fgxmel0g67Wq79TzyDu38aVInK+X
EriLPvB+ioomFoXvtacPhC2a9umbPO7DzniOm+g5mpoAfRoy1iOO95mMWmlY41xZFi5vbaRh1tT1
HJmFllbsuCCm6obinyfBL97uF0IsukoUtdYtS2GTTGnrr9Q+9wZT8x/1LjqSxhX9ei240/HYUXtD
Qn2y0jZ3vC7WlLve7fa+QhCt1BJfe6aF2lqGqlzjNIPlFot+Zi3O0PWuYX38aj6YY0OBRAVPYRbG
kQkUf0Hv4+XjkmM88SfaPdGqMeDs+pAV9uwss2AzQ/ew7OIh0aLiy51yoxxinUFkBo7e6TVZnrMO
L5QiMbsA1wo/9P3fJcRTG09LVmeBw8s0lmkKNsAhq77eNS3dmjuUJVHXLrQdVAOkH5Ham81VGksZ
1rx3+XOyrZ00z2SEfGBs5EYoAxeaLNOFf8uA8YC9OUxDc0JUrNE/71oMZj3WboBmDXP6VfJq/i9B
Pj7eY0FKw//44SGUUjF4eGzEdK2Dy2WyM0L6JRds10mj/W1iw2Cmwowz/BVA52Wp9CIkaXCNxAc7
EB5tAieeGR3NPyXD3x77LZuRV3pI3jErGmuWtOOVM2DHV3e6hFjOqeqzL2HX9O39H16QxkIsZMg+
DblKOtMjlDWlq7w3mxIrM8w3nCxrUwuvZ53h48Urun5D1N5qF+IhoBfrHODUyiXt3Bsb/vOXAN/j
QiM1zv4vi62QSf+bG3NXi6NuTWHqfWLdAXgWBYzY83Jp3EPk6CS/GXtC4GoyYR8icJ0q5MYsI4cE
kHK2XskNLCq8NzD3HQ4SX0RveeSeWHLxwUQ/oxCtvvRNJY3hW4BcvfeKJuWKIh+lFcIWF2Q9San2
BDn5qMwLG17mGs77ZsK1CSPLfXU5CSdWLsxYUgEGr5DFZTxaTxEHYegivf9YAPtPzWm5CyhHlgWM
pGj/n2FxX9MrgWTE3ykuqDyxj/GHeFeJkYAAB5q671+94aXICJXKwpRlagGB4ok2jdKlVDva9dz7
YkWyeu0KZ741CgVX/DRbxHbiIBuCCEZ5957qQ349jhVKvX/jwk+BZEEO1KVijm42ua7h/DgE0Krt
vBYgVMGRdivK5v43uOWwNeaIUEWTvJdeSbyCuL4BpB/PRXJJ+f+QlU2BAgqlyCisG/b35QGIBjEZ
dCjT2sKpoq9ZyPZKMWZ4rey4iG8c0clpggIRFAs809UofzVuxsI+EZKlqY2LTeDG+XM2WCEYsQYD
Rk66drJQM8N1i3DrxTfSd2pmTv5NhG4v5cVPdfL6N8Dp105Q0UkPOh4jTPjqpXf7pQgqSBbW2r3+
vVv9ZJj4qjJkmhUz4tbGhBjc/kDAtMBecp38kD6B8tDdJ1NBZbHUElRiw12Jt8NoQDGZxYRCZ3+O
EmgeHzLsVU0DaisnbeU3ZUvylkgsbGXIjPNXNvRTCS1YYQk/8iHOThauOUH/pL16SXzi6advlFYa
qaG1NrqqZcC8SZGo68APiNk+Dmm2et6bvPcaFDJmRprhDkXo0jAAhD2SPyUSaB7VCUgclDxgdCI7
NctPRZ4oMTjGlxYT3bxLXxXmthzB6nxZE58p3IK/XzM50edqX0JknwJAZ7I2S8R48FE45gCM6+gL
PSGKVh6SlRvaPqT+piLcvv2+xt+A2nl6XvSc7HeFIEpu9EJITgTUVwldKz1Y6DHeG1m3z42SnGZT
nDWo5p43EiUbSx7SqJulTobcbZzTAR0AFaioBnsj+gc4eCwjpKgp/LHzuxHZ2OryxjyytcOC9b7J
kNcjBZBtikY9vPsA1YgxvRHhVg+rFUVgfB237Xcxa/YLsru3YVhLWNdywoOGm/bF/5ftes/8qamz
XpbIJBUqjBCGEAGhgYwbX7RtOQSvFo63pscKbr5cnrP3BVnwlcyffSIzAAAOabAoWrwgTMwHmjHu
ZUjf0pAJivzvm2bkjh1q9gZ7rx4QYajrYAx0r758h+qJEgW9vo7a0VuYSQp5FJ/zfAAM41Wf0bMH
dUTRAKsUOcR0UHrEkXf04oGFxHN90xusrO1I+x5UPphPkcuMJrFz5fug637lLdkAnlCIdStA+6Az
1K7J1Sjm1GmQ54JnXAHxhlZhMjqsaK3bkG/cq0YG9jeylvGo1i/JZH5+GXK3dVcm+osv6zVqfZGz
Pn3K1fGo+10owuLhImaQqNe28CiheBo3tLb8eLSfq2goclnmKQyptYdXWsgQRjhNZNxjwl1k0wl9
bKfdISos3z4xk/FV/azv+2XlqC2vpAaftltO8gyTboVZWhKNvmfEYvxqk3RnglfrN0gVSnYFxLeN
S5DWpltqt4w1babJGWao8wOux8EuWmpHAncR+zT8sPdEtmSQWAJ4fbaq89MO2/JKhIIqLytwk+O0
wJ5kHYmLqt2LlXdXDk0mBDsTDyRfWUEDXgBL0eX6n9FZcR7hLECn8/ase4AFf9mUUZoeFHDDwwm7
BCRBJwBPnl6uc2fv4RwP4AX5mp+rpXP/qxj1ngN9Mm3g2i5LGyQ7erk7M1iZYt/fhtg6L5j12s+2
tZn38RSvH8/ksfjLc7qXIqh1QReUvOMh+1uGWcIq2iu1OWAOqTxgWsCxel/alcVK7tZ8Kl6QP/mC
vCxHqjOI77YVigCAPPzxj1ElHjaiG6ofvN0CwEVR64uo6KEPiX3yeQ37J9KCJfswtZ/Wugaj1iq0
DnPTGGnbVmG8xyIs0QtMOOJttOqJNtPlcaclEzG8PIrDqUCxV2pijSEx/d3jkNSQwzkbKLJaIYSX
lKAacLd6Us9QQd9NwPOYtDEbI8DNKDR/DYUNq+NSeoL1KliMmWHcOa5EVbrDs7RBgu8CqIFi9joq
Vq3p494mnfr+wPyOg1yiyFFcR2jDOZeTwbDe+Wmdto+eTeLfOaqmHfcwdc1dK/UliTs7shHzBAc9
GL6hYJq6XzmTaIzuAFlsh9fWRSYvs6X0bMnqwEkL3TRVHV6Lc47cKFBpvKHauRF9XEwN63LwpseN
uiqjLT0ZkjCz2FOJzMQ2rvW0ikwes+xYIdjXU21Z049L7KfQRBTSl2QnlO4NBs5AC+TRVACAbRsN
nEOWp0P96ZTbsJopGJ2lbjTjAYF0R2NSVmEioYPwMZoFcdm9KrpjT6noRebunEMd8aMntpK/6zkv
jKwLJve4DLB9M18ayfu5Ug30kxGeJunsQu5f9c6QBh1YzhcAcc394TI0MWyF/b2HYCjixCoyFnhN
l8uX8N+0y520+8bB7D33d4WF58lRmrxy/iS73mXlgnONc/M9R7uGEyQgPkTOdJCK3qBIyCYPKrbY
HPaPd6YPhhGXKBmFA6CtSaqxXLUTZMeCAB/rOhtdROnijmQleUXdHIHQzMxGTrgB5oMiOmSsR0QL
JvAOUgIi9snaRRAMujxRrWvvDjgObzrd09hXborC+xSd0yslZLndCCUA5b5O3NFaO3mMWekfmdaX
tiki1en+lC/LjiwfndDAI5F/3xcLYFDO7GkLkHtZbWp1QkVqfn08lo/zVeN69kr7WAowmfCYTrur
BINr1m85kaQrtA4LacsUWPqEpk9iyGBVD+k5qV3VykhJFzvo+9XMT9XCxfaNwupnJ+OrisQu6KXh
26LIkhEhsXDNXhXequJR2tFqYXWMgpSEYt8fZBxRIjjOCJrUYMXbZS4J4vMabdvaX3ZFueL/Xf18
vhY6cYMKlnoRFSyajC9HnzkR3u9ejePqMIs1DX1lleMq+gd5xi99rIbf1YTIx31MQp3gPWy61RqD
blmzKNK0ADXKliz6LlobVRVujubjr44+jkqlx07Px+EPzGcvNxnl4Y7Gj7jzmoniTG+uh7ZsFkuJ
heZbJUlzY4+RNVps12GVTXjpfor3x1VjJapLip//6WU4IrIJHch75KfGUUSUwBYo1rOT199xl/Yn
yse3roICzN24F2fFBDU6CFjGs29K176u91glf20rNyZhVaH9MU79ozjsYNZcpmdnwl7TL8sDvJSf
mvIHuJ2a0jizScIBUckN6d/zQrNLSMPChktYnUVR/3niF+NmngewQg1YBnZ6e78STdZVnxGQ6Cco
5XzTUh20Ztdr3C+Z59eYynobINrNWQpnaYQQuK9uBwa5kf/u09HsofoGiWt2FQXLv3AP14P2PzII
rWLolO42W/8kOAOB/bmhIWurdfLyi3FJjQ3WV+h+iYgaJA1olgwmbo4LW/oBAjWmlcwXvY6Akv9l
5m/mVq2NtC1GFcWsq5AQtaKyZyUz0SmQl/a1KUVNHLOrc5QsLnJ4t4qKXWWxeDuqmd1gl8H+oV9l
npH/zAtq1sIwQDU3PDQso7KCdfKCJP3zUj5Nd/dmqvmCpQ4fzF2CGG9pLmG5L0wd4S/svHxQQXn+
GzWdHK67sCLQQUNRY6heyzCFOV6lEVgfvqzKS3c2U6CIhmx0L1JLGJHRr3ImWC0YU1/8DDwY33rb
AX6MfV22e3vYrgEQz7Kv52S5Gef32LNuqD/PP9pblVz5lK9ftUCLvikK724Mx/kE3FW5jUHkY9Vs
A/kZ3klqRfSOxCg8qfrPC/UTPzCy9FGZ7orpCgQPZ63ZlIy3XCZ30U1leL5fAtgMOcOxn8tL/rbF
klTox0tsxongbjJyiRl3ndfqNd7MHs7O9vm5iEJvq7sGCpZC3eXzrnUFcqzUoT87KHD7utyd24pE
Yd6vHD9maSDICRCfJe3AKCiw0GL/1m7AHowIPh5ajTSI0RRNMZW0m/0DMz54BVYyolqCWaoJrO8V
A2BBMbNXMvhZ4F88NhDmoxCbIYXX5JPku6Gph7y7GNr/RZod6Hilb8OcdZ/ffmMb6/JgO0z8b1CZ
3IZABi5ISzSSOFIMbqks9Pj0ikuay2o2NEgHtdh71ousiZcJxndeD18Jce+bhH4G1iUtmWGrm6Th
r5aL86FMWqHXXpdqDcwNOHyhkWAwiU7SwCpFNFrvFPPhv69hYX0+CamhKrVAXnqwN6Nm3eX6T3Pl
L4uRmMUiZBXT+ijRQc1+frmsB25DKF84d6HRq5lDnO/4uFPF34Ughmp9y3t9p31KEXKDEKewGaDX
Tx+EhABqbKf/9y2czzkUqBtKgpkCgJkHTlaCc2oe0ZfTgF2t0UpAS2uZBRF2UdvEO4g8t1xTHCvM
MJmK7shBUSCIYgZaAYXUis+FSB1CbBpBFQw6BRjRzNFXEaAzjecrQgUAOAO3whErwLAGB9epGOHm
mzIfHE/nm3mFbXvTuvnRZFOU4rxOmERrQWriHLe/WcXhjwyAVkyszOii4s4KY1cQPbK9jlCivOLX
jUN8TJgAiPgirOWNYbrox9bidu39Hvsy/SdhzRlZTitdLSiufWtGOTIDaGA/5bMV51rHGF2CLj/H
qV5jHKGDKKA38yExA7gtXB+tBYkMGFu4G4ZDN0014XxKQAzSIaVFNTkIbpIsFzZRsjbuWtbcIiIi
eqMfqnM02YXPWMlrGgswyEFtyTQaNlrzKH9MmMFSb6HOHTy6o3xe2V2bPE0KUIvmPECwosDWYFwM
uIKAAkZd8AlZgC9wTKVYoWQoeeF/h5mvkPtovFe5wxOFnqXPZsCNREAGEsRjqRpOBfxIFVZuottZ
s13iDzFRR5UUWUbqNnywPpYmye7FHpfR+pyqNOd98fymlH6EAIdWC9Cki+cZw0nR7dJ8jhQBDVew
h8sGucEEZFDcdtQXkMsNU2sXIrvklWbCV+bFupipTiOSHCtEmbuympr1AhnkGajWDsAv+5ylwXGl
kdXc7OZvsQn0tt8V+Qni4Q7gaLd+bHQv0Y0gNQhV1ojPMV4Qpjs5fyQZHR5hgvrB4lftnlLHQ5nq
0n53u/kjyMhSh421oy0A8p9LGFVotDiFGEDdJMA8jIT6ZRspLzJEEpI95PtMi+adZjU3qp1nVLqX
1a18mH+HHcwI5b04WYMzYBamhgVM5C74E8a6ccjQXBdaqvMaIC1Ubs7hQU2qicZ+uGRgzRPq48qK
Y4JliK58Jebh5RKCgDS4n3PYM75a+468IgAID6WRSIq6W7zLk+dvG0zud0KNQaJfgZtNbn/KxBHo
Mf+zkvhFZ7WRhLAkOr30vMElTETXKwX3uybfhAaNgr0mXI64fG3+RURnKNHEyPcJukgLz+3q4Eqv
82jMbe6QZo9XRDUZxHz8QoQj4xwbmfHpxhqTbYqh53BlHHuxQSB1pVRnfxcNIe/c62GU89+1PFMK
qSjLtgg/hE+Xa1xtpeqIkwPJoYf8k/BgZULDKg12goastfiS0WqmgvMSH0xcPJRa72LeOzNKA9Fo
8jJ3/GQcMOr4aeoavNiCr1H6+dynS9XctZTgLYb/WwAwoU/2G0e5mBI05qcpixPni6jKKL1TZRLG
UlXzdcMUP/6DbCwLO0nVf4rn+8wuzCXdZ0xOtPxCinP/NZRmhMf6eWHcw7xTqHKmne2xi9LeNs1+
SMw5cqK6v8BQ2e1PF/g/4n8izXDBMURvxver/t7g3MCz4YhrMLgBrcDk4yRAG2oP18/EFHKAuAHg
FQkJppx+f0xeGXNveQy0AEbmh3l7NvAtfIlTvyJWmsjQg0pdy/UiRl4Zp44DyW1KkTMz4fgLhpqB
Sq4PdAqJO1DGAuN0QCr7MrD8afeEUQ8HldlfBYP5kUAYOXs0wszay9sv3qQf6zcntNL4U0Rp63r0
OVOJ5mo8cI8BW9ttZqRDMzxTmM4jP7NOBaJlxI9dmoyAsScuLXzNTTnoc9pmJh/CgldJhCT41edb
jAobkNtCcvx0QNp9C/zmgjEy67wq4g9CqjNeWzVt1nrZy4lBgSKnqZlXduFjpZ5ChqUtiusknkM3
KxN3vnBeFfyX0nO5y1zR6yZZNKW7CYylU0Z8qbYw4NW9OzIK8xw6ydu+g4K2e2n2cLRIdxT9ny2z
9xVAvbBHk2OeURRoY0xrEg0h0mhoEIBm3h+YBnaTbCwPevFFinlF0SiQ/53BupCbW1kakN4PDl3W
BmPGwceHHqKO+xsC+mFj+T3qUIdCDSRKQEN6EMx7pVLwfXOORsS+0QADjhh2kCvGau63xkuR4c4J
cnJubaegAiuTQmUlQO4jnMAhnOa7/j4rxzd7pXjF+L75NA/h5oHR91f4dhRNpoP86YjsfUsaguh/
7spCCGRBoyNZDr9uBc7Ey+Ac21AcQtcSfZD9Pf6ZzzDshFtdnTG4l3ZPSXT9ACfLhei7sOEnhTBL
2S98gGPRkoM/UOk1XMiG3bWvgir+6mlqYaXxBSerwABnftWpzAPEZKGSljNX1WoxpeSd+xRRCXKO
uElaMMi0OftRDILbot2q7BOCGsBeuKFVx9zxVqmWqq5GPIDRsfDwYkHkvNU+mAWx+F68zixhM4f3
iO9atn4H/cefMkLHC3RWwhVFMZMdeRI7acAv4atwfbKTBVgjmBiC/ENaAJHGAYBARJF4xCyNRhyG
l6TwZS142QDqbOhsawgeQkRjHw3KvUcEJjS7x9c9kLUfgM91ePqQnfSyxd8U+nHmSXlTi8o2lqeI
oVqnX9l9Mm+qIpsMQ/fipQqKd3DJXqc/845j/RE1jP88otsMCOfGWhaLUqXQCsTuRDgGgGIADJnj
WYXnCyuOERgAjp2B4np/XeEiW+knk7yz9IyYlh4otpNfjO0YyCymA766rDH/8oDYLVo3gZDDphMb
IffrFzengy182+PaCCqmuprymZxr/MK9FwrJk748GtZxXe+vLJ7utDw4r4ao+YzX2SWwt8r+JJJh
+yEavLlIkrENAxsIYrq5chMxGtYDn22vnana6XJXq1aFT64KXNHkw1yo/zp8dx2+uH+TET/mIgqC
qZTesGxXUEMKZSKHpStkGJFcBZPEUTLa7fUyN1NWlk9KQgkoXvVwCLJFmt9tmz/ODPOhqYhSUS1c
xJAd8MNplVHhh5vIrM8+U4z0tiy2FploMbopaoLu5tpgIHUvC5AWbhlseUotNQPCbJFfnUYZAsMI
6dgjXsS/MT+T135on0W4OuXoH7npomPvd3yp0H8mRY3Qc2mruanqIE6UYuFvTygzXh2F5HgbXWHO
3+INQXE54TEf9BJ98cNAdviHxAUaF/XcyWrgMKy2dgqGNNElb6ljqGnHGRRUeAd3ukwhT64j0lZV
+KIa8694E5ht7A0lFjotLtYghcaJJv3/VAd5QfTkqLvapw9oE4i1RsPkiZYH6rvOtql/h8/ggzRK
2HmdKQV0oIjIzo/MQrqqG4rUvGS/95sg5cp7iLYDHbmP+nRQ27FWcJkUJc4zMMB/YvlSPo0Eu3hH
Ag8d+qm2I+syK/tFkThEyowi1gFDxmNmrLDuLdXezHE4bBpo4fDTUDKa+ORR80373MC6b39/8tQo
K1t4Xlp1zvt9GqiVBeZ5MDLpye7eH7lyAKYdJuo+ZlH8tnN7KzkGVGe8K5FQs8IvFYfG6I+kQpdw
BNC78oNUr7a9Y5jLzuDJQdmCXsVaoakCWj4NheDlN5J/hE0RDNbsP5EzrEhz/wGq/rzjk5ttoTVU
+9C83syk+3E83gd5oBDDWWVVjlfLkKBkF6wFPooS8tL4H4N1ve4jfAKzRLa4hMDhW078LorPDqLN
SFyoLX/V+RfEuPOh7sKB/Dc3WeJY8DP2W55iMxguZ/9gzVdiKiNxQspPrg3P+8DyAb+hQedTPTW8
rUeYxxa5U3dlrOcOLBXnzUnMywjqdHbL/G+M+JuY9bAgUgOgAjv6tEpTGDsvyDvxb3vDXnWEjF9w
TQx8o9BJeNe1CCJVP7LTn5NmHpq3RBniX7JedLR2d/Yjzz8bMcY7ifMa25hU1agkyOZUW/CaXbax
Bft/PWZxNECRoEe2dVhY/FzqagdXfk7oxNhvDkvVKqVaE4kkg8G6s777tJ2LYdhC9iXJNt+dT5BC
EopzyP8v/WSMJhm78sua8zASlPy1L4Sq8c+k/ywUJ8E6ZIS9SC2eGHedtdm9fLD7v+Cq5SY2YHqE
okgKGMV7UhScv561Pe6kXz7cDtWX+630L969bXtsfvzW0sFrXrqWvC6tOBa0O26SopT2/frV0ges
Rvsitkud9sGX69+ybJuj7zlZ/RhtfCb4lzysrdzjppPVmOXUsC+DL30vqMIy9P8p9u3GMUtd9wCU
yxE7PDecdpV5iITo2WOzruCCczrrkziu4qU8lhJ4m4N/3bZIiaZ0b7O15Ch6Yg67PXz1E2E0F+yQ
cBQprF+RuUTHCa0mWRu3CpVtcr+sHoRqyY/zIV/9EWOTm2Sbx58KF0kEXw8gwqkdTqQa9HERTggB
lYuVjuX4iHzrDRW4uuv7j6+5DnioWeURsZgyqMk6Wz9B6zA6WJfsRG0sZiql9KJkYkQG3OQSgmcV
w7trT5nY4Sgiq65zYfWHHBvT0dt4xdKaZ/+M+vUPDlHwJAMUZUitlP3m91pWz+NAWOe860tghbsB
n++nH9Fpo3mwCumNgIjl612cfCTlH6Umj1+ji04tIolsWxqNJniqJFtjrujYsymd09YFbXu2qR3y
YylFJNnsslCUHRSOyPqfOhqoHMQwSACFdN8CjUEEu/yMdaNCcLXEPKKuFmew1MAER9Mt/m8hfbSz
PIIoWhd9DzYJUmwwE9mXUUUppBSYyMZDt0apK3xOySD6C7iB85hZ0gnlQQUODMz55SEY3fTgXZrw
x326DVI2FLX5iKgP3ZeqbqiYBv2i5ly7X7fIxp2ARXEg4Flu7YxWXuJMeyRhPRmXrSCcR0T4sEKg
Fv2MhHTaCJ29Wip5+Xsw7JbBgh/Str8JQyDAj7bk0h+iUD2xoVaPHpg4t6uoVgQWVroPV+lFdgNr
wgaRQ/9vMKN/0Ml6cOXbE16zBGCTxLtnbBobrQrSFiiNMOIxy9Gc/M49Cc850tt1tF4V7VN8pOou
ywzIxO7e/311QaWM4t6Km8VkQRWnWIVKGQWlCeAMxjBlvORJoFiU9l6MJLygmj8okRPuXDsonTon
NeURnnoZrmUfV8BWTMSbv89SMLRnr9oqV2a8VqxQVphQlI4u/brY5xpsWK9Uge/iT6/QmOPdPjVR
rH9yAGN52KE8Ow3KnKXuze65u0P8deQq/MvLeAUmNYQfeDOK7btBr66dJWbI/I5N369byoYZUByh
Ozizp0GTngd97KgpSsnIZ1vQ3wNO76bVVCRRA/vHmg/XSVotGx6CvmiHFySdoE77I49Ew3s8t172
GnQNqH5ZFdYR3NwiO7q4mN9UkTlpbngAS2wetz09XRls6GlhiYQH45qLgS+zGpvgIpnk4zc9Ad1T
EyWIctbqJPXOztC9hQ+ilo/1I+HrI6Z0cyck0hdV1Sc1cCYuBlm1jFjcrppmJFyNd+6fPcbJ3NIM
tbG4AFepGtPkAa8gDgob76v0d22djLTky6xC4WpBlSmA93zkHDIUQZFzKCPeLxnd9zgUazPHrAKR
izps5UZox4c5D+ood6g/1rtIvzyj48gKHn7qDT4C1UaNqQTSv3ivHPSPoyVmUigHzFCwvePhO5Yy
Tk/29LUkNc71FCqChbxxrsVCQWx8e8Ztc9uZ8fhINhRr9eSIS6eXv+/u22SfKyDwOy4tjDMvApic
HZvk00AHyxtSgI6yUNeQrm+HF1/NAL0HNxZe2j1Lam5rvK7KJQBkv7UfHt1o/DZBBe2yRxff00DB
ryFwkTmcsQehHSnuaMH/lpGZ9rwrAmfgQMXwT9zaRgwOhLlJhn9XLRIIgORIhzrAx2tuTsysHNwm
V/JGSDNDZ/Cg7mfvxqeb/Rg+NvnIZs0/cmrJnUzAyQaElDTKrqEoiYSDln8UrDKGihwWE5zrHomy
joMYdYoPu9mRNAR2Er263zXi4PrwwEmxHCCmMJTBAQ0kQkAs7xoeKrUHDIJHQuPrCThkJM+ddna2
wvIfkrc0ti+gg7dM5AXPWwLC+aevCCmt+no4ldHXJDvaYALcInK3Igi6qs0VMeZ+OFxlKGV71yYc
rssK6z7CceAKBZIGZC/Ogl+YZMLnxQCkBFHRDiQXdlE/DdwC90/jdQQ69hw6v8hRR+o93utv/3Ra
xHo7vlCwRpt176iDTi/w78iS4x8dhksNY1GbU44+iCihptH7cg4d6qSq4oEPuvvdngjrkaHPq9Hw
Zzk1p4cQ6ghJHD7OsHjGNIveXB9qMB47ZKYnnJ0zZU0WgO5wt0ew5Ll1pNeZQnxa2+uFwrmQ7Ssw
JlTGAz4DUVI5Q5gFg85XlBeN3/JlwlbklZKgvsjj/fuCS9XCbaODZW+Y6X1DnUAHZ21NEeGSKrlI
dwXXMremqKquFFctfmYNADNcCVm9kJLMhg3WAiCKZrNbHGewYRpzpX2H8ySXw8PUJve9D2ra5zem
pwnGKC76SRkRdPGp+kUfixAayB2NcAOn4cJjefaec81lvffXqFSnXM2Bcco3gjZJE/Jel4K5QI2k
RZ+y9eLHesxj4nY4Vt7BW8UgInFP2P0hvt4uzJoA/H2fb6Xoyht9+RXWqsLj2Anq0+K0Fhna+ArI
qPdohjH+5XNR2NUdRVcI1zj5QrMru8D6p/rcoWC1qyNJpFS+lOR3DlKzFAGis0SYIZajLNBnp2XU
chhiC4LyvK2plyEnZW7VRk2+ZY5K9WTviy6Q+0GTLZ3e/6czo+PdlGpaUbAWwJdVjHFKnjCOc/Wg
ZRylHc0mP1p3TChNXZz2p9540ChqDg2d3xb/c4pynJj7imHTqRl++0WAS6+vEHZqBDv2bIdXbiS7
bSYtiYhpx90vFptqgLxXIERmJau+so6JwrRLXxnZNo5ypxwiXZjeDzpEn/3dCzAlDODexHHn5img
m0LOYY12K5NaXkl2A/PIOJ/GA18VR7Fg28zx1weUJBOM8t6kFqN3luizru18FavJZQqqrnPNMLez
dE0Y8AtRKZTmaj44qacA34Z6aD2RLtfwunByD9xLHe30DoKYNEB81lB0zKR4bY+wo5imSY90KYQE
trs39NkkaCVpSFvStRCt9JIBu3UoQQ5fSX2uyMPk4mWn9kWMz1qnFaWAznZLdVTHJiBUeWWZVtSD
4Hh0EpG265vmumphBstbwUgHm3qIg2/OKhQwiP3Lf/hJhjdRpeAIo+FGxpVDeLlsddEQqz2b/eY4
bUpfgjOvMUMiPGzswuHK/Fvy+XfNwuuRfFMZm+07i1kk2Mee5ldF3752gT7dk8W4E4dk4gsRxHfZ
ElvQPwvQfLpOQaO5EDOYowZkj/Xb7fT1nPWgxI4ZD+qIHGHNB6SQv4Bxz4Da6I2YpUYk1GHNNhCN
t40xGdurfyOWaEBpTn3m5spO6OE+EHl29BQEz8OW3lGjFGOJJO7rlKCzDD/q5hmTbyzqkSrMEyqd
PNbYSjXAd5nH5mHrcLm1Sf89sSg+6VGkiLoL+JYZysl6Xic2JkMpAVp+e8vdOKN1FqFCrP0k6zTy
MPWl0vAN+UDzYQ9XCt5RcAljuHmJPt6P1v2FSLFWhUKxygNGuip8DJo602lrGWuIKZNYQnHPCVdU
GEfL4cu/7D91UZuuBJNlKFrKLdGKssEl9eZuXub3+K/VD7lijEEoyEoHTjEzLIBuSOzUmpi1t6hA
+9wRcoeHhvQcyFZ6ow/zS3HVMhqg9iDXpjysIqmfaY8QjF/yWaIu2wIiYJw5N0me1Ef5h8Az1IIX
j36Na0bdl33NoYEnY2BCH/Ec6jrefxAoQxg7wfkfA+cxa5+Y+IKJH7I9klQKYXQpllFycMmnGKwU
tUSAd/Lty1p5VpGrisKNfL2pWy2Otd24O8xKS6bke8Pc9dPj1qQBSO2CpCvAkM3mOYz6jkYPwZyK
Zh4ZbX4yBsstI6yG938yo5jUjIKz78e+UpXRedeWtbtUyS2+wItzKtH4KcFAI0Cg4f1Mc+qGmsGl
b+DCrSDtbUv0qT5r1ho01Mj24v+Ipdtf39acd9fjGEuxIcZFFUgFbtAjD81FIMXU4XUl7pjKxUzF
AmVhBV0XwP7E6BNqiHFKVAWdPU+mSe0znrDCOoQW8FIfb/JriCOwSt07yXJOhxqBo7qRdcnQDz1t
zEzH89pXrwM/vz0etl7Jww9loGy3w50xZkSSWNXhnRQIGlvFmRelVndR9uyYqWHDAcqf/WuBYps8
SEtA0H/nWzlbt+3S+gOw3agIK5l40XMIaMOgXA4ho0MXCE8d+om607MQf495FXkQK1hcqE5hSKZp
ruSwuPyhUPiv3jN6dDpPUwTWkUDTfCHLg8ZeJvtjn9rl4W9+hvf29G+ANLl+yogrSAUbhwoh6qfb
AzhIl60ArXHt8dodIB6sXM4QOO3rOmffnPCDGqqhh7ioBZF6j5HKa+UZ4B96/2C6FWk4yaNZLudy
Ydi+YFekYzYdwKfx1PeFS1mNC1eVh0Y6qxYlPT0GLOKuJ/qVIT+zNvTdJXgLfJToZA9w/Q8kbfCU
1uI057sN9BwMBbxKn1zWJC0Yz/MJkIQb0rvI8PaciU0/St2Ggx8f/dnY7SlrkkWQ5i6yNeNd3Zn8
P6sL57hmHl0m5T34v0U5B79klmnWWzsTrC8/khVEx8lJVuY8h67+rNRl9U8DWdcbsmNh4GAlVPrH
+oJQcSjpJXfcIp/ANl59WmDIoCSv95DbBPzv+2h9zPaHufElHZZcTOprvRgBqEnye50oYKQpCrcy
ihxzx2675Au8LhlC2vCOz/rdXjXTDMkgx02f58vuyizlkcuuQx5UtdzAzvOkxWhCO50yhHdwQ0GI
hCD3vR8RidJ0mxtvNzpZ2pHKnyN4aIFkU2CzrYu8oU7Qo80CEfok1VOQdaHbq5I48gIGMyt1ssXz
g7FUr13lwUp4L9ZNPKr01htu4XbPSenbjmE5WW2VovxMcxMSiCD+wSy5c+GQ5LM/zewlEWn0aLFt
cwUWX4MVtLB/3XlnLh4GCUKgnu1Z4Jb1WcoGokqj4Krwas1vN7WX12SY6XTUhrJ38Z8/Q/D8+k8C
pGR1zK57CrRQjM2HFjDuVzfnm2yqQORyYi7gk5Pr8AFxEG71NKu/uPfp6JTtiE5n0dEcJDdsPqJ7
hQS7OR6a33DxhElg42xmdEnDsXCU35tubD0X0oXcKMjYsB+Vbqkjj0hVAbLgcariCtntZ1SkyeU2
8Qe9YKs/CbTPnEfQsQSB4ch89mVrGkvHT6gjvdKXjar5AZOUVcR4800WJy5jlXK3zXpxY6I18ohj
H1KkklxZ0PKU9blhaejhV+IXP1S61lhfFjkb2o38K4Mlb3QHmjBWe3/WnIPOYkITj6cETn2C3i5+
E7UeXweRjz5xUHBMobJ8SFMH0inLyXLPBay0BJS8fQBHvrsIzIS91CxfjAVR+02F0/GAU8OxN/CA
1ln3uaxFtQtzyHAfWJLMdXeOp0a9HylIR+jBNyzb5wFilY8UoNFjcYx1WWjf1l7mO4boY9RmSUJF
Kk1/cBbJ9pke7X2nBf9+23uoQOm11GtZiHv5dFCj3VJgUa0uQEa2RRDLwf65lHNcKWEDvcuTpdOe
x/+vRY5DGc9S7EDx3om/FNfV38bFt0sXGgfuSOtrSMoXaexvb0q5I6DwHPKY41sRqWHYE/RjZS4C
X9m806bGCI9wKisxbjY/s616ky90cg0sanm+l/3VX+qo9JGXsWvNlp9RMdRlpSlen/aUX29qUZRo
iOg6nwHzuVZtU3b79dQB+BlE8A1Nq2vCOn8vy0O4yUG3yJPJEhJ6cx38i4p7EK9BufRQ8kli22oO
jCaLNnvtLzgwasNCXiNkutHvAX+CGREcz5YzZZgyT9nboZPumoFTUp7A2Wx3vWzgS37N2ugtOreG
Ua1ei1ss7x8rLRfh5yQngoPU50ie0b+fXKKxwhOr90oqNp42GPPwgAXmLYbVIQswpb8BvE320vrA
G3MPcEjxqhxyBauLQb54icI5wyfrwT4483aOu5tK2znZcr56CS3YvVzH7IOlzEgjG56O5skAqT3v
d8iT14hU7ZfajOcauyg9BfBbmU/UvjqqAGW9KuG9qCXWFOKDosS3/83v8iEP2W/7YBSX3jOtM94m
U6Dm34hdhxpr7zk6Y5mWYgn8cWEvkDZKtGd8slsNszPqZo/NrXO5Sv764GDpJK/4jPdrsfq0eXVB
L8JGlb3VBDvdXAyyZQ7LU6ZaEBW+q1H0gJT437HLQlDK924UO6fcn+NJ3knpq48Vy44JeGx28bJk
+7JzVrxQScz/6b0sBG71wjHKWZbwmrIoifGYH7O04wF2+1Vhvv2TSWRK7d0NUZMGGza9g3IAyIDG
mBB95F0t2wKKQ4wN9DguNK130pn000Tr17f/GzUbYIPoSwntJfFlGjotdPofRkmn1MobkVgYFsNZ
w+A68OUoV2HusurMFtRN6RnYM1Rr6SPtAmDuGmQmCW/rbcgFECdjPJkh5Tou7wF6t3VS90qw6WSK
87zzZy9hV9TmNxkuEojgq5WCMluNq70/2ysrW8JSQmbH5x2eOlp77IhNr/ePxG6rbpCnYV5DMloR
GrmnL0hGO6phojJ6p6v+F8PMBsboN3PvHZ2KVy4pv7lssNDcMC4wyG2RoC0VUeM1d0ObMp2kmt/f
ifXtImp0f9lhAXGU7XrXyNHlkxfSYiphfSIgQWDECR/UccJm2dS8boIPcfYtgL2WijkFkz1JOwU8
lGAWLW1XWNH0EF/zv9Ans8cEyHXo+BWx93rbCZlT4pDHokK8z8yjZRxYMRf6qBDdgydQ4/GO1PCq
d5/jMeHLBi5R/E7/R/yhvQYvZOAV2Hn7tqwxkvRm9fWxKfktyr7YJKAuJPoiI+S6lbpvXmTcG9Uu
ssazBvBgn7RCGvgsXcnmvdnn9d/EAWJ0izax6sdVuwmioTmhGBuQGlYzx1W7WPIWA6OHnywgrreM
aXyZapbMGYAhCUq75VPf0kCH4rJbKTAxHFs6DWCvLve3Uk6k2JRzaHnKWbu2dqz27cWqBB5oCflN
Rq1UNfryBa+uCdwTEcunHtfhRnqrUgxm7pKLCCIkubbM1TZxcqIIHNpywHa/RVhKSZlbGFUyiCB4
p7JlpJya+SrYFV2vdc8Q656ZGmvZb8fXJWZ8E7OHwdIeN/mv4E6dIEjHxdGuG+BFSmzt2ndELk64
dPqZ3vtuKltqDNGhppzgsgGfiVFPLKQ6VNR2l7ZkNxB+F5Qq/GjH0lYEaWfVJu7/NCmnR/1OlSB9
RUSraL9REE+N7RfMNgdAII1fyK1gVyvOkc+PprQHYZ9Hu6dCQytpi8r5ridrwZA3kAhXhFPR4lKQ
MrusOBtsVrCjQeIYaWRnCc9hW913/y4Dcn17+W2txaOKu1796mdtEhC+XPuNYNhcoYYq/AuPAU4F
igxDTXDfaD0bZK+WENZRC6GmHhl5NpEZcIM61O3vJVn5Nnk0SIwJYUf5QNsFhfpx+2Hvo7w/m3jb
0pc/uezeLR2yfjstQ4sdPIcdmHwiSCRkZCB6EpANwI/eN4HxBc3v5OSPfXM5wa1FANgjwBGcTPee
yYKUye9Bl/AO5V40Ae1u9SRbEECZgenRnbV/BI7Di2lFFExbJa9a7N/Q5D/6m3w7eIKQHzTniwi8
U+Ns8fxZxpILvio59bSEeNaCg8F3UN0B4PNcnpKPxnEp9wqv5qRN8MiPEJc9fGGo4NTJO1meOVuv
H+lWevzvldEROtxo1c8KbyKfvJLunB8c8hFeHgyGV1WEN/kstvdzVbCEaODHnXqEndQ7kH+lbMUc
X0Ae1jZT4SVPwjf/38c1He4PRcX7j/lZIP75kse3UqSn8JaJt16Mazuh0dR0gU3e7Xm5pl05bARh
7TFcuEvtUc9v1dxHITfXqlbu7XJ45ZPYLktzNSYBdz/ooIiw3Ad5HiA98SfbeHk2Iw+dk7elOF9w
XIz+xIbXeOVmR+fmA3SdJq1cGU5aCOjIQkd8egVuGS/IqVqvY1KWK4ipx1L8MbeqVlWSq0svcFpq
lxos0WBusnjjSkjjuV3uZjCUtUHrAGJ4p8c+Qw+oCBd0i1mtAzYTyu/t+TuKkI8cKQj8WckaREgh
5gBoRHOXUilCnItpnB5HfwG9NIz+HNi2JyZla3y+iArAlfqOj0kKKuHstbzDod5YxAvzycnCV7Cu
GFlU8xD78yPBX5zEscJ/9FImxTfoNcPE6f4moC3fhEN+4emKqKWEJv/k3y4YEtSgbF40Va96rZDN
3yNEaYIViufccKWlBPvyBDLfFoiGZxWjZnlwXaKOBqgP0Xef4UtzJd0jwPVgX9AOby7CL+9hYCTz
wpUtoAXNPqGPrH5bnMKL9JfGzYXXrlZXhQn1Co0NW/4FOs1pW5ucRVlsHRp9qjuFqSt5HbL3Jgjo
LbbqqDnhyRX2x1WrwBTpZM/btgA+SdDpAr/kHmoQtRKfIyJH6DQdpPrcn/96K7qqk8LdKkg8jCi/
12EkapasPsUodNxq9s0e4WRVniRiyFIRCf4jymKlfoHLsMqn4JtMC3Yh0KLwfvFeDgIyCZRuFaDh
CL/9DwwdPLg77uUGpv4eomDXBiOzuhQgZ5lqLlmLfjQ/fLcUAX5JjSgQaeJ2vmgOtbuZw9VfrGjN
yPGhBusUuRdiI+j4+defyq0JXFscqz9rcQc0N/n+IIsTrtzbwODHemGY8R0o5QUs5XBsQJ4dEg5r
hpeD8EQ1lrL1mw+5VQBeK0EdS8X6Tj9s/lzMdOzikS8iCuhrkRUQjYCfW81NsbIsGYc3+eSmYVG4
CMxZaKQzuYSB4Jz1T9NYJ+B2CBMwe0Md7NcceTWm48udbdmttGPVNP/vdo9zaN7dnL4DWX6PmaxJ
4n1vRVS+91OE1DTo07RJMOzDc84t6hOvYoI+A0bX3HM0cqeE/7Gqv8YRw4sHTLQa6hwcyk9BA/m/
tlOfgZ+JfrydwS5ZwSbdQ23zFvEAv+zhAPymgpO/r795cDJmrIxe5cielK9OTs+qkgiflfTq6htX
8OkxI/5CoQNbVxVrpV8KvPt/dgW6/Vva4rZerMUH3QNoWfdacPD4/rfqgJDuScL6totLIOblqPuI
usMTS4NsgAkLnJBu+EVtGmq2yy1tfKAlfdMbiynHLNDE/giKBPZ4PgbVXkHULGgUc1prwqgH50LR
jGJkW2lE3N5V282tKwM61SIh1JbjCqEr5da4SKrUaXNEvTkFgyBUHKjfU/7YXYW7RCTVH2vBD1wc
UpBH49MMTJDxVkNKEdj/W4p4iyWebntSzA+YAEu5CmmGzQ6lHkO1GamfjWokjIMO31lkEUGqiUjv
XJbsfVLuIQrYFIlz82iF9izY4tBRZF/qF5wDRFJNzT4pTLwyxlamgQHaCPnyQVCdT7012RYxtBxj
/0ZX5aS+Khd+jOPog3MDAfXad5DCJe9DQRKSfOo6zPi9F/J1VJkU5Z2gtyQVZSfM5xQM6xZIuSFc
JdqVhNKA9AGjNhq5qCbxoy+nzh/8UVwijou9/v6pdvZynQUbYlaIhPWJ8wc1nkcs8WKnP7aiFSaJ
Lqefbhlj8FpE3vdvHEmjNXANab0mo0eD+bJYkmGxEIf5n6iFDLv9HjcKwym7eCdZk38KuVh9j6H/
ek/w/Ofuf+xJTIJGvLG0d1kAEbdMAk4LMiA5zDUZ6PaUG+bxqWd1SzqyjEPhQDsj/YY2L/etUxj4
aSDeqG0HRXfbZMp/IUSdfOxPGchoiaq5P4qP/uZt4nMWjRkfrsKcLcmpXW67GTpRHN6Ah21ddmQt
ApQ6RgORtbDzUlCApV/r+8h9/S9jmqMioa8HRrag+s4fEO4G/DkC7/OBM9uwHMx2DVkLH0fBZbt8
g0U5fov3iKGeQtqWDu0ycDAaLoHi/adoH20XKZr9fD1bYPNll2RM604SDlCbuPTnIygxizxc+pjZ
LGKClhUnfVrtmpd0dXsO6FuaD5dYDY2kJVvCmjSpzEoh456QjN+0MhHLchfeTP6X5bNabizG8SUu
XhCEhUw4aBYgSRVeR5nmmq/hND6qBV4Sl3x29/rsWagPcKwaB3oo71CAPKMQZUS342zZv7T5+Puz
lGgLhHSj5M6D9l0NUSEpsCA3xh7KJwtS8nZ4bPPUEQ0Jkre/rIDE6p0E5bcX9F73I9psQfss6P4r
il7cSf29EoyMSDwN4SqRZFe5i2+BRn1rR3AnVQkggG0M6V+CL0qalySSTq+4jxMYA/omI+tLqWds
oG7Gn+uvp1L07sxrS961Izf6ob5FU+kKJ9G17zUiDLEgSnsLdXHglkJmJIDrulQnkkjVUgfVZcT+
LJoJVe1zteTmBJw7/n8+KJAs/phCyShHV1/Guys+EOBu9QEWPai44WO1QQAWhnMs6753MhIFSzPr
YLlTjIZkomF1k3rY0lkSPVIxDWeWOKkZcI+7aGPHaIoP3J2QhFZSIkHu78l6ncCXLE0F3aUiRzTJ
aosTJX50fajqCpdtG3Rpo6931B3lb8vwEt02jSWCRJaVwWVJbCTRhBb0YGmJu4/CSxAlnNrocnSv
Dhm4lwqBJwUV1wLNgQD0Q6CkDalQlmResxgkSmJBAXiGN2YOrFD7YSQGnCssEwQgOKBr/jCnMoSH
9IH7Zcug1PzxCihkGJakwtzraRUGFEadqG4NSdsuOLbXidv/ynxZGLXtkIDj2L+TPX7vLG0Vickz
uVPNqzGaNjlu9fpt9kagdGltWOAIgGSomu3qK18uccSvUg3QGt2viK37zaUeR198W+PHv9y3Nv5C
CGIaz407Sfh5AjHSHbHM5ler+jVAtGZKPzMZOlIr152TtmXMLiqDu2Cdn3bpZ8eL0+jWxohzSQJ9
Z6i426wSsiGRbvRZDScaaxURr5xeaFuCejULfIvOdqvRAM1HxV9sXPlQOWJdGdZEAOJaKx+HhH5J
ZCNcBoJB1V9TnfZCE5mjqzr7ViA5WGhQXo9/trIxY8ZWDtf22ihhGTXHItV8SFme4T+f33JD4zJC
U2LDlGH0VgZ9OUBALdUe9wrBE+9KK9AVbIuU4ifgOJtoP1SjvziEA70u+cN+kV26cNyVQbYSaZW2
IM+hlPk3IZqpUQlnPHU+OoYNtEODg5iLNcnGRTyydXI2j8faMKSQF8HOmAFP0sns/91EC61jVjEo
GEGBvaNhHxRhXuQM6SreJoCs/WhzgvGF1Oc+XUCJt3h772XnPdCN7qx+iviogFCaLBRmec2tOgfI
H6lHYNEPhxIfyzTtjetVeiHu1/7VVwUmiy6nr/X7+G8QiZ+GWOKgShj7SjRrRUE1kwTj57VjiyMQ
QrpPK0bHT2TRe2tmCMGFFNpIscWlVUJPRh/gJuPhippt0yF04E2CvV+SOeNvSFZYjB1zRLiFsEZR
fXBcCOlpKep9Gj/Ot4HOepZLkUGQ+DOn1sExBjeFi6ANXQubbD83RrCSsqVcuIbv9jfMO1+gDTWw
fwQHvzwCeKpHRnU3MUIcjy6L2Ga4SJa1VDzZRQd/Ldx2MuH8km1vfck4J97wbCyioiCweb5q/cLv
CcJc1Yq7vfeX62ECG/H54KKnwUbtSo9EkaCniJuTh8HZjz8FJrf0umu1ew5PSbOybPd5lkOXKrKh
oyzaBzJ8CoXcmOpRXicl9XemBWPsMgi7ntd1pWEQI6R1yllLX3NOUbh+8eUALi42xO+LB+9nOq1x
BxZ2ZPmd4VeUAVKlqg04mKBIIYskMgGdDBrHluF2bTL76GMJBBBlj3+7rpSI6diyyVb2TmC2InTd
JRpEsh0pRvoMajqArpOsd94s9fLMx6dnfzuW3ecvLvilcV5K2iBGn4Y+xqnpjjnkd9VfrTN9uYfT
KbBGLOZn238jaXk/x0jlR2lcIMb0gDU9Ii0iCEHNs20hj5E9yyUud2clDjX8TQGRT0Kdt/YVOI0f
adaXCG7twYG+e3C5rNloRzC9VsBpPw+pS6QvhNkEHtJs8rrUCraJQJNyMra7dPMyvi7Aowsh9mzD
ZTQtb14SjSDWCHpaW5TJSzNSFTzPDUlA358BrMHAC0ehIkM1kjdK+Qajvu2Q41HntXUfQAGqEIap
rgWKZ0wAwVcFZVnVo8ZBLZy/RBsZ7DhiLlrTIiu4hGhucX2jiXrKyyH7AdymkHoN1PQyYXX0pibp
KHpQwiAU5HtSv0b97rmA7QsduPHfETxCCm821W2NHzjIySxSu4wUd2gl8UiYokuM1KNI091xXBLP
+x0CKnktx8MuSLbR+g5bf00myU290Mxr9jAUPrP0at20mDOv43BnnU+NvdGRx5lW+gofyOvX/FHi
GWzb9HeOXSrvlWEpo2b/u0Qk5xx8QBYsPb+hnXpQwe1duPLMkxv2/HAixH1L+X9ygkRrMedUXiyG
rnV8Z3zDcQMML3qGwY8Lxpcjomh4W90MuwHWO1BtRFw5NFZH5rnmRDuU/xGcuAkHiTg6BTc0TMF5
ARpuEoKp4l3G7g8edN3J0S5izxSvM93VclN2cfsiQakKSi1uXIOIXAmUGhjAx3yqpH5QhgY/pkUV
e8DSoaT5JORe/hE4YKuz/OtwhUFyzquMXoApht8SShYbVfyq3t4xhuKvQedjeUiucrE8EYecY+Oh
afTVlFAafhwRTiheM9SL6/nWpCgx4N9AmeZb6QM8P22qoQTBVLGhsLZ4P48mSQ57wlv5cA7qmbSM
TgcPvJXbq5EftMhevPJB8cw/f2RIYqpMShicIdH8i8TxGfFQMY2gZegOAoaTUcoGLnt6cIGBUdSa
qIphu8w6hAagVSrItNM2df1H1e8e92LcUuncI1P7HbdHqNK+jBSb79vmuN0SwPa1QNF7DI6vYJd1
wtE1GYTq7a859RNnPfbXQSsRUaLFY8rj/TRd5YVyyUmXZHxyL7EHFy9dQQFB/JrKa5B2sxAQcrfO
ovp8m/NgAZ8PN8BYU2FC+lK4A3etBNncA/1LecdmY6/3lApPuYC03ReUv8T7v/7aZmKK83XvXnk9
EOGeJi1GCFgDy/umWCXmgaFPjuugl4eEiMOy+6uC7RSvu9v0cCn9bpfI6Bhd9+6QAE1DnfYZmgoB
ymKQxj71n42sMl9oVgMhDtv+yNhY7WSMxPUNxZkJpY1U+x+pXTjR6Y6d5cENMZiKbnQPigoMHPqE
9pkq5TSMU2B+Gr2qoWkysjAz8psFu2E1rYUvclzGwGj/O90ozIHqr10I5PDIjJ3hbCVPmrIlnwsR
WlrHo/ZFVVAtptZnbmws327XEBy0qcZDgLSMiWpFmDCz4CnZB8WuoNT9E1w+ZyIS1cShI1aXw414
xsbAcfFapBVupzjP1ANfO0T9yRTnlv0+4W+0FSxHfkoBPbi/83vqDw9T3sEknM5COZ/dbbtg6ZuX
RdlWppgsyGmibaUllsQ4bt+gln3irMFoamL/HXvlX5mRw7XeHpza0Jimx2Z0U++APgYFDFsjLXO9
DD28oJ3linB7BVqWntsGmJKIzhk8FXtfiSwQcQr/s9f1RpOF56A5EIxFaG7q60rm+ztVulvU4a2k
WvxB+X/aiIMqFLCfhh8KoQcoaru5mtxgBi4QO/aX6xO53+BxzuGuYrQptkQte3Hq3YFVSwaJD+he
LtUZtSVWtJE3gJx3hO+9bzzhTeuRBlwbw6uyfekQL/QbzKeGW0vqO/YVUxt65mdvSFMT7E9db7pJ
T/1MahqJoywtM/isj5Lg11sIbvMwNyCFOcqgtewOPjEmWsFqCiIB7px94mpncT1LeCk/FgnZubkv
UJLOtZicG7dY2YQrEGKS9ruOrS8xsdV5nJlrAVold2TMjSp264cB5+NJjSCRMnwB6pmpiD5dLBd1
OIlJ2TNpeual61jCyl/tikqoV3xfNB3Oay+cuUxBCW3ZEEznDk372Rwk2GGFefBPYvAF5TIooX8N
poJ5ZGuqmYfs+FdxQ4l31XKqtFutnSUI0wWLP4T1OFuTStnPRqzz4+dYcpa3/olFjSNaBz1spnvN
vpR0LqzkvBmeO/PeyrknfYYNw537BJPP9iqKxLSREBva4OJT8lc1M8qgi3ODv3M4DZ7RFDixKTOh
gYAoS65qoqfhUrtKLwy2Ln8K3E0xWcYOpard3LwjU21doZWpI4bjUoeKFozrjznx02V6AJ5SiPZ5
s04PWZbmy8bxUur3JHj7LMwZ3g+RPX1/Wc3WRkd4zViptfUWrz6V3lSCyG64ZiTE89Swg4daG//t
xLRfSZEeaZI4dulpLOWVUryxjKo99cHPtaa4dGs0Ig1boL6VuOFEpI4oj+6+O4AyiANVPHUBdAit
MJVzeej30L67ZBYyhhRzV9604Lo9T5y1E6kqcK10Sa6JTQcT2jF8k/Z9bGd10HFgWTct7zXMkRuE
9AsPar8qOaN0M1UK6GhMDFsKOEjxAUtZbhoh/BmR8K+1M45FCVqcUzy7yRK53W9IZJB6llXx9QZw
xvkY7ZlUq/b+ab8hAyFZxfvy7vgPgYeDEnZSfimnRQIh9KmRstOdQzv5MzwhMFcsEEL1wRU3WXFr
1uRTy2QR8Xu87ffRyhfEnyBiYnIVMQ9RwLKfRKh9h2vYoQaUud4W7ZoX3odhpRrQcdvEvv4NrFm0
T7XeGuGLgBQOhWohue/fmCdffhVAGsCxVFpGePvR59j5ht5yUjvxFHAAWCyc9qj46XGKl91rC+nP
cszHNjAXmGVc3SvBu2Mia8J0fNJ6Ct5Bf2N4HhH0oqEV5tHxKtjUKFTtCQzafl3aiWck6pbt1P20
eZfEAAfvMzSyQ4EH87+j6RuNOng75Gv8vFkEwBI89GPaYvq1tof4WOBJKGtqn/S2Lch3eNZPBiK5
w1mSo9J+XPcvRwPWCDOWtFVngkncerfucPNpoP7DYQPmC0GUIyjQ28wZd93IteT5JtdRdhrAjCU7
xSfsNVeoa27Q5tV4aUCFB8yFRVYYoFBcQ7r3oy7JtyMSRPkaGli/Q3lnpgLwL97fQlu9jrVZE6Ss
3On44TZSF4dKfX7opt0tlaLZtufrD1tlqL53IaOXsy2LKBe1wmwLYJ0U0bNR5j+CEp98xKLFDpiQ
ZwK1/3ghTO0lE25ZlIQv2zcLunnoypXMNmBbMuQPLiux30oJdB9xCrcnrXPxJNZDqzdoBO9jUcic
En6zvC9ZLNQrl7mOK8pd27h2kj7YlcgJHe/UkkLB/vfnHnswxbVHArV5jsRVzPIiuG8E40h7/16V
zvFm9o8q4xs8p9C8J+Z1BoEmyvVPAcotSK0qfGjemNt2D50oEj6+o40Rji9XLEHprkWowb/Re40h
AV08cvBBHyUzEgyjHj3g7ShHi/O3qhYvbhKPenjjaJi5O9PEVoWuOjLyRA1Gaj3jAirtaKhdqPpj
jFwJGKIjApyHfpcEeDKptfrxMQJgmEf3Z9ZwsyQMdH4xjf4D2Ea55fA/u+gU0xNOSjV3wIjWN/n7
Vaz6UsI4jg10+Nwuzx2ds8OOhBx1cCsNisxldu7RbuNCPSNnI5pccWiAbwKdpTM2GxFaiu8C6Azs
T10V64Y7rdvu8yAtDha2OOi6Fjc24XXreTjV1U8gfGtRSgaGYHGTsDiLH217PwT22bo/Ble7sRZJ
tjhr9JKkuGzLxIuX8zIHZHWNJPb7g/WgDV2C1wClptOAzDpQK5giRQWLFlaCEcIPliaLfo3w2Jwp
zsHkCuVs7P1d3OikVntbYLWUmXe2QNi8/5CcOcZWCLQSXygi/MvSIGmIue0AleOi4gaZ/LjWjrRe
tr83rvUVZAUzt1E638nAyUbl6AvkyO15LVl1ZEpkOf9lM5waXtXHpOIf39gt6nOrT+HEwhNKuBOx
zj4t5S6NW0Z0D+oa6KNX0i08xXg49Fj1cIpzntYwzMVMdIrcJb6gn/3WGvh01noHZHKFxmPwL+si
84eu9lzJgEJXwUnQT2tU64jrRF+PcGyHX5PS/9qt8l/2MW7TpIPc8eUPwjQR/7dwVL7Jeuq3kmMK
KPczuxvo6bLzE7XKVWfnS9vNXIe6BKwPUUPSzyoYoIQ+ddyHCyJyM1W3jRjcMQ70384hnsUq2wSU
1726kUsJNate64U3X5bdUzJucWbLwyV6OG5vWjPntMNBGbBVwnsTMRiDxeWYW97ncmz/wDEJNdKQ
7aTc1GLkrdwKgBZqEHQ2g783y8Gq6dOl9Iy3y+weVtQaXnkCAyatMCmhQ3UtHedUiqED8u2Sjpm2
MDn11pa7RokJOKO7jaQkirJN2CHLO5QllKKPQQHo3EdKECWTzGMY7nZ3Sm8ujnptCiq6aaR/bBCi
Gu5QYBK6EUvqS4T1yBw0q1hDMxnSiZ6vleTr/bknn2Tq6GhoQf33SVOvNNv1aDWzT6zMWe9F52wi
1TQcLtmxVvOS4BlaMSDlSD4WU+mzrcjxVR0H3KGfWN+1KNZyNlYIDDdv9jpTmN218VBfacKS6Rpr
loWTqjZX3bpC8VCsgGjvUzikgfgu1oHuApZMmhE4nKYDSRW1wvxXulEeKb/QHBsdeWIoTLdu5FeH
VAsB0VP+VJP5Z1uTApkjC10Nz+zDhWClP2AhMBcmcW5gXPmqa55AVZAR7VWvG5b/PXc1T2aA4dgc
6ZZ2Wf7iVOZ5t6mOfpkAkWAvLNoVX+px+nlwEPcqgQRkTRNG3WL+wX4M+YSsh9j4h094nGpuUGIJ
BZGjEGFLTM9V/hwJMa8hUYb0TZi10oDMfkv9CviolruSL8jwG9QoQfHSZiPj74rnoO3aspPFsPI0
HdI/p/aNHruLugZItgtWBFGrTJLM5GJYTMF5ERie9cMSdGlZinAFn0m3qfqsLH8MSWof5xONmI7e
W8DdJKkzaw647To3w98ZkwF7dGHXnf7+2K1ztawqFtSgxET4sNjDy68Gg5I4u7RthEhtjzXZuqP8
3DLm4n/Xr9aqRAcD5hPq16Ai9HbBbo722XTaxO6ZWzbn0pCmEtoyaq21tl1/MCOJUMDwvy6zwc38
ES8RWJ21nM5QeBdhi+BJpukKwnY3tgTqIfZiy1yPSvH6WbwgZuffkFlNhTZOLMbjSeCBcFN05NwP
NMxL1qpOqcCFvcF5R6W7M2D0zI5xcxt4rlT6dbbppyMBlrr7gemLPzY+vEH6PXsIn3x6gJiSJ+QB
xpskwkj5qvINrnH2DQn70A7j0QUCVokFL7HF/TvhrKeGEZAz9OuzTH1scX/FEZWOkkOKkB6mmNeQ
PkxlXvAz4ffQIiMtd4HNW++LQaYxuEKvh+PVySibv9nXpJw+c5qL2ednHp59XMUPgDTGlKS08HvD
0TjkKtcNL+fCOTFT8MsjGBzpDqwMjhjxTdBWCjfrc3J7fCg/tH8ouLMYc2oVwOcVbFtDbVr9kLj5
fOGZaA246MPiNxo54qUDusukn607W/U728CaKrmYIo68nut08Tf+gPNzfKn7ZdQQLs+Bv8i/sGrs
P7JL1F6VDNAoPdTzZSSfCY0r75gpgWsMAMtKNupv9chtFCJ8mU9C6IzUlkpNXbVz8sMxEs9v2NNK
IOyhaGHxM+qY8df1PkraIMub8WfkZU3i7ck46RW+WW77sUBOjrgcH2svFt1oB5ZOWZDV7wcLIVqh
kNASAH1VGFF97Zj6t+T0OUX4fzKj1SO7MP5qQni1IlKW7cJyc8sIaFy1oj6qBStFCaEOk76DXdrI
Se/YZWxYcxa8mJ/W5qF8do7y8yO+rue98ncSjqpeIYRA1T3Uti2DHUE07gnOvyeEiZg23J9thq68
fJq26Yre7VOjiVXdeQ78OH/ObgtxBPRhr0wqKikIU5r0yxXFlBkCgPs3khy3nhoWR8QQoPMqoPWs
2mr0MVtNvqL3WY25TtQ6b1cJIE2l8bl/PjOiOpYnx3HhmaDyaSNVo6r7b+SfZAF4FgMkn9JwMZgh
pIhWEoVfCCwWYWwQgigFvgq4kcbyL0tg/6pzvddhflIKtcJ+3hz6XYiM77YSiob2NSyZ+JpOR/5G
PoJM0+hYBYJaPTJkkWnMG5STPtgm31ttvEpvW5yPQdt7CtvQKDkDRzaAAHDQ12NYTMGxzyP/WetY
4iFQUQCo+/i30EbqerW4UuEQSVuPiPrlfZypUIeRub359qtZgXpeH9DI8R+KVij1d/GeIxo/zM4+
GrpkX/+wBzSfrHXXkP6L6p040xFdc1Pw3y6SdSSQLJ+7UkANxBIzXGtO5dhAkumye4W0r4n8m6gN
9kAHJykJ0+/PvmZgNWlTj2vC/YR5pREUoJA+Km2u9QD9VUZwNExdH6vr08ianlgg4+RDyEZ1nCz2
5BGZwZLZ/xiYvlB5evJ+3+0VPsjoDsjB+3+57Z6lPVYkoYZnSB4gDjvWY3lQYdP9AAJqgdrXvVEb
uF1suTw7bxP8au8g7Qg6T4fIwiq9zWpuwH44X/Z+ZMk1Z/RjstvdzUPEKC08wJoL0xZqXrE7EGhh
EqEzp/H2w2a9sw0LRhp9YCtefr/aniINDWzy9IJCAbvab3lRhj10prA4OkC+TaBcbJOtp+hdPs5W
WWNQQLMqdnlRRDHhE7y5CGmz6kTRfKzBf/xCz5WklNEeaPGnz55Z+CqU1sPSHA8a9tOacNUfo0ZT
ksjwv3UhXWbaFBDdLcHp2Xkv0YyuvSDGRPy9Zut3FJmIJxO//enlJQd6YZ7mH8Lqjuho9wGYgxJ6
NzDAOLGFlF8gWF5Cw9s7cVur3vVGuHD3JB+VVwidwFCulNoDU2saAW72mdM6jcrH2YBZcG7dxgZe
LhThaXEfXhxSCvIojxu38leN9NLaYAGqmIzZz0VPUQzTCJQBcIEOYP50l94JnzMeGpNZgibtKXr0
6rfIgG/bjEuwAfUk2RRCJFbw9QMqL6+O+x0Q8ik8wHu/wSm8yaMFgjzT2ZPAbzBZMtBlg6e4f8AL
Uo82kyp6ri3Aemuk2V+FcGGItUk5QmaNWUR4VTkeSjjZuVnery6gI9g/Q+fmu57Qm7J6GPew4zAY
2lxAYCbmfQSIlVioConyovAs0wiaiXGnB7TmvdMfiWAlWv460b4IcHxlECjZZsaoAXtH7NL5IMOu
O1oQX78xpF/qaBeAE1uK/s0MjNWaSzQgMG5GefICMhE5RB1ppV9ulP51K+uWK2HrdgZV7sxwME4n
QLRXRvDEsbQBAdoE4fv63vsclhr9DK5+iElHjkfpF/IvHaAOFL5XjT63y348qhmVnY8zUJVydJi9
IjlHDR3mQidsPTiI0dIv/x5QAZJALJl4hKbg4ojDwgqkWuuGeBzcr7xydffq9wRpxloX3XW1Z4MO
9PQnR+xAKr2yKUuzrUA8YJbdt0FlD/4NDmeXLprxcabch169DuwBf0DkdK34qivpHewTys0Dr71x
9Eq1k/9bcrgDnf7rEbZVQel2ZoMOV85tQHHTF9Sp1FhjAH1JcoX6VywS/XgFInFQMxoYq+pKZzKf
OL8UgYm4Gpm+OtKsXLbtfSvFNeCfAKFlvOxOjJzIMdqVX2Xwqf7Nw758RVsag91E40KN81kfhhar
rPUwdAYw/w3SRI77JwS41a280FJ9SA5sQpAG3fYmkx7gQLn3tAVzuk1cuxMcyF8oN6BrEgWCTpOr
Fie780LVEey3fKjjC0ggWRmuKAvM4f55WsLh+LLPxW5hek9XEKxbaBnMBp7oVz9FgF7o9LOcVusn
/7JDZpRmLISZ1Byu3eoz40e+nH1ZqeMdA8MHFj4yebLOCa9G7sUQbh5ECSy6+zP5jXuhNPuXnH/2
C/F1OGPmSqeaVfAwyEkU0CAL/8EoCsuwf4TU8l6/a/aIQq6nY/Qxm5gOr+zqzkExIFH2uvwrMPZU
gK1hdkv5lyh3U6gdk1mFZZAPWnHPGLy/pk8t+Yzfb67nRw5BwSNx7OqDIHnCOGQA1REd/Gs5MBUE
Ri9an4sRByn1OBZwM8xW8w6IjQ9u6Sr4DPO848c5/OSeqYzRaT+7c90ReuXWY/zTL0dMUD+GCDgN
qI+TbpZgooDybKtwo39Q4GJh9J5XdHn+uVCX59rDN1NS+jCLgfW14g9sZr3hKzVwxqOmW4EZGrSF
EJU79IqB+uyACZAefgYij99YZAGy2k9NDsgJhIueJH6Rnwl645tYGFjg16A18hiVsc+/rhbKM5Ri
4e7bZBqJl1L1LOKvfHM2coiZ5NOUCrq3MsMeL9AqTAKKAj+mHpK1Svo+7QqZKkTRpsCUv8eMHsY2
ng16Zr/udVhSKpwh8ot1T3hxEdvXwfFHNxGmEXksCGwUtImOUlv/t0CMdTowJ2CIY/fWeV0g9b0B
6cMqETqjSUCw3v1Z4sPuc+S0EtlDOG8fH4nWb/ZEBWzyLwXyWvojBf0ls1QqI4aZPPal8MxLzarD
dLe70mKvtufNEVplA1FMK5jRC0vviGc0bdDj7BrwqxunOVqX5i852P3yn9G6ZclB9p2r9vpD2YeY
U7raUpjQSqbn0To30Eg+s8ypauDjkycqHgNSSt/ExfDQiwjpLvOg99wyu3h/66VkbcohaRrR3ERW
2meNENoeHb3sCcvouT2ybOBLR+TLrng9E9bNSWiCB62RRKuEHM0bHgJJx1YyA3ZCvvSMiSHBKSw3
ql20sppvOdvoRhvUp/XUvq/nxk1KwHg8KEwDxHxoVtVr+SdVOMMQS2fKDd3dw+GCrW6aREjvZrzg
7o6SUkvzPCXIwJTXqmcvE3CXaK2VppZs0KINQDHRzN9cSCOY7NTeF4uKHYIrGpUtDv0A2DdKoRDE
b2DetPIT1mUSaOZwiQyMuhyINEyEsxwwWKSUQ7M7QeDq287qGZXWYM1yKKtdGVyTIKyXt9mugOoq
2M8ytqBVKvXiKX7vddPRLEyECH19RTm6sHsWhgQW8ARAT5NBpMfHuR/7r+eCR0Mg+4QAOFA8fG7Y
IBufT0vy9YUrI9bi1u1VsOCSeteLEvmxfx4i+GLXCMh7dJkIAIutOasgXvxhjz+mMjeLDqb3lOn+
h1Ee9AQIa++oPaAnOSNsnGoipbfc9VrZTrmVCZ8+k+GraB8n5kb+RNS9KEuoQ4/tKu/D0m31hds9
CYLuyrGe0C1+HyPKKwzwpQi2vwky69hV61vT1wIW/2XLJUSPkSqtlyuaw+29elCZqVAXWge1UtbP
x8bE9gNJUaWzst37XUz8fs/qbZX5DHbPjpX+zXjdGjOugDRRu5KHMUXxJL3RcLclM50iOqpEP6ue
lp7OH2ntiY4vC5fWFOyfgfaLH3nSwUsHmsk3lGrr/NLD5P0vCHpLVJIjG5vGK/yKII/dhVhFryJf
RLwC5atWFU6gugCVkjQh/Qu70O3A/2JxkuUKg7VLGkZUJXlWeFfJ74RnV3ri6ZSO5u/jSpIlNWB0
Nl/+01XwMhZZMm9TD9N3XuJgjgmwQxRA1Ngc7N3PcNAjqQ1xzqBIkD8CCeoV9bq6xvWQJxPg2qHA
eLzUxpUozdUgcv0R0fqSZ8Qy9gKY01oWEBcgrs4vlsv+cYUKAx6Iiam/fak6GQYXhZNmXawI0z9X
Y0zJyGkL3fNvCaC1KgHni81QMIM+hH2Qa72tu4L6S4hfK2FmEUxD/oozJpW/9IstFAIt8bGzdmtI
5S/FU0OLz5WUbDQWI7vORz1ypHLNFL2h0RTpMLaEtp5xkbUe+rnb0n9P8VhTOQNlenRbxcAlIOdZ
Ig4NlT0yJunMH4dBaShcsVkQuZ1BeBlDkUEthOk/grWn2318HmK7Zhr3m4FqYQfenGeFGmGNilI5
w3cf89QWXXW1ZMSysD5pwu+/LgcEsOqgnDkJmU+wYSEBbdfa6iqjVHFBdIfyOnhBO2sY4QYRA/W/
+CdolbcGQycdpffaB5Z2Dq0dAR4wCIIzCbqPWHsdnn5nVW8Nu383D+L4Z0IOMVKzKG1M7RwsV2Rr
XbULDKgAPnWqGVnx5TF923W1DprCcBsJvtag/dOyS33r58iFY+K/pgAiV9d9P0VAsdpJYOaJnBv2
N4goCasBMOiHJHMveDo8ePkQFOoRHA+CQotd2BWBB7GGBAJXDlWJia/7pp7BA837K1/OzTPj1nSh
4QM8PGJRhgdi0SR9lZknGBEvXShZY0o5Rv+2DNpsuGszgTQgwnG0sKQX0f3F6gSLSvRkKkvcL4yX
GQ7WmJ2/WrwbhOTSHKsH0ECvQAey1jggJLPMqdnjhq61wJJH3nbPMds59NcNHU24O+WFZaqI2d3b
Ed107ZuTM6aytA8fzFNj5X8pkDmxVw2SIYervH/+/HOXTERpXI2z1M3D0ieDW5d4jJ/2vESendEX
pHZXy+IFgQxLX/M1LH+GvLAfB7A1OOF94mSMkXOLGOIoixjQ8MpkFYf9WEcV+VlZzoQkzDlKaHgs
efeXocQ6Jn1q9YY2q26HAI6flJLMB2+dz1V5OBzsb9qHhebT0gWlSgXqKpnLiS+mJjwGDqYEq76g
4B9POXfF/CdDqYUKPKlpc43RR4xrzYfIHVvjZ1Hd+OezBX/ZukvxBRc1Ljhpi6+cCuvTbog7HkQY
Tra3h2nBl3N2pj1ePQQAvY/LMYUfnSTAfk/NdlXOWo2+7U0KFbt3g5b1gf4KabljDrTeluNIUoHg
AkhhLagmaN526ezvB2PvBWPU31EUbgfOD3i6qpIfCDpv7NNRhR0S5v7CQkMSBUA3saeySYOpjz3n
ayNuRVohcxqXpd0Kq0v5a4KhULzQolVT3SSepHLe8dCDs45CWC/LC6Gn6lv0YgEhMGLo9KiyqVqa
CE6hOq475/MSr10q5JPgXVmeQDf3RMAeqWdzuhOn4oL+t2A51hZLnSCz6pQZqbjU+G2yU/9KuAEy
Dxx3c5v1sSLs1+th5vGa35xU8vgQclIDQ+EzdaIn4IpQqNB9MfQz1ppq4yaxelE6JfUEIGgnyrFA
FKYoRplhIWWkxZYp5AQU0MuMN2xG+Jvo58OuHZtJzk8Z0dryfabeWC4natHajogFXTkCsuPjA/8q
uuM41FlnIYCD4ukCS9yFadV/yNhHPjFlSd493Kh3cJq9khgFnsz/Ygb2Ke6b9zxJOwKwtoRV+4Yj
1oyQ4xEmWnQVDsf37+q87PfVRATbGnt2XITdffqKUD0RFUjpsHSgFJ/A4VIBIPn8oni56mSa0yKO
7aehUkVZco0XUFIFSMKNI+y6x2apHj5RR53sumJkP2bBWavn6i8cpSA0xmSV5I8urSbG283Go4L6
kG3921LTnrX9jXXYq0OAltKlKgm/mosAZfjuaVtdFBRN3S3Fgk/sonTLS5IYbx8S//hZ585uFRVh
NpAcv4Ounw80QIVhrfvYjFx0FYu4VXevWGZtZ5bD7oi+ABEDZSED6aOiClHfQ2tEWuXZKa9AsDeC
U3l+CP+QVkuWU/bGgxTzECx/89r/YjAC03/MThFf34j0J6vYRnDoUF6IdCeGQ9JqvgTTm6gKgfno
OgDXY7rvD8JpbCJEc4WVDUbNxn2LbyywJBzAl0L9ohGtXbzh216p79pJvAFy5/+ur6/STemhoH1+
FvpvAZvRlEfG1FJNT2mHJEDHp/YKiRSJr3xgTUBRl9u1zG0gTkFsliwRE8YlPclxAbJ2SnkheuW/
8oK2jtFf1oD7KI5CVFGIgHM/Ecc8KjcIk4fDm7JHVV+i8TkPimhpykMtTDc3KWSWYMFF3yOi1CTE
4cX1+u6qa6G3keVVSZkmUYKKyiPT1jOJh7UND5cAHtMZLW0Bh6LocPCpMgvbx4W/4ZXHNI4Knyo7
VvwBFJltXs5kaeeLV6yG0i4NKMoYfp4UjbCLeIMQMSy+qHv6em6a2FSt+4xQX80nj9dChyZ6/Qo8
cnpLwWL6UY8DRNQg+FaCAf5Yw6kASQwRAhVOGOI8AVcKHG+bxhfqYqV3fH0UgG3DLCzjIgkmozjE
hrfUFAmomqNVDwSRi9E52xdAJlOkFFxbKJpjQt2zTneJ1BWQyY/YoQ5Ljxpy0tGUP8inC5b3FsZV
6OJ0ysBcEg07hIM4Y5lNdKWFM9RCp3ewuE6Fte2XtSW9n1PHDLOVHlE3mYJoneic95GjAAr2Xwp/
Qm0gRekVA/NjR1BDi74j30YqkK4FmiXKhyX38vBLplEdvaKAzLAcrkvob5kDz+URvMD40LnSwalY
djJGeVBC5TIjoh97GiflA5LrGeQ4HO4T7+0M/NqM2rh3fj86LCTzwHJOegm6njpb59gPVJTWr87N
7Gl2/driv2m2AdeaK4xvCmKuuy9R+p5DAJfA8PZZuJg/KJu/unNZgLkc8qQSCzJdodgmqAlBlaTC
/2VhkyR1lMfsDNxyRBrCjLsmh2q/SA7vkUXvbx+ynsIKp8n4bODVjFh9H3YwAjWK9VOyx3YKI9nm
TsG6YBcFiNlZrkKKBlT2qibyWcKnu513qVUp0UaxYmwDz3UMqeHW7/qY3v26F49IkLNsIw+ga+sf
cqrmeIosvXloTEzREWzClg/jy/o5TpBnqDZEUE8sGDGI2ef9PVXXQCjPRLqoS6ZyIYJxyNDaT5kl
XajmztKsjZF3YyubSiBakhZ9N4X66k8b48irQoOYIadsBrEfmTlb0bzSiV7cdyTebFE+vA0sTxJH
bQja28BalKtASjUV4djcPaJ2BpTmjvt4DN+US6fcbMzPm+Ily3wrOClNNMxfav4J7buNyfM9Yh/j
tuPyn18tumg0ti6ghv5waYUYxJIMJHBdhZMYwFEB8LT9fqVGS4uOCPe7VJKMk9cjlUt2ye1R3mht
L5h9XZIrR3XZAl+i58P6E0JM4vzz6WfcR7RdycEq3GjoQeQnMvh6+I1+tHLLP3lqTxlVVE41a/Uo
VBoTCusme/T+izWfaS44cnqtsDiUQtsxzwUudXnS6vherdmEr3RofzEe2oHmQ1+I8VwZUmSSgprV
LUgg1VlFjUfuVZO66/zACwROqRIQD+RUomth7dcLoa5hXBfEVmlxamc57cDIGTL5YHQk6GkB58wR
2PEcqOOlDVv05514DzGNkyfqWNW4e9dsUsl2kbfN5CxKSfQaSV7J/+LpyV4enkluPvIIXHCEi+k7
jFJOn/LmkiNX55l6kU9CE+Kr3Q1S7miFa/WveT7Rz3EOUCFUn8mkfipDCG1ivNLaflHdjcncnFSK
9n7j9vdoL8DObltiCcxNf3o5udGnnGwtc4jclj39MGOMkKGXIIL3sQNAHo1iwPNUcRUx76F2v981
SEao22FIB3apbVRUgwwjZi3d52t9/WK+nHbdrCLOGgRZbkGI7Swwss/Tpau8VQs1B1LwCikLDzmW
FlET2+3F57KtPbqNATR6j7SF+LxXFP/WwXi+iIfoQWQl+Q2GeUnJ4xUspnnwSv4VaXiQDL1ORQou
/NFqRNVerha01wT3pIBeJDQ99DdoksFKnAKgH2FqIuJ3Mbz09cKRCT82abIVLaDIXUjFw+C6c2Y3
Z2fg4IR1TTVjo4rRa8JcGJgwFYOf1KdFL4F2tq4HOSPQ4X8wFTuzEhGN/sfi7iqnOeuEtoQnHKvb
TY0gfI7OQQQGuxV87OMrkpfRX8aY6L4iCyZvRilarjg1pxk+UjmoTAcDGhWlatg56qZsfKDYPTQO
URvTxlmbJSGRkR92XtIKxFeOj7Ah5Sc+xIXvrpknZlxXFvwykJjIP9dQNrPv2jJnjsNeSe51nK0y
Xe+7/DEXa7O8IdJiXT7Cybht7CPyk73t9yluPfTYDSKj25C4glC/8N+NsCWsfu7djHbdYa6pw8PP
Ajcu2z1adhTv+yUWaESqiTsj70byjWKAUEEAMeITYmwgtk+yPP+m2sNcIacq2MmZ+k7g3DKNf/JQ
IrkuGe4JVah7miZHEzZEzYM42lxqzNRKd1kw3x7VVghag276OW1NsnSvyDNF31UDSFzg3oDZ7Kzt
wuRSX35WFMbzKCjBmfFIepDZZcyeNdIysg73kcg6rdnN+Wpfmf0CdiRznEtocUikhCEQTavAKzaH
W6CPE+QWHGcIuvE5UHPs+jLz/SUMx/9gb6dEVl3q2r06udFjJp5cJoQjp8ZiT1pXqp9/gCp466WM
wCYU65GxRfZGJCUeqFna7ewKRbFa0XPxsZa/HpqpeOjpW5pAEZL56bGat65Txrjc5q2tuMJPq8Qz
KztA90D7uYM/JuijxlDXocKv6WE59MaBHyioyMqaekI6DSA+ehb2/I7FJN4p8N1OUPm98jPxcVIy
ReBvN1a44ebu/dY/Ari1ZpV9VHBX6q5P0s8SUWAHoZsSanL9hm4oSpXj7DYgb4wv6qiVLH0unsgg
cCmbgvRGDto195VTnW9i4/XJxjGKdyicif8EEsXvSiNVKiPVNJMa2b0e4eWzn50W8EAxUXFjV9Hz
Aq+SaY/JmPw8esfS+zc5ttEa9Y2XZZotlDQszj3LYdBjUcMKcefqycV6Ygd76M5PQwBDMJaVHuhl
n1MRgIR3XnRhVbeqVZ2zLim5gPd3Hy8jT4V8P1BalLdLNyvZZQcfIOXIlKWVFfCXRTeKjKFU6X+x
qzeQdAMToawIAR7MU2fJuJifw1frv+2LelnKL0Dw63wg8P9eVuqjFS0xmcQ+wPChc/+yHUR7xu96
QzCJfE+4Tybq8//emqLCk8zvXK/fdcPrkiezl4cS7FNqzcv+7X2UJpnDHGyGQYsadbFeuPSveuY5
abMomfS/ASs3F+7vyf9WPIErjVJwNJ++Rn3eIbW3EQsLeqmdrWBQ2zRcnpQFd7zPryoSONGUqJJ+
7EmbXU1RoiXBWSG9SdrYthLAPHTox7cC3r2A+78fv7yckvQ4H8s43jzKrFb1nAy8eKwy3I0Z0TwC
3Wno9As3Uk9VAvMCrJlbuBL9l6PB/j+9e8G8CBuEyh0YJnkB7oH3uGlFdfUzX9AVvZaW9G3MkV3L
2C3A/A0AIanY+Ry36p2mvub3g0r7XUEi6rd1an/u1Y+l46Hvb6WDzUEecH6KEkgI2fvB/LvQrzEp
zVBEVEEEVicisiaqQ5OkQRp9MLEfOeseZIy0cRBjKTTNwFFSK9xICCwSnyYnf1q6hzXuni8xaCQU
xMiVV31dRm1zDwlBGzRaZ7Bw8hmikQCqwVUF0Tu+9fBxDpDYnJ5ziJa3JjBiaiu8YdZI20+KyoAs
qflLAh4VyqyvrXebmslw96XlEkiT0x96TRkyattY2rXmLrrmpbJRisvjfz5EalNmlEQuahlIG0ws
XJmmnlHUeyF1QYbS/+X8/JB9cBLL/nOfpED1P4tMTWCrh60svVSVkR4vEJ4XrgO7svIGIYIhms4i
IFeCARmAHa1dwlA1OCNAAPBfQbt+FhwfKUrwvJA1TFXTAnE3dVzGN+Qn+DqqFpQLQthdBTnmkXDk
XbmuXRN+q8CFtcYUkhLMEfJpZ6n4uPgWosqM8XEz7PPgULnWR6117kGYs7bsgOYRxRmt+6kWTP4w
u3gvE0YdLDAVNbOphPO4tRyoRWMBGt6Iw70XVDDwynsorWw6NnemZGY+EKk9vwxgwWopBgCIFGRM
Y229iD7XwIccsCnqNzwm4zj1r0NE7crmZ2c7uxtGw0y/2o9b6RIDXol9NjryhZMtDgmV7l6vcsc8
R5Zh6zLav2EJbdZ2jW12xelES+tuRXfs/SakEL7MFPrA3hywmGx+by53s0eTxfzp8q2GLTQxvZjq
ofPG27bO3o+SAzKs6AkqMxlPs/QnjOi0ahYumGIGlSSJR8AF4I3e7gd0p0KGiyadi6KbFiFhwxzm
yc4KXSYyVJg3IXq65ayW/4cMWqQ0h/m83Y0ONyfDlGoafXIHgyunoHEYR2nfDoxa8ctrwdLt5/xd
ZhV+1ePZ05DMfvfN0WgY30T+wHE6PdFvgwULon4RU0vS+C7/km2JZWX9WzSeQuXUuu4rfjnU7uwI
aYlLeHgIaKmTQD8GC6AHOppkFJoE97t2qLDbTlVP01Vus+TPU7g5DDXkM0Wd0KnEx92nYlS9RxiT
Tf47I2CnL3zJpAPXcZr6pZymWVsou0pUVE2U6YamgseIEFSzjk55ounyKk+MUEuVBCkmuB90qXus
SKpsrOBYu2KNBiFVNv21RpKV76q9WPduske0Heyx9vhdc0L8DxbXn4Z/hoPVRRse7UfjqObhpMox
uPzd7TRbTmX5ygSo4t2t5dL4XnlZHvj7bfCO7Zlv8APJNkcv04XmnRjKArUA+eGzFVwvrWIXdaJV
88OQJFZvXIXqNS9bulBrxHWAxCT3jrtj123bdehF+yft3w7wEqMACiHbxZoaMrU0iaI6VALODeCj
yhqxwfnR8Aywcm+LOb7+x8/VLMCJdF+29nDltyNsfbsQGCkU4r2OP7epeK3EssNpa1rNGg80duel
Xf15hCyHC/62rgtNeXcNDGzC5dqK4fex4B5emndj4Ihu/gn8Y2MkjNlX9jx4D/iMH9cv9G8chIKP
Xpsr4WgfkYfs8LbzQlNk+BXCc/QRho9XLXh+ncPgBGU20pX201RECkIi/IMbNNU5lmuVQs1lH303
MD3i5U0bQucSfa9VwgVTa3Cw7LP4SfLUQmTknWBesoCzAXejlPRs0fBrfdyF6f5azoUqVggovX97
oBt8xF8T92P9GsJlq5siwfLnVblZyWlAdlGA6/Jt1jWSfUvf2al7XVk4GezaxugvSMS4sW7rYinX
RS0XUmx1+mWvup7ZkRoRJ0ecMC8koQsaUIxJvH0vOT8jZJxsByLAAcES/CGKGDKALspSxMNAprUb
JYZC6jlY7/o9myqXWxt1YOwYuF9RzmEpN/3VRf7B/VGR1LwVTnunR8DkhGmgiGJrHbrduy95orL9
x/w27Mo42xAkxyG3VxmHKpZ0XYdJYZ7nHRBzYHqjhhwSWaW8esrqUBt+hgDC0grvW84vG5kdpgCz
Jqgw13p0q/k3jh7sR290j4LuIwnwe0X579Z0yparvlJSZQauuxqktMuHH5gchz/v/JNI25u9z3/H
yiyJPW+pQWXYlzredqlSnswJCpDmffAD3RpVWi1DCoMjjWzJ/jGWNmTczIH2C/Pgh+Fkiz6/5Hy6
XoVQDxLf9WiJS6PTe0kpOEGgMIuN9AvVzto8HWgTmB3EiE1U7Iv7DAhJsxkyQGgigerrgiQ7P0L9
FE15ECEyIw+Zs0FbpRgKb6K1y+5U6OtRS280Wy9MKeA5s/KK/l7eUdFGT2dFc1yyY5W2JFFVNdt1
b16EHBrT8Cb1a/iY63OjWOHH6D2Tse3hDbuS5FXC8SEWbn4MPdvVT97sIN3S+v4KMFmGSskxz/zI
zFI6aFlic1JCnjtzl8ohJX0XX85ZGSseyHGJXk9hmhDVS9Fot40t6oCsdrVrO+cnU7qzUxVDSZ6t
19afTBVj+H8CPvcV3bEfsJLsvrt4IGwEpT4FXgTCZq3MNSTWjIE07FSJ2XZ304PN51/OxBdiek5/
JegBtn+2o9Rcx8DqkHAafFo8V3Ely3Dozmg8G7P4rMP5yeS23ZcAzcKfpAT4DRb+G5CpJp5JHlt9
KbzfymVcsyo/x9ZQzXJnhbW+2XRcyhsCtH0L3P0rHRWDvKG45/Uspprb2P4BXDGN+vHnSxG2DfX+
4uQeuHwEiqW3T78cE13/+VbMwN2t7KC8wQ15aJKFaagb4PGO+O40y6P+kiXxajuC9yMvVw8TH5ek
/HrWwQetu3qfR1G867PI+hOebCsd8t2sC+uCErXRoOKp3zPE3uHbartImAhisd6PRvoej+2/bFCy
U5I3uWDkEQDNKcf/lavF0154a7XdrSpAaP5eQnTU0YrGiOXtsTHAQrEQTwjMQunMyUhQqrYUtEVe
YIVbaFMg7ekzDU8TlSj5qpqR9eXayFo50j8RW8T7NC0OK9w+viJKaP3mgdvOjsygypXjuTT2mBNt
Tb/3SskhM+OFag+HvhBL4sRjUhA7YQixs2R33HiVRZrdb9rhfLkR93FMzBeuqubik4X2eHLBHLns
H+toGgrPFzrn1DeKLFIjZ538A9aEzoRPSqO4iiyb21T30n7S1MLsbCTe7HGECV9H4SBDr1EdJZZl
67kzleiUdRdRO5gOMFlX2803ygBs/5HM5DfKOrRJmgEA1EK6N3Jfv6DOHzvUaHVTq2ydX/QaXIo3
m3KnRkpQHur0fganDUYf5bfvk2PMhjIo9jc530PbimwsYX9IH4hqeViMgXeXThqSU0aztUaTWaEM
t0BXPN8eyqpGfNJEOu9cQVnGsrGPimJz8sKMcZpxQyC4gLCat4AEgWZZak5vyv4AHnjGsvvHlOKu
bkiM0Y4Ak1R4w0uHFcm53CwE514GjzIkOd1qhPnB705lmL1gzvC0XOQis/uO+xsVV8CEreQ9rc18
sG+SHtLa44b1PCRQAhtmq7hL48Pi09Qt0JbKVXQfPXDc3axWF8prcy0FltF7qvVYznHutz8KOubM
sHm481OvD65us/n9QGaWtz0D9bju8Q5oTbqhnmouPdbkQtxF1bKpVYomQHTBFEV75S3gxPJNpFr0
FvMWoCFa2Lb2xiDi0qIqqoxu9VG2NtjfnT3vyzR4BhTsnAzKQJGhdOsiNRbRgmX8FSz3+PWKTflm
95uyrlvdoKPv3LUSXXOZqfqR1JNarUqRIOCJJ92ZMOOsn6T6wTfEtRGDWfTSM9iFIwS2vOczxLpt
qwzeM3qM1RTSrgBs1ISDOHSggL7qcbyFzIKJBxYiJiI0YE+cXNvBYRGVoq1xnki0h2y8ANJIyF9u
7gqZhQZWxwb+0vVnhKORWRfujub8sRk1dkfjA9o90ksoTXelY1K2N2bhbNiBEQzh80RtqhLQU2g6
PLr4SmbDcuTXQAUFtVukB35cEGdc+OemDDx2ZIXEC4lnQR2KprHVxtEseQS30VImjNUbkOt8au7L
2A11ILUxZbp/mKm/PZKs34Wbsd7LHNyC9rp8TMNLOZWZC1K6coBtFFc2E9TBGrx8RHAmkpPWuim6
XLqBPtavjOpzuOYgyLCunb3aDiwqyMZEnxUJShrEDQ7gbFfbPQ+0wV7ay1+tG7Cj48b/He7XUXMn
SqKU72nWbtwlHCO4dDz7D6Vi/7fj9pf8c+1cUu17kZalAj9aSRdtGxlOU0c/xd6uyg7wtahJTtdv
6aB9M8D19Pfu16mAE5MvP4f2JwbXfcR6+W4/umJQv3/iqEH/8mZkiV7LvK1O7LWgQPJoRzP74kqd
safq/L8g01A84ncsCOUoN4jxq+bowHofZ7mIuSF5bSA2S4b6+XfFarnzrpUtSpT/ilbq7rBcm2aV
1NwzeYl8GItZr6eZd0B+1dfA+Ls2HHbfoTxS/hUddYLIzEduKVox5HWzM1digFYQlME87LyBOgj4
IYVWDdHVcpiZ+1Q2Kq9R4pgOVXXCeULiS+VIcXAqczjISDzu8I7jm5DBEUWc1OO3GBkWuM0BAkoP
/EGz0X0p7k0qTHapvmc2sRLWYzeHq6UpESAXzxEYPAYY8VI7u+2qi7jWe3aVM3JyTK+jw6ton1F/
bAL/Btd74SZljczHYD+IFkbq5RRiFuOwhNyQCzyrCTWcJMt3nzKkNU1j19FCMH0GfD7g4EJAQPCP
v1mh7V8y7iCuItcxkSJgYk9ZiDtmgp8t/kcmcKnuDF+uQ+EkKd8LXQsaH6gC6uGuuqGP+xyxauQ3
GPpYJ9DBLRQTCNQN7oYXR0WrMBlBngkksALa5EzPueaU0payp9Kktvooxp9fGFSU7zhf4r/4OlL+
v5znDcHHeC/+tq+SFz3bMKayVTW2G1NIvxTolUCnCIjkCkAX8bbGX+B5FxZT9xEdS/FZPaiZhBDA
SLWE6AOEm/iR3Uck9P8io6TQ6Wg77iSkMybDvWyC+SuQxl/ftcqadQT3H0CwNXfH5wOH/McakZWU
gbxE7sbW03DscjqyaUpSAjr2FJSPC96ap5cSoO5ApmecP2/ZgEdjh/+ui4BmldxD4KtTSjWd1NG+
qBGdXDNAMgbOPQQ30oNvqxk/FlS7T0N5BjHY72APhdlf/CjXOU8isNjeRRnL14Y+Pfq5e/30noe4
MTT5SBWFHc2qxAWGLoF1a0hOD/Hl+ZTap/nQhyuiI+T/Hr1WXwue+MJfaINU1XfuHTxoq078D02n
DQu+V58keuOE66ze4ndmigS9lHxxhWPj+HwVMuUso7qmIxeatJXITv5JS+08a5vjMFD+ibqxiCBG
TwnfZlk0oEVTgC7gwZbDJj0NZjY3/s6Z4mTTmkRoIJZfTcyLsInt3NkrSMBwtkSnLMyELTcNcFrE
OaubVPnMGD0bMRoWBNqPDtmV2rvTHNDXzWZAv1fjmW4MeSaGbXPI2nNRjrx8wxpl57iF1E97vdnh
Lnv7Q4/HhX+LqS1C4YQIoPN5NIfuEA6d7P/1LO6gVYdtamBk+lxBPA34xQ3pRz+YDMxGdlUOUl5T
njnrJ9c4Hw5vWzJsF324GTPqV/EYw/F8Ces2+EoPTh6iG5iTmKZdpZ63DrTeD1iI/YFEumwVOGtF
J+2GhV79D6Kf/IHYLVM+sHi1CDhp/u/144p7hybdo9EbInPJiEnbbizwUW76Pmc6/y5kFT0aeLVr
Bg//Bxep+6S2Yo9MZ17/LxRxeTs8vYIYPq/IEL1SU7mxu0jgXQi/JElJC1oSYFM637gSkLNQQeix
toaVMpWHAYWmB+5ca9AbJAWhQ5BDupPX6nuMDCVbnsTESJ7z98uNq2ej9ba8HNuOXMyWglExQ846
3E62vsaicM4l4YO2Lb7uUn0vOcB6/qlzL1HbFzkHGgZWRcAxPIt/RenEyxZ4OFQzDG5EY+VFvgv+
M0CQ5ZPimQ9ehtlXxA7gNoUFJ6qhIJug9NhCXBdGQHaWuJX9khrYAJ0INjLWeCoA3/TheZccoaM0
v17nRt7TJges5y+lvSZrOq3x6/fv+sI+cJKsd5aw0hzDjBB7A51aw2E0etRGgz1dQVRPkedJEIrJ
MKRorH1M8DtpZIk8Sd2R5EgbLgYREbvK7okc5AlJsmxkCvo9FY3oNG6jOaHolXAH0D134TnlKeyT
KX6ZI/1z+xQr7+xWQ3Y7MN4I+dtWkw4FyGu96ht3Y5Pqrp87TMJ3u45MWUCCbXN/t4QFfLo29VQJ
clXQhaq1yYTvo9uywPWPOGc/nN9W5Jt2OdJgZ7OjvgnGInaYeU5S24YfWyQhWk3Qmwo8ANEPy/lp
y0VNwIBX5dnjP0uQypnBVuQJvrsJycM8EL0v2VINiuDWZkp/gi5fmyU00nbJwgM0MuVdyxY4+0/V
MI0YZhae6Rni65ly+8UmR0zhOBJxkcx9+8NlF4dt88L8WGwe9A5iMZolIcdrah6Zb0XMH1cN3A0X
xuoThbK9itCYeYcE298GF2a/uEYk5ZCWv7+mmwRayTmthmmpIl4i/Zm9bHXnQAcpszOTHIlF1zUX
t3GOlHpFTQylLUaYsmtO/b8JCfQWrFIOJMFj7tWTQ8nb0tZN+6rDrR3OqgNXVIPexMyxRhkQLsz3
iRwgFSrcp/Br44T2MwjjkFyLTlb6MDVGt+YB6shU9glPhivAtls9DVdGZXwU3Dow153SmXikwAOw
h8g3Q0tE1eDkmiYFbATGzDol1l7DQdEzvZxoicz6ASWibbjPnNXC/Sep7CbZVY80BH1bPFtHrl6L
alB0zaKrGPA5WnuCmFi9Xr6WjIErn5t6VWVaGt1AGOuFSy4idI4NJpqIWuugLokWxpE+Ay0ZhJzK
mzwO1YB6qUQmKbjSyYxp1EeSE3SujUHkw8nIj+WcrFl8lO4Na06OLpI+FqUQSrWzl3oU2iPLVDGM
XzzacJUm+oAf10xPJmltAtLKnyIRIqCcsdx/jKH7oLRcG+lcSF0MPffZa0xRveh9gHKQ8+UbNvHX
PMDQWi38V7IgQX+G+EUzWMbZon6pKNPMj4YazDrlDHttpuzt55lb4vJT+Ss6yLvcn/Xskr8EMht4
AL4Iq5Ad0QHf36MA5fPRc/n+jh1MYPhTU0h9klv6RPPkS4OkfSxfdPkiRmkV+PRQK4nY4ydS+NKB
xjowbdfuIpdmgxvRArg0Bx5zoCDmLXlN2ipqTLRzu+9C7mmyvfiFSlSeqityd/QimdzCDDaA9YEM
x3Omy+R6hUWS1Ac5pfgFZ/K5E8xJ2WqpbSFvcy8tykcrugcsy3/2TViJlUAoz9w5kK2doXnus8Ka
GqVqmhtVGz2OE5IdVRmjJdvkxNwbLfsylRNXeq3BtFPizgYTmQ9knwqovGi9nvKkp2+C8MDwz+li
a9v8mReyLYyuunzfV2+bOJ8VwpIVu/s44fL64BoikO5bZRZTNg0bNgxo+DCK8x+V15XK3LmoPwlY
o0kfVQeuGNusP3MYHePQxk1ZWEf885zYr29UaD36GY7NlXhK86l6hXV2AFJgZVucCTxv/zTBM+ev
TDvWeNoAW6VoeHcCaDGnXJ5eBArl45r64G+65oDIZ9pmiH5VRORXX9M2L4dqt7Sy8eR5tfA/3dx9
+GTBuxuY93hMt78NQ0FXgleU/n62vTHMek9OQ41LxRaN+Qq4FM5aJ8bAOCirGs0Q0IFIV2AY4elj
RRoehLdvRrYnG8SJP8kAooxm3f+2i9Gb2RXPxXYp81/aP1tc+UWLT02JRstBwvFJVYEpD56/sT+K
4bWTllgknjSASYz2gywZnO/lIb0L05QwiF+w+NJKpowxFb9u7sEYOVL/eE4p7PmW6h3VNx7ZbiZy
pOAm6u8vfMLnJ1BuCjM39XFYSEyhYnNrGhJbRjsPoFzBkX4oqldcjxpttzGHG9gwjjXcx40993P0
EMYKaNC6VNAZ2jzlFjR0lYFl+vVx/ZEvHQ2ex1q6+T9tgl2kHlXKH4ZUal6H+cn54Z0apVVrCaTs
TkHND/+LtxHben15LIqvzDESGskIU0NJ6iw/UqO1mWdLc8f3TYTQgvfD51BCtcFeN7QOQdOPydn6
b9gz4gNw+j79g5JoMO4c4wbejwMjTEVY5jQ8Wb/k2cdzoG4c9gXxpkXbOd3xAkBGIB+TQNenmYxC
RMUAmtSTVIgUYU+kib8Y5GtwpF2KCjAd7VT+pvCLmKd5nCnfERCbp+auaX9i0MCHDf47Idw/rd39
WptQKfccNusl1ubyliJ5v0G+ezfZpdadzTx5vlpHqk/QXF4y0YpY1I6+R5u0YeQ0PRtfC8QrLR2W
jMmx/+DDeYsauRlCn+33TR4jrJrZ/vjF4TBU1Jh9BfH3ZOzDswKXJRhpUV6E9KipnNWunA1j8fTQ
D76lrnqoKDIYrFVOQ5tcA46hbTjzUUS+Nef0WM3vJlQHXXIdCOn00jAc57bQSJqT73vMc6DydiZC
jd3ccsSoSjrI48tOazjzXoOFDPc+XPm2F1K2NhZ+b304b965nPlk18N2WBvmYij8B6uwVT1U56q8
4Id6ZlZIVPRCysm4hhA/T4qobmW085qqckIougS1TBYkRP+LxBNqtnjmrpdiZeZ1N+9LaV/zsbNB
6jjDAUhhlxdajopSymG0VmdvXxi4FkvqeYrF49vc5sJeauPfLR4H7atwZ/XUsgkun149PPOmMJbW
2HFjMh++jyVjW7jJijNzqQr8OD+Iw+QI6PuPfploYCcRYlxHWAshVlME8dV5waiu1tL3wQRp2LMM
7nn1bv2X/iqIp+kuwHbSPL5uVO9e5eLS0a3e3B0dX+/TxBi18murKRMPStW8n3P8zZE/laL6nnr/
lJBXzK2CAv+z+8BrGAtf04CGI/SdLNNkA/laUPTmXIZKdFwT0xUYKE6c946OzYxsFZmi+8v1MiVy
Tzjzkn83exrqVui7ykcV+8bi4MS9smE6RFT3uFtm+QoDbnoV1Xu48L6dZ4DxAioR4hGP0SXED+va
lCHS/Cpc8MRmGhYSHEJZ9YV9nY+0wXYsFQV2HXfkRixyzs4pgE3vg22jz3rI/AFKwpBq5sU4RPcB
HDXNgBKH/u2gUOGo+/i5QIdNQCN69FsHQfH8UI1bGFMRL95y+s8P51fw/VrbHunK4RioKqp+uHpP
pEnbJOmenIF2s5E2V4vW+N/C9AGAD6B5MzySZ3FxbTFpswbmFhYaCfU/bmG2NhEz9L9Cs3clOzU/
RmU+TmlNbuIOjcFkUw4aZ43X9I1HvNYJcDJOdVpMGQ8rwgJVtrLuDVcQB1Plde6s0fP2AN75MJoe
eM6jDpSInV0Wq3esLAL8gKN+qkbzQnBxZg9JtwraN7yU5v0NABg+e60WHzdKnDk2QtxqrN59r8ht
FSTy1RJq0/ssHB5hRX/kxygu3dVK3bM1OYv7XJN9ke58oeLI0aajggmx4rZmBiu6OopXbzjwibhz
8VRyzJGeklUU0aVy9dTrw69vsKk3a+MRGBHmwvJIKQYvNu+kNo7ZXuqDTxP2qWp6PC82diEudO0Y
VpHwLgTlSkLEMhpS/Z33URw4jT+PZ6sHIMFVqiHaDFmOLsFbFhv/9TwtDqWsg8z9a9RQEZUe5Bu2
e+0+kCotP4NSxmXeBWkUKRPwcXUXXgUQB7gQoceawKBBu00MFIAzrUge4YlYIdblXtPhSRet4FzP
SGJ4RDSJGiI1/361tjKkJTIjq1lr5TLpWjeXHooFaXzJ3EKCaIl/RbGciHgvb+Lk3Yv0zymmNDLr
7zMoJfqPtZu4QRkYuU6WBdGKm6sDwYXy1FDkA/yO9psUprx1RJq97uwxZjuhoaGLAG2cIjkE8zal
9xVIRgaIwOKdf7DzTEn0BASRz/3Fm2ICz0TOQZc48Z3knWXsEwTKDv88/P+SUfC/S4Ny1JjKLV9s
Uw+zcfPJH3QOmogKRAGTJ6xHxfHMPMB58nP/DsXXovIlyUU87irt2hf5QT29rZ80bkJr+xzCkQMZ
pNMrZ2uAY8fZ+4bNcUmM0OnVs1SFgZsV9uLJvSmAbtvfEXpWb8INTxD1lq50X46gkkASgGFKV8Gb
QqDch4q9c7UMu5j9XsLSuEZVK50tf/RgrLUf2V1kq/fg0ik6eWEcG/gUeXbxR4T08KTAerNQtfxg
yvG8QrXattP5KapKXyj2WsxdfpiuUWKLssfNxn9petlS5luGZE9sriZ5fHUcew7zGpEktM5CSEwU
yLFd5mAAa+SWDzNCPaf/tiYTyCuuC3pdgJrT+kL5gw+67xCwLpootNFCbdxeCKyF1fNWbgkLNnhP
BBVi7JDMQzGhWmcMlSuSYVvBvCXrDn8DJwoibAL1iR2SVfHJCGEHUP62u4r3eyMcpWiLeokQfttJ
xmGgGpOF8rHWGuRS/69dg++5/oQiyC2jIwWaQT3wa4iRQ+18JDFmrlUZsLO1bg81V8136j+nqzUq
6gyEc3ZZjNkbsa+f+CGpoliJaalplqhtm3eph3wF89nFBbAqAtvJL7R+TJWcTw6Ml3owDn31Uy36
YAIORH7MYNu6ClkE6vAaDAW4Ymz8beanMc6OsnMP16u9mDrR0gKYoSEJG0gIuNyBAD1dJ23gwg0z
G6cb/H4Qu4AIUSJnZ0Ml1bvpRMTx0GzBdrtHY5oXQDDMNjylw2u1xRuId1efvhac1MVQ0gk2KYRd
KOlMiydj5O0PkGOpfG4PGL+H2Vh7uqv+A4NmcUv6EiJ64uGq1s/OD3RzT9TJsR3M47KYORVNDMcw
2C5FOEC+ssu1Qfzhma7VuiBYI3xNNuCrQezm9DMXa14027xzKzsp50+/+EN28UnIQsr1U/KC7sPw
gdkhkUruMIaY1Q6NYoN1r8M4K4CgiuxNlR+0YxX6aizdTsvpxHv4IcAhXSMscvYa7zVeMO1VDt3M
K8wDbYLIP6GCHzCIDcEjo/LZiE9FVT9YmNQohBp5pfNDS5u0gPZ2EvTrorFjaLWo9U+K2BgypBy4
upOf7gd8jJ0ghHOTTyUSvZpI2XV4n6lMFZQeBygDqM8TradnorE2RqMfQQ9o389ugCqj8T8nrkYa
k40nQQJ81irpOkNybs4ppGgWOh7xVbV5lYsIAFAv+U/2qIB+UwRPVsZyCzi/EldXTlEja2crWqks
R1FbenOoTGus2YVL7ZoxXIBqm4z7GPY3OwoEjiXg7U3JSTS8+DCwoStvM+E1rJVwOLZvFntRFvT5
1GUQDGRRBwR898yJRmA2X1K/8aw6BruqAIffvCJN3kbGK1fyKJGF+RgFCeSzAKdINevXflfC9S5P
ve7rzofuHNcBBDa+iK/3x5Iy3gsOSUNth9ANC5eh0uxlrgJRcTasIyqBnSVbd4p1Ijr1X4nQuMs9
OIrB1obUkhoA58jeFmhhGkVZJjWqwk1+Z1H7C6R/ZNpwQ1kfddUbnym6QuQJkYfXxKDRISkayJej
6adA7BHM/UEw/DUeBT+dsS3v9UiRxvb4olTw7K2kUGOjegzFlzns+XlEgvvxZzEFYd/PWYmaPlmA
Ds3gq2uPCc3nMV6ePA9xarSvzKdyHJRVTeQaq5u5jiru34rXC2++uGIuwboUT9zU1Cy51UBgQR8D
bmgWcgNdbgR0GdIWeTxDN4dxKxbb6w8g6DtOvdyCZOR4Tl9zNTIJGnl3bs1fInqwER6/AtW+EyjH
q5X63FA9LT05FXm84v/NlMEiMDMx7rHR45czb1zBAHC+txHn4v6QfukxD5K4q7M+YJdHRrsqWlkA
w8PEZHGO1C5oemZYc//Wb8KNX9jdQ06lEbRCAnCYcFFm6uXSmy0QxNQzGyLU/cXsNsCSz3Bu4W0b
sJQjrmoC73AzQ4uMWrOav+OrpzcZZgyNBSNw0kSdTzAoBmZ7nqtXPS6ejYNnicMwDtrK1hIQhxk0
9d0M55QfTvDevfc2zJh6KgW8166UVspz4kliq/Vn8uJgl1GtuTeg2dQl9vuoFCP2Ntv/JPC5V6EN
YUFfmjv7JrlagGtMrP2agk7UpFi+kEHGCj6lHjxJcJpaUudXGqeDJvOstAiXDLIHAiI6ytaD3GOc
Rg4eufK6jvhC2J7QOz4tRF1dozOQFxM9VbOaQnEGUHHBT562RQx949WOdSqKeFNyTp6Qdjfb51iz
l1Vy1gvhvepZFXJ4ScSIKq5EgHoH/PhVuN0IU1ze01a1ClvjfIRXhKYuScnB95EnqqtA+/QUGJQT
5b35b/6x08IZ+HcC4GyEwFu/wS+qoEcqCeAds+MO2pwlKoZ9jlr4oVjXie6GX6RrMHPbLSPDw61F
zGEeTW+4ws0BccyktHpUOaiyu3blYRdykHoMEaz0zxUsoN1xAOsdkd2RAAnKf3qqmj/nwkyFVVc5
1PG3gJHDAGmfusMmwQ22+gzZLOriEV8o4jes6l0Z7W2yryNG6ck24YLOS39ZdW2gbBWePdOTLGrc
aUYr6ZI/zt46CzMtlZhASqOOlJm0rBtBfR7Awa7eijDROPTXC9AUu3+3kI62GNDjw1wKvBa3rVgo
4QzhCKcRUH1WeeKpSDae1TslAL/ZK3ooF4Vv9DAPzaUaglIQhK0swg0kepjwn09M1aRuPbcJ0jEl
+rQ4RYfhON4FIuFspn5LLh4Pi37Xhr4Jsr/DcpS3cBVbGaelweOfNjKFDM5Qj2De7vj3ZkEllyio
oBVX7FyQXvDnfdt3MsGnqiWTMQiZ1pJyJAg9f4JIPJRjbqIg6GF7sVcBqPALpinq6R8FEArhHcOj
dMp9z1T1potAiMXb5N4AbMC/fpy3mer3vNRUhUAQ/pAofSE/wgDY2G3JNhJd9pFORGXUghU2CADq
E/RK6Wz9SLjO78ePO1BaOIjb5x81nAKlqTpTQw8xqUs22seOCiFyxm1Gm3ZQPJ0LK8KCfaVMi50Y
+p7VS4Ec5khfYJ8V+Q09dEqHUWj5LtzgYbHgmBp2oWvJfRrlEv3P+LvGC8mdzQczjMYUD754J/rI
ls3aB07q2+IfvBCiR1+dAB6FQ1QeGVZrPWilLV193RY0lBJgroKfnNPE4eXJAe7BWd3b8sV/oQJv
q4ao/eQQJ0WY1yqSurKjClohUiZ8l3Xl4KhfEecsECJHEJaqB5f9eXdAxuV5tla7z4ZAx98ahpJ7
buciRc/e8FlQdKdQfQYQKEghfF/SmVShuLZVkC7OV5Pv4Rz7kykh82X7jwOE5qxnhOuAtw03ROC0
Ebk+Z4vvYIFLekmN7nCw+ehe/m9uQvE/oP5W2m1CPcUdWu5m2MGy2/KOY9L4kqVUIdOWU/sGqfPV
UbTiMcuvUPeoQwaqVvEM03AraZmu34jzcgDnqCmwYCHMsvCefpT+fHqj3l8TEz7bRpqWmEt4YX5D
M4yabpH/SbJeA2OhATuI0sfLIljqBzKVXaCcHGjCSu+rp0Y3Ya6itsO/PWhSNS9EvQrgnwrc/98n
xE5k9IpB0hSLyklfTGEoTSnoNL8HSpewuOD/8/gd6HJ+tuvhNqypOPmmlYhvKThOfzG8hJ+eTi3d
XotmLk6ihEjeFSyelhy9gtxY5XOXJPa8Yg9whpM30QAHRWZV21NnrBi9xfxw0XdqNi7Aq/DQw7IZ
tuUKMjjM1jz05M8p2USo9TQpd0uSIQL30lrjP1umJ4j26YSrUAJ60BIAtvnNCk2v+Vr1f78URj3+
3oJNqQ3IMX+86+ZJsY5riTdGhe0dQqXGaqGHGL/sGW+Wvlp+Nzxey6hfEYj7nabwhSeUEiPXEt9W
PDIs1mqYlxpRSHoQcK0DEssmmhK7LScIg/CFHXAnAWnlPdMYN+7gp2q3L4znq6UzjPD7MaFa5lfs
d7VrgB2xxc2bTPjXUKurQtpKy5XAqb+57xAbDO/3dJd8fVyxtC3QV3iFvFKvevirSR5FVyQuIn4K
0QmxX34BGC8v0aZ1gkZlZYKRJilB1Tg0yavW53KOhIGV78sr0WNYLYrgzN0pv6BGZxj69EK7GFdV
ZSKQ7vUAQqXg5FVNZEDZ2z4+0Ogo3JHF40piw/TrLQOjPd14VUrYDXh/M6K738IN7NP0GAlqXrME
lnst6ovRduXUmYkUSOUrqavtPrTJU8VyaGXwgI4O4lqsNNwzs18RfhGQsPtu97wrIJgtv9ca924n
hZCrzkKULxJps0mfF4KL9cYT1svVmQabgHV3VZrjk9y1nR6oKfqHl26C8DTEN4YV04senpiHzupC
Gpvy4TmZaA14x33JkMVGZ9Fsy1pApyRG3k+8FJlgP7EDvurqjiLoRUcoOQ+DBpOnRUpjy6GPe+86
lqLmSP/Jv4m6HdJuo1o0p+rLEUiDmk0TW1NiOk2/weC6kTCGUSzP9b0x6zgXdE6Yfn2AncGTvbew
+YPjJlZp1E8Ztzbj6Z8fGzkqiUEiIRfuH0huiYObtBDCTPcimI4xW8SHjzFLP9EJTFOjKYAiKY0g
XXk/2Q57eTomFT/NNVEcq9LFUe8WjkM3kg57tQIciRS/R6Cvu6Nhw90H+EOw47kBWO+xIcHh2Zwm
qF6ucv9yBMkA08pNFuU2+d2hbQ6rz4oxtMZsiFAFmWHAcyg2OoSsQmkF4rXBIJYrxORmNz6cmhg4
7kqNu4jsnAqB4wrGoOdZlAudQQrE0zjFHe3Z3zSKdAEjjGSkL2040JTHupz/C4JN9+DgxTmXIWW4
E48EUeuHZjucYlfpnmDt8YbpkLjekwCfU3N+O6Hhe9snROTBlYn5+FR1hg+RnhXHn71j7qHLxw8L
eFr3EWHbXMQ9zvjBjpr3ToguRbiWflayLRKpYYJmgpuyT7nR3xwO0Jm+9kX8n3fyB6repRYpkMNV
RQdhxWY3Zvg8O6+FvD+aV4yyKMPm+6UY7AD3W7v9L6v5BSH+L7sS0NYvtoTp+dGVojv9WHBDSlI0
Hn45vwj1vRcpJhpTkTzoJw3GW7LyI4JO3F78JCorpEWiQ7ufkK3XL73l5UNYM03o0bTLHj5LA4Rc
KmVEl8aaytnfRJMKkFHDu+X9rAhA2RUsErQsDnSgIsrVJfqnOnVzwgomkfYbESlcEwlaTorKvXPt
pxFA0lBFyjds6cGPSeDrpP1bxOfhv/dk3VOwij9euBSjMxYEN2mIkicPYHaTC6wmRlgc3/o+Itzl
u87lKpnbV5oqdRUOIudrfG0qUK08eE8PcdCqtiyiKAzIGswfg6wIAR6/HIsGsT75ZV+1dAgu/ew8
u53QwuLJsBjh7hIpH8xw7DgW7lNJChPdYls/wX6nSnhhxO8MM1cQLDOgEr2XW22lHhF/rYTz/49w
G6NHEtXtc7/kZ5XzTHNS+0WQ8FdKGoQEbtaLiDfiSQj/fyEusbNADUlvBTSAB+y4nolTESxi8u8G
IDZC/7Sn7VYCkmDYwjhI3ov6SQWl6ZJuAiFlt9OnkTTqRFiNfoXnQbi2rBbCjaQt0r1dJM9DYeCQ
z2oTXYzrnoq83wdWPP3HaSIgqUFqzzOMZgZtFqeAwlacg75LNXdR3Q+xbvkAOIWdoeGYbG0GgPm7
dZ7G4dmWmPajeBf4jEJ8VMYtdbZT9q4Xt/981F9R0qFdhnNXfFgELwup/1HMhnwLoBZyLBnXhnJv
+dR5LJ1QwGZBb+r4CnWSWhMPzlbhPXiSp2q1NLqc0Yjja9jJeDPPrO5lyRj5qsG4q2UNKSAEdtjF
80v2+ApcUhvwTyuI8Q0fzidN6jWnT7msCGyrd8CkVn8fJhXfj/txI+k8ertIvnl/+zsYRSwNaZW/
0sa4+Xw3fUpoO1kpljntsmJRynyh4B/QCa3XEwzE9twQ0InQGBoJLSKOeSQwMM+LXKOb/D4+OCaw
rFNFkznsL5KG+anzzjCjjHhlpWXRu4Y99KuTup8ZRdRBqjPVxUIzP1899wypcBTiEE+qS2hu9gM4
UaBOT3U+qboSOXUIkTgdzpN8rPGXJYnDD8moD9T8OmR3r6EZd7+UeP6Oifp78l17WodT0UOe9nDR
lyzTokBVYs7aGSAFX3xgQk1Hyl0pbUN0HESYZCuJnXKBu6RoGbFl071B15dzwmX0mEmBnVcHb22o
2j4DJXIuGIB4UoxwlT5wN7aIPiJD+Gs2cVba2bMB63WmVZZi4o96Ju2u0XbskGjeYnjwGdLxbniz
5SE9XkJ+e98UAvk/6OLVewnx4ATucHh+YwyGMz5BpUkC4fug/9F3OmFzO0WB7BYDI5fwJ2g+CRNI
fFiKQ+4Go0NLctb2kFbYsg02w24PvieFOowIrA5yic7DkIMnajEQ4r2iy/hHBmpv8Z0T+u1ctK1X
dxXJFjfvDNlWSVb1rX6uF5QWNOJGGqar5b7otts1XSSrmzT7n8C9k0cdiuQm6eUsxaEuOQZhA146
USUzpk6vXq5nT0uObyhcuMDulyGwEirE65GPSLqH0J+40stWI/PlVj1+JYT8tI4AXzyu/Nqk63Fo
/5ApBiqKzAdwNiJlHIu/+kuq5oLEceb29rE6fCUDFwl87qV0Do0aa0WGWZHrN+7HoUn0YxIa5udu
zf8ojdHGhLAZk4SdrQxr8O6GJQl0tjCWsmoeNE4cwpZ7PHOuLagi4AWqji9WG1rfYh/yLUG6D79e
sXPVFfg+/7QH0afotBEHuQ9fnif+qrIhG6Kcp7snICdmclSjV/9KUg9wPeUdp9rH1hGfpnQULTN2
fGIyOtg0p8TU1lw1tyKMpXiAcRyzDPMXlGKNOwsHLoSv0HuCXxEXLNlcl9YMhseVpskRbZPY3CJ6
w5VCinTwoaQw8KVobz6pXfJy5Wz5cDaUdgbMcrr2fRe4nGBSzroG/Nn+aqAzVyC1g0qhWE4YeJW6
mwWneG+CbFROOwKOYAwtekqzVJ2okXBlcAITPyodO5WHGHD09mkpIKs7tThaRw6Km8f277YdjGWU
PvL2s/WZ3NF695bBi/d0mUVoEf3wklmugF856d5CH7OG62cufqS+EscxZRgNLea4quODV/febjLG
eAVA4BM3HUnLF0kohn30GGiVwzZPyFpVHYhz1nXqpmyltnq/nl5sSiSKBQGMyHzjZ9PuAdiA8IZ8
jZqGmPl6DNCFqiEThXRCzMx35NmJr+svHkHQ1XlQYHjI7sfaza8WAYyb+5rqN22foEt2HP4kLWBC
al9e1ndQYGKKc4owXWfxO2D2GO8LuPqU3kdEI5/yxjoF5l63WPLgJdXYj3YOC+4HYyNSVxA/zW0c
j7DFllnL7jAzOPVdIB+qv+EBRCvF087wChipHBAT2+O/LlllNVZWiX7FSi9AN7vaknYO9/wL7thY
x+VppaG+jNoGrpysqPRC6AtAovxmsjOMLDLkv+V4VA/0T2hR3aRn7LgiKXgSW40ZtS1JoGC7pGDU
husm/d9X9lxvlFNsrpSCcaCIBN+peiCQ13E2NejQlecHt2Oa9dRAGkd/FTlLdEYV7K2G8GxcDdtU
qp9UqfQ0sdxFPzfqI1cLilqxJYVt3kM3g4oErpyDWPQYpLC8Ga4rxitIiTU1l1lmBkrAzyODg2WZ
WcwNxZTEIH6fzYkMombhEc8KUv5TDRVgUrcdSbrRl0ZxmmzYe5sgh8CdK+mWJ/N/2DSz7dvT04r8
PBpMI5KG/sHacSO7PqrM/kK0qFIWASSGy3jLyzvKH916p6UfGJHYnk9YwtMPG3Ohj3bqcoN0tlLY
VfZwo/1b2YpMHoceN1gP9RUnTg2k2j9rfMasdOD+KLuxyWpPtL0uJ9esr4C2vEYCfc0U+pJ5FV1W
w22HQKDW4uZPLIa+JXVjbLRqI6Sg/FJbssMwX0Hz6OvJIvrq6nS7+L2ltYvbDEwW8OZIUHyxcccd
lcSHxzSEk5VB4OCJjlPdKtuw+NsMU4xayTpf/kug8k2uXFRkHYiLWxhHjQ1IRuX4NRxuPDMoMPHE
GnlIjyavWSmAWr2GSH4ba8XjqBDemq07WbnnC1iVhL64jftvlSjelglYfjjDYq9WrtpYkQ85WELC
stARB0UQrIw3rDkBVy+nuSyWUmv/9q43cdPtIhQymlOwko3qQiehIzkA2ihr3s8cv/Pex3jE9dfa
BmH8nTnP2NQ5IomYPQfKKLm3tgMBCXqZGSuGZKdXcu4+kAtF5wI10/c5o7NQ5gTid56Quu8mxtWo
+XC6a6xzAvoO1cnD6Osm/LKfurpu9F6XmCN1wvPiusjT3eQRaTDLaLBOpZnYq54J0/xK1jFVBMPr
AvQStoLLmndQHbM4uuPgm3Gb2WBGwncmjsncIAIXP2FjDBhehfTNoNlk3e67Nqq8X5fFtzV+Muh6
D974uTbHD8lrbOt/O6ZXfLfAmv/UwFoWAyBM/yhcv+5yifv1Dn3WMDWSl0d6zfx1WRkx+4RzkLC+
T5dJROxvDyI5v8pnHh+gAyC0woCB8+wJmK+ZQg6UG4UfFBVcIa0rrsHlwfaQ1I9WYfrIAl8CWJe4
K/Dk8tLDgGzQ3pPWMwy5disolyYOopmXSZ+/aEbatO1oqgOBNGQCZPS2R2AzdC7LUTDqZJj21Rlb
4Es+/ESx9Hlxp2s1BixDZjyJK3asrdFvBiHS1kHvFRq4V0les8dvhD/ue8SdgM0NktsL0nh5G+Z4
/qy9m492WCSICZIdo1ESA9UaUIbzwpUbNa2G3psZWX54S1rZzFKZq/JA/v49z1cKWqeJOziGZ5dU
veyQvQ4RD6Z0/W6kvTHt3k8ewNZgyyBVnRWazQf/SuGYexIJJ1/DMs3KocxyRauNSgKGCdgzmyqF
UZQp1dQ5xLqPpQ+A4g4R7XKOHGU3S9cXstbo63VQ/dYR+VK/E9OFtO5cNkRaVL3niTmOTJ7sjDZw
CT7bMg6vc7qHsFirVS2aB0+7pmi0eg2rFNMyLzx9JRsw+8sNma4fHBdi3tsTyr5JQSGLvu1j5Fj2
iJRcycAQw3Hzf3R5u3XQrMi3UMRDy12KY2U+GDLXbcy2RIOAB8A+BZwUAqcB95gNOH/3JJsc0BIq
jElp18chhMK4Bu+KmJpIrPZC37vpSRu2VrMlnMf9wk1lm4v6T9WsfuIJnhoUH9fyxkYcfr3pKoQ/
Fgu6P7tv83SLkXsyyfDOQY1BnmJR5jsWMkakBart5vdKbkRyvtJYhuwe6VlYUsxiXOWImLzVbQln
ONXqB8472WVinR5BL0VPjfQ87B9VImklAwFb7Cijq4gVuzKKYTgdLufUHOV/rclE9toaMfDrP2yw
v0xcdgzolmlu7RLa9Kh0dJs2r+InV3cNi+JyLVkbFDGB5qp0xIQTS6VL/DdJKgJmWqLz5KMtkH21
XMVhY/5HHJ+7FC+WYmM6hsX7BQylAwk4O7EVbV7uW2H+BMHrZ/t17Ha4kKxQxoImuzgdB/PAOCMC
+prft31RZTb+ZK62MG/dYn7Jl7UyudnY87BVBSYfpenlxHaW0o7/bHLA+TfPxFmObFhmthA8bxf/
OannFiNYQqa8n7DdjudkFGB8DfnQd6+XDmPdGJPR4G0ktiL01pPa6b4NsvTDk6+KWH3KkLNOYMCA
2oyOIRkr42eSpCBS1XAgaHDO0cu7d+Au7robmaL0ZRu3p9JRH++++zGwgYXXZX3gumSJmLMoXWEr
hz0FLCS3DbA0Kx87Bjfq0JXb7EDrKRe4GPHLV+ck+C+l6xPLVAJVVahynqA49iuZc8ER+Ep0oEEq
bOTy0vAEtBvUn//N0lXTh6HjvE4G94B4IofbIdpySmWYV7fpdAI7Lbd0izEXxYyKI1e/Q/I2imLr
uePpBA+6VR3hR3q725tEa1jEhrKZDzFsuq/+1BMmB5W5qCGEZhMN3M3xKtsP6FYx/VudwpvGLMDg
+G/GWb1bUfw7sNdpskJkpfKbXyoNrJlXc+etXKkr7XuzLQY68rkpWF34RhmJbOHg8PsyPKIKiBcX
LxNcF9TNSyMGvMRXx/36npvT0qgpmmokJ1if7FvkjnCULsBIRDdYdpDOCN4OeCdzHO+7syWmeARG
fWenMOVfHdvu39HNf3mqKC2vSTPx4qV4AWFhIVhbjI0bmmcDsnClcKy1NIZ68WQeqdbEiDq8Rqgd
8enwQ2HcpeUXufc/Sg0+CxgHvm3oh9nqEtLscP3KGQA1PT4jIZGvyye3s/odQ7RJJMYH/DGqElr7
+0NxIuhcIAp6AwGHwx89tOpE/GMM4POwCO41f03RRwCxgnbukqNURdcT0+pT8QrItORVtl52B/aA
1Av9kedT3QTFd2uT8QfP6Bm89+ZHASCOGzLyWiYQ9DPXwwuM5qnqp+yWrVcJOprcluGMwDkq+wXD
7V0Pz1RC3VkVEFdtdyPG+i3NMRWC5VmfiEbSou3hd0ezp/oVcaQMYhq1xJUTQwhW4RKyuaCx3mHV
X0LSgHLgNm4G3ctBrcb+VCUUKfhiEj4wOquVD7FQ2w/lBekmGxegBsjJjoUArwZcyttN5GkHCTNt
qGYAIuTe2dIGOr/SnLrrGUQJ0JTXXWMzjgy3sTnXxS6X6EXRUbvG0HiPzIRtPJ47uGzMl1RIkZsc
cbce5QXwKx4FrTIxZzZzPLDSU8Eo27r57wI091eXZMddyp1/SwZxT+jshvJNvNT1fTl2BGElpmBX
OOOy8JsyeNK8i5PiupMzRrJrVznKpRWX3HHPUqHhcyi0d4GnjI7jJRTC7XRJV2ocN5N+4jG5fNeN
PG4wYefyK25hHZo+SZwGqvRwS7DCWCuO9tbKiZnYSjR/gZcYFusRk0OLdmmZD7IM+goEgsDNW8Mg
IZG5SFgvkBAKUUyr1KCtlT6oTLKCeOcRN/PeW0N9JNApayepbG936rg7hMYQHmWWzfSf/a5fRstX
l6I0JxxrkSDEqCL7jE4Ppu+yL5SgSnkANEo3BvD14sYUwQ3DPqd2cuSzQTBK7UTdVENEspPiDMkH
sG1Tqlgi0XqTQHx0lou6KxcE08OvrAX12GG0D6QHHXzBVurncSkv1cKOFCuhrr4oYN8i0c/I6T11
YDNNR94T5IMqWwnE1v5lQvOhXBJ/GnOcEdJ9Kh76CGa46G23UqfL9PyGQ9/rkil2Y0PYMB+Y36AX
3LelnWJBm/BQ0w024GmxStVktBAaep7UgTYn3uhAhhIX03Rn/GL3HP/B1/OexUaXOQ+PpNbKDYEF
MdkLE0JujC1eaU4TKnfhEsCwsSCU5IthblIF0qIr3747Yom5LyexPpn3OOoEfOFXIYKbeEfPH0i9
vEx8h9Cv+tJhiTNzvtCWAzNn1tCq7cOpRt7PqWEYVRkEhaUPVV7J12jSDNL9XeXJ8mXfbg8hydNV
g+0DOXeetG+sovaOIpQXHnzJMFy01GxKaJY6oCEbysk5P/cRGzD0daM3vxcwfqWNjd/pRH+I8DTd
7RygvY6w1aHzNs5+I+rSG701aRDSV2E6N9oW9KDdhdXzVA5HVDQujFSa4drfMXb9UdiQo7wEvzDU
39SFd0meNzBkGS89uA2RCSfzT/NGWYrsPeypgdLlAF21TUGeaZsjbic2RrvCkTcGiIWnuWw6HHwl
fG+3l0knNVujeJ0zNn2SKFzq7OeUw1SCwoh4lSvRXiA0ALrLCXSSIN59BgjhgZwwiWsth1nk9KYf
tO0yIqvvYv4sYBIBWwp32uh/4ri9pETrE9QzUAxcb/4uS9ym7fDuzHQXJgxFBKzCgtqnurlzry3z
vrkCJQnj47sKZ/PgsJFBP3qHrzkoM5By4XiYXhCFvfLYMZyeZPkZqh2yq47llUT2TomlPZSYwBmQ
DmivLwaGT9V1cMI2jN9ku3QCY9HXrlfBBBwn8YEGtAJ3m1mxXLczgCGlZ6E5fcXvLwfReNJwaG17
LKKxuxt2kWaW9bcy4nL8zasBoxQuFjgH24UOp35BIIc/6QVgsx7VuYKxTai9l9LVCAjjfsgp3Y5L
SDaTewTPJhWzngE6qzSk4IGioFxQeyo2FfioXYJeTMv7r1aXy71yLdAbBkZaTVZ+vcvRgrtSc0t4
pnK2mXiRb+d1vOphNfkclESeX8itBpwiMwYn1/HqO1VGa0UykQkx9rSY4bIKiAIezrXHlSQjqTMP
1kdu4Ody91Sw9m9X5YtsxN0cQIUVsRhAKiTWYkFeD4wbebZqKOD+jgcqs57OcWyyrT/hQ5Zr8Adt
0Qa4c3TuPbJ9YVkTzCBtUDX127PGl4m8VMAOHcQc9r0VPUV9xBm7qWBTZUIEGwcX3lM6x7b9zq9w
qmgXgdb0hv2DQX7Tg624o6m7D3XbJD9OlDkiRvdL9GZfGLFmrsMuk1flyg9lHd7hGNx/6j1vMQZR
GrD/uOU0rrwxy7/4BqCFZEilaCqK4ni8zxrLobBDD6kJiGz0Wt7FYVi7jW9FBLKOdj0/dpd9j8Dh
PgCqbQNhiCF13mpkZVkm5BcKirz3YrMu5tHhJFfgJH4s1bLjdYh1uVv4z1FQ6kxGvT2roQcOwyFH
Elk65QskrsHOi/ywpMpsNGargc91SRv78a4pZL/nkhyDzNjJjjJ0atRSaWpd+rQ33Ye3s2o1oDOL
hNPUZLUsGR4zKVU5Ua5KJ4pRGbEypdvePTgIycAFt2Z+MAJQtnIqe9bBqgSW5J9JtgoZm+/GmVjz
Wm+eXGcrkd71+PlmocMKaMkHvuXBT0uEmwjgw+5U8QUQ4jP+GYJknMPlhxEpfprxQSzX1dMBCH8G
k4BTbiH9rkNHDBLUcPkPQ9bCqAsJfeV9A+CDs7iV2P3Tn9euYGkRPGRBKCa5kJ/M9E+8PU+fqwFL
kO0Y3FBVcGtXQohv+X9D0QPPno2nEcXv7MK8rfhR+pytRWjWNtk5JJOOyLsmENvh9TySsqkq8G0Q
V5iv0lR5j9gqCbmJXNBxoD7G+Da6WFO8+73nLWzPo5qftRRKsvBJYdv/MOq6/botLCnbF+6DuQk1
5H/3QJnwuAJ/fKY7BV6qleyWXT1wkY7gPBHhcoE5KrQBKckMmLLb9A5lCa29VnOnSHWdM4vSP2vn
zXx8BpPvUDip4F9g7oCHpMz2yedHrgYsXDNDkXc3l6eB75o9Weu1oglOVKtYSP5F3PIg5h7AiSuY
uHj5nXjz08/TXxUKz/TPfW4OzIpwypNlQdcIx16tCE9YpckNrXde/vImbkmeL8cozcDr1GuCOqdS
o54hTPN2O4Q/3zxOgCqn7pIh1FXj6W/wLy9yiQDYB5s8GoAmi89rmCYxsxwOS5TpLrdxU5rnAGu1
rmHKKZSaZY1K2PQZbP8pb6j+g9rOXYAuTi+ePl/lyyMQl3JcNk1LikA5HwMJPfKWHsDzeOu9RUYn
lIqLNJI8cLwUH9Q46hF8jEY6oZoFbfpVPot7xtnPWBuCVb5N/F8wWvo2GkhXFDmNIFTARBAbqVn9
WEhKKja7XLvWp4fXeWFD49I6XX411XmxCy07HJNzb28W0EdMs+jgXsDwq5Yj/YMZEZ7yKuaBnpBP
7cl5B74ZZoYDuF0WVJtChxiakZYfo+Q998I9NS20HEkRFnJ0Mgo7fkQDUejV21JRYSxsC2bjR6gU
u+yooRxNVfPNzJqSaOAh7mRS2aPlL6D+rO5AWPkCXJ87RhxYKkdKP9umz1u4bXKLTUgrxLT4J3I5
qGPa9BbboMR6JcQhgSoHXN7lcOEdigeFc7+8tZ3KMF5/WAhPxWTVcROGIfV871IU6DJFJti5TO1h
JoY88bzhfH2sfOWz2HQbbhyXWsLuKskFSHOpxxAK3j6OGpDWrPMuwZSNsyc6xdfyGcyPHUDF3rqb
28eEmxSmpL9FxANsylqhY6vec58FJG+lwsrWspjdUY+B0dfeDeAIQDFWASb/184NMRDAZA/TR5jK
Slpk/YM4zEnowsq+jp5eKgs7uZi+mardP4+k8ZvZ4D9nO/Uo2kPWQYiq+XaVa16M4SrjyuIwS0My
YfqQfyIkJq671cQpgBDQhYdpBXyrKClK13E6dR9mwLlwEbRMFpru8Tz6GzN4pLiA6hxV+kPjjL8s
hQdquPFTO/vH078vgSsVA0xA09xrp46EXlWaUYbwMX1bO/4eZRqna72T8hMT0mNdDwXHQNOrFqEt
4c0DG+PbHBk2Nb2xTzSzbicnalJBnGBFkMBNYA8bu+tmSaXgZyscW7WnUxks0p+deGF158dhPgG8
NhSvuWLNDftNFyJRVAWaVsXtkZm5EKhtOVR6HQHSmKUDh/drym6/+sL6LiuW3FJgjUd+yAbwbwL9
EbYXVMNi0soURvZ6/RqrvyBkHFEcKgBHLGc6fo34Es+SyrQgL8u0uPCcnyEJoEE8QeAyuevwbpFu
GPWjlFU0fH8Qe6pIFitsZ5jO4F5oY9Is845nfoH/9apyM3aNNPcVb3ijQUMHUD/QoZZzLpl/9Nzt
ur7XhYvIrWGcvTtdgckyAoJ5ZitOD8cxxyiQeBXfrqVrzr1j545xt2wjteJYMY19plYQ/eKRXN/q
8760JLoieY6JRJB+FFKDNCARars3NJ9R/WpISnKCHt5ZMPYmhZQKqklvKc7FZWD2+qpC/lYP6yuc
RsalRkfdV/jzjHKnGvijgk+E9f/3ZphC+iZ7A64ds4KW+c1dnBqTsSBxOuJJLn8yhmkznSODuxMB
Q97lsmaIdrKgQ7oBqtWFXJJLlWxBG8sgYn2+ttCzptPMENzLkGej5n2JEC4QLLzh0ysYxlRvWPjZ
cg01Iq1ro17ayTkIS/VeJ/Fh+B/5XFB2ipuKitTzcrO1VjD2vcdSEpvzXJxoWNY8rvGK7LyyL/eA
N7bfUTpB0x0Z5rYcfUMPNrrtHyt2q24aVMAAN0sA8aHfg4R+Zmz4fwm4C2W1Poof9XKGqM2HCYoE
isKY77707+/nneuoZDJ6Tl7jxk4KwyC4266w6z84hu6CWKoQe7PFwVYTXcsNuSxYcG5ou6MyGT9G
yDPUbM36kqMXep1TttA88aCMKAeUipL0wVe7W6Ouw0LY0fZ6dcGb9KQQ3cYp/SFcrJxZekFBSZit
cbaxQ5SIRqSv3weCXSUF0LXb1XOGgNe/MCxBdIugluBoN3gAJxCBIOKdSIrZH7CTqFW4KWXzK4M9
x1xnw57mi6l0OwNPk1Wbc2oneFyvp2e3lOraHTdJOLQn3kVx4KSdhJKQRpcf6lJxI/LSGQisq7AH
28nCx/49vK3TXA8K0eD5IcOBevDw8R66pYt03EN0yUM2xmGuREN10tUld4I/4CjdkDA5xxPiC0Fp
bemme5j+FnkB2C6Vj1oOFpwZtoJhC+LyXtEqOVrliUY0jVuhe5VrsP5vmb7PJSe5XDlRPO9QG9zM
PNwdE3LNU2s8YFcT5/KclwbOGk9970v7m/Uoekx0vrDC7GvxgvTeIoOV5qSipHUd3+17uFHiNqGj
yVklhs0veiWemxWbhFeu4bcx7ha8tKg7lIzU385ZLVVJu+PGFytoCmuJMMvT1pJkGFqyoApsX30f
PqYlVQ1KqXkhn9uP6bPcdkKfv5xh/uYh+nuqgXR2gPqggG5NKrMvGd2HFOjP140s7LmcXsBS1YAQ
uoEQg/NnF+kRIzW17g9qPmkESqKdZGwoSTA0826IMQZU/tzUDd6/9gqGaO6TJdtWerKwZyMAPgAq
wGfrwuzm19V7QLEJ3lBiNYwaiOZbwTrV/p7YKBl3/EoJzHOpH9d1sOCh0yX0VY2FrNw5a6kLxXvl
gKC22J9EhB/efHJXY9XRqleGGbnH8cgQ+SFrEyivrnUo00GhNr8RsNTa3GR123BP7mroRt4Vorm3
HoRu55e8Fg9sM1rz93K9mzBsVsoBBqbOW7WmnLydNZe0AJaZP8WDqutXbL5cn7OT7PPS3BdSMyil
xWXmd4OZVCOzK01K4KldrL/CAoxqbbHicZNDmrhE2GonFloyLJJyOh626vIpq/+c1AWfGQ9X6Jtp
RtH76/wz8uXy1lVA8qyxS/zDnjMB6wqeJz1lJImT2GVWM1a8qO9qO2Jv1SxL4utTK+DC/UnjD6S5
M8YvwXpUCpEFgVwzkveb25AixRHAIp3M0Xz+n1tOs3of+ewn9bTQc7fwQoWt8tTL4X/8xzFzhMNw
ls1/6qJwUQ3yt6ZVgcG21YoJW7Gx58xPO1608a68Zttwq0Dd85jQrTBBh4G+xMR82NiVfd2V2kjA
FVxBnkSMq2WN2u71TS83rYUZpkWh3FhhMSOIdcShr4sYigMJt2XirwHTfEEGl14KVF/n+3GcfX7G
j28APdjG0JPffDRABSICgcytQY24XS9BCX3DjJZNgdizaAG9aloEhhuFqUhSKuxPoMNa3UvNABc2
zqcY57uAXsSdGUT+M2lrcMuShm4xqxSHgvbu8S22zTo3xwJz7UfJI2hpb/uqoPD9GHNW7iEgzZ+L
KSk1vKJPmP4jafngZsm6EJFkK/qt6oXt+1YyB55MNzYs17W9d96mNylUiq5ilLwfYpXrqHxjbb79
M/g4jM/dBH9skdEKzMmHMyk4+/qMHcsSc87uF0dOvQYByAHP1Ah8lYmqbiwh3D1omSgtn3PfXwQp
ophhlyI/DwL2kg0Gf2hS8Ku96tmdcjgcLCzux8jcX2955SCG4e6ea953EO8V4zxrTZX8QF5CAHGE
PWsV5R+a6+55rTor12zFL+4MtNajAsOY1+6hm4+655bi1mVAwFjBjKUZvNrQrKVPMgnObJjCs0Rf
A51rwkLX5XEyetq2yS3T34hHzgQ2IBiYth1UHUpJp10JLRVy6ZMmgW4UqkcZyonHNoKWSXian7xv
68dZGNj4zRtCF7u8NkQOm392vuLGUdYjDE26mbzXLISrpHohRMII1gYT8tXMxowl+zSvHvdrVaE3
5DnGfvPcEozPL6iWoTw+9mtebRyuquz5EymbRiAl+N7EstYosuKfjXKIhQAX+8MA7UHoeJ+fpobT
Cx/JieueGW9/MlOBQfpulhQo3LPnZ4lMLMcs2JBkwS95EERBf920HDM/agUAX25LNYGz63gMMYwo
cb9N+7CNGccUF0MVJmCz6P2aGSsXUNqbz2bOr4FEoASOUax3Hk5Q1UceiMi75fNGq0u7puHkhD1/
XMrqQL3pHMmhNCEOYooaEfl7E6cfhzd6ju4SMNBADhsOvXin0RtiS530DyjEQDqrrYWiBNnLE18k
mKQ3K6ousDng3QBU6uO3nyxqCiIAS8kv4xLz1oKVtwtEdAFUs0CQ4pkNaa04htH5UkiMseqB1JZI
T2BNNM1GKHBUphsnM3MtGKS5oQ2xRR5Lgn1615l/Q7Q1pNv+Pc3VDOI9T04FGo/wQI4bbbX6QTiR
mh6v4pZZhXD3rbI02XP2BCUF92TZBO9CVl5hTUpI9dOJ4s1tnc/0YL01Bg6eDWS8WdGBVB8ZVCwm
0IEUID/OZxGwV76c0m9jBdTJ9ibWITwbTdPEdHaVjzv5bo3YG2iw2RsmWR96ja2tOggQz2wWMyWu
cHw+D+Rl2Yq5ZqATNwST5gnrB3TXNolzQfMmMKX2BPIIML1o9aSXpni2dyxgvbRZURXTetIuehgC
eeVAxdZ02RDSIRqDyFemLSrw8MBDLQoN62QvtHjGljAKu7jgq6tRNs/DFw+hm+Cl8QXtmSc3283j
Sz9IgUKCjuFo6zyWi+oJA00UuIAAQHV0pJbp7y+E2J6Hd67AXcbpzMjtywF0+vFha6lMm6SGf04L
m7vtvZY9ZDKoWC9VSFAMAgYjmutub3IwOc+6TqVJi2D/OHY8EO2aJsbHTXi+ZhC6aGw1ITmY/fTA
5yzQOSj3B8nXLc7QbAnbAcsvkc7hTsMUrS8rWnfx1GrQ/Xf2mVzSo1Kq+QnL/oPDjXEFNgoxWaJQ
kDEu7gxX2SfL79FD/uRqL6wvKRp06pbcw0seK49hAGMiaA1c+3Ed0CBzF3yBCXO7gutbAqAGI57m
mvnNSRJdSn+3BOq2NHODOOMq6tpD0egfpdF5SxdrLXnaf36C3Srr1aL0DbSzpq0n8JsPrszG0xwS
V1fh6pp4pMckWUJHeCQEtyoq1JfddelFd4XnviLUzUharIAB+Gto4ZndbK8pxRYkdXYmQBndQ8RB
1g0FY/BVgxPXu0fcTsKTQW9iTKWLzuH4BLSn4OBl4MIYPAvpXT+Dq6b4Y7zYDR16eNtYbiyLst2G
ZSUBKzRlPMwHSskWYGLMXjtzMRoPwhXAo2jSUHPHoLvNEdIPnicZmoSyFCP0Ea1oSKB64fXICwkY
r14UtmpQqLxfbhLE3tGIbkP2n1pmAJNtLrACAam9ME7iPkvjIryhtx96WZqUid63KyJqg6tpb4uw
4vXd9kE7VnYzT3aQlNqvlpApuG9mn5mlTdKJSgPAvc5+8mVpxJQh/j5NOBuzGxNaS2YzyJRZZRHM
b/tzGff6bhHQkfRaPJvScao8I50CSBkVipMlCT1n/KVyzTpQXXtythm7lN2QZtRQNrHkBBHQQY1H
GVBCWuDTX2jUHXJeVd81QbXphLQ6/6pAwihMgk0PNLLIfST30tiQ2vEG39pnE7P9lRNfzUBm0HpA
ExRJVXMs8+qhFUQ6IhA6F09+jpdoLFoDKyIfaBNmol3q1JOqQLD7rUGyfpmV81Y+6xEB5GKWenmU
krUpw9WAR9+lJm1KXAT2XEgh+j7cTLNdd9HRUCZmh9VSASkqvHJDr7KnGMKf4QwdUVoBZWvoUKrj
KhKhbUA49VF2m9U5KnPwfqm7oxQNfWB/knDzXgah6AXz+7SpVRDnZG1ppKvue6Ch5zC/PCK9J4zN
QG9EayHY9p+oFiJ2zfZlsxQUU/XcqSWikM/MRaJChPKTkwOglE/XV+iBDRT4adbQUAt8t5j6cPoE
asrB1/46u02MNuST3s3BalbbzfDxBtuPyM3o4CrabmGO4Pyn1gAWegWWIzcxHnUKebt0g8p1deK6
QFeeihu5tq+Y1Y3NKxpFDjnbHuWrmWqaM+BQWVnpAgfo9EjIaTNKIRsMzT64aE+aHeQmmP9rSl+u
WrLrzAx4ZEBxSn9W6uF8QMIGx3NMmq/ptpTZvZ1Bz7NhW/HI9d0xZZkJz4Q+5eFdWYOFNz3Xgc84
AMKp3DHovwUtQTd2zMuGDqXriua4ZvduPeWJZOUkdd9bP8KK17jxLiokNzPLvn4Is4ftMw93Y/hf
DQCA5kENwiIuiNyl5Xf7tdIqM15K7Nqx15556xqWKxjBScw7armSF6H3vCygBQS8PZTmtRxT52d7
kcJ04YTcBkLiWcjG1FfAbhwePN0enxfg/mZM9Rrs6JNa3zVpEs8oJlvbYOC4oRUp8WNFsHvccK++
0h8hrvB5EbCUapd0Lr4er6iuK5XyQm6b9s+FPzDhsgkCd/jZMgfKEBZ/e3hzLFFYrPJ3skBdpXhZ
VEVwZr7JCWrA7xdj4cy5knf2Enxf50W/ufnffqhtakEpmhJ1gEBGU7hG0gNTQVduz4wKgBo8Z8ri
OavnUq5TwIVuNEkTQYemC1wFzvzCqdmD9GJRYgMKpe0RLWyG5Zzgist4b0pBHq8kdKqADlTmCQFe
yrmJWmqDbCwcruIl5lGzUIIEFKYSTIto4zGXW9EbthorcUfpJm/igJClAgFyTaAmZNMAE83ENP1F
DsZ9rqnxxJ9CcKj/P81ABCkuc9rPLfTbBWSpPn1e8fMQRDJyvvJ+4saFOrCyKYwy8aNiSh3jro4E
swiPTWQzIyP/quMlVQctDVeu7Se0M8hXwRJ/ppK82IY4NA+8nswCAojJU9HdsnhZtaT8YYKYgqDx
nmZnZ8bup/KTh8rtFi3C3m/g4ufFHABdGvIiwI6+2odA31q468uMZwc+k/t984T4QbCi0dR87HXn
PTeWhJPpF7EzyVx5QfVeHDhMdxaHD8ea2VONbfAFT1vhWy6kfKXYXFCfM4Ju3XY34t919saILzXZ
xFTf3tdUKbCqzSPUcY6VANpbjsoJq7vbrwjjQcIveDEk6wSl3dqtXFkijoTlXB/WQk1fgATLlUZj
EEVZFadhhL9uosJlrLHZL32CRflq7ul2BTCLXlwsmKOTHBmynaQrd+aZFUo6N9+Sxdsp5miPSJcW
3DNWdkHCkEGdYSp9cNfB1WKUH84OymwrnGpsLP0IQE5Ujzp+KzvU4oTOAcZbW+gUsdgqG+1/gvX+
7TGLmI150GY4hekuSms+wN6R+4j/ZfYO13NnG6z+2Ien+FejRgkD8sNkJxAZMS55OyylzzVt0GiX
u/jiJslyOtCHyBeA8mRcMVgeBygt2uOOXOI0m6r7w+Kbrag5OjjqGcE9D3vQ/z2vVCDfJfuYR9H+
l3iaNfkRNzjWzfJbU4wXLwuHVUwKIzrBtFoEYx3h0dIHqOGeqqTkKl9SP67cQUkFbSzVKoYRrX+0
K2a2wNmrCkxFQh/5ozaOwMew2Wfcmqlhp0UXYK3n0ItMuSj6H7DgfzRBWjYH4PPMLPUrrVep51Ii
SNc59OZW1FZNyBJLSWlU4L06M12XwoZQVoYvVm/oq6j/eeXkADgrfFkChatLSHPXFtg0MXO2e4p+
KVrj3o4QVaLpdSo9DI5JrBA+qxaMhg9t2DRz9kslE5zqsUh8P9T76yyQDR7NrR4K+mYFSVUBOYuL
fMev3+JRha7nM8NQjuVIGEFpu64/hk4ooDIG93THclSIAtXOPdiTTXwKOBP3W1Ua0aWvaukfv59V
Cu7FN09OSnlc1oo69l/pSmaGuDddtib+DU6HZaYNb+MKNnSnFei8mje7N/krVkM3Vc2pMwQ4Xnpr
2mKidAdytezTByZNsp2ml/CelmMCskPYyLwME0zHwR4pfqqG6PfONibZjoM0ByZxsxQaBARaciNG
hHpS7C36raM1StYRJwyxRdju94vw04RDnIVx458zapxdGHPCIuZvQ+QBrIDOSx8P/FZyBmUMZQhm
twWbDD5rWafJSrE3l/D0KS02FEEjw79rVsfga7VTPym9/YzpFtUBfsRYpd95ic1zgdeDBZbBRlCZ
1lKyZAD9wPjEwYcDJKgBVFNY0Je01n8mNz5rm2q8lFJRWV9vXAvwYafJmO1mucTMq0iOamEYfJLH
Pw59cuU34M5rhiIMQAAsUCWZdhARjTgITZuB93Z4eHHdqWQllns0Lj8JZ+L5fdDRa7PG6IWRTMz5
rWMAwxsR1evVLZsSHEoV/IM5lTRLfwsAEtlUMXzMgC5c5CgfwF9Ojuvc59fzlkN6FOq7K5uqoaid
ARkpBwUuA6oItaarjEjubmMO7lICO2ZSxuS5mURTqAjRksmgMiAtgBhdl+swX0FyYtH70+ukyMcc
hXrMpd8lIEKgKDjC7QguugqwbLHfIwEZf2uOjWpKVPGBpIuzwqQiws5SxIWbPrDmkXBAZOJ/XJXm
COT2NHvpJ6riUm3nFsMkbNF6mGJhMbpZP45eE02nXxLRYPn4Bik/4oAvMU8R4tlD/xcrcZdID7qL
3ZyVATMuwwbygXuh88nxMiP32c+XLv0uaDdi43gQLlEXe7YsBX11ijayht9CE+QShazpFU/dtbCq
iEN5U72hl17eBH8C+VmfK7+53YvBMjFktz1P2J+qOTJ6SkuBdhHXqgP8ONJFc95RkuXqFkGGPGps
SzGoWLaOkwd9hLG1ih2aQ/7GzWmL70wn0dP1fZLx8lfucUbQiSQKES+KZgbyHaHUxrwy9lw9yBbn
n07mw/874mzkMPWKHYIytE7DzgnPYcvA3nljnm8thb6ISIFN2DzDSPe4cg1aW8LEzH7D7ww88F5l
X/aGekqL+rHP1Dr0LXWMqZ/0I2tzfWAYOER0JWQVWppkjrAP+eI9DyFRqsFHqhkPXzArrwCPNoED
jcY/AwU55xlSRbgTAsh1XKBnJIzuA9q9ULEoRE3ayxKct8co7Zoa8N6Au1o5Xvdon0MrLxIcpHqO
9ZxoKhs3estqW4gUydLkb1ZRBlTENhJdHgmnN/RPRSGTejDwCWXrrz2ypcUks15/pg5bV6HZJmRY
0GBWrSNP1lf//lI59dKftfN5dvryKdxw2El4JTR5gfC0podi3CId96ZRp10eWhzKXdhCrsoDW2tO
V6B5fmDBCLOdUYkAXRXT3+7u+rIposaPHb9w3Zb9XCupfOnE4Bu/Jo8HKHEwDNY0iSjLf6+SnIeZ
hutm3GXJzk5tpmU5tDGjqNzbZx6w8pCaSQPL4WcTiRUt8cYUVKGm/aed42mCIRmj5Nqz+ojy0gnr
x67mDySW9Kp6QszUTdrksBOcmWmArzpx4dEaIniVy/BR1lqPFsGviLEWWBn6DSGb8iME5Kq3wgrG
vgmJKuZugJLeHTToCYJtsP4GTnSBX0eCcerHjgS7d4wfCJ3V82ao8DPcCGI61Xo9jNbUTQSeFXfZ
NRirvPKWoo0p0R0bg/86zUuQQbEjjMkpOAsJ01XfKuqdAGESujFVhIxNkx/Q8UwBsPOvz6qDNLvy
pDJvDOBX++88x9+jf5mufdpSYLpqyHlzGCr8CfP52J10UV/1bo6OxZ9+urGEAXbkgmrUnNAbeDSl
mkywCkCbYrFIxHzsnN5aI0RUVzi2RBRgni+4LvQxXo0WzZrIpKKg9TIMpfSCoXPVsC2RRio5UCYl
0gl8j9q2BEZr1autlL4ZNp3GZAXIkE+cWJpthWPCIdb4DtSp/qNosSsDQVzlBAq25WGKkJ10+4e1
xK4txjE5lAanmspBSoO2RZaTLNj+joj74b91zmcXNVlhGbHXE8QxQO245/+QnNwgrMhJ3qurGF7/
kHJRM0eYARFt4tVwr+TjnZNQnBer5VwhRYCtaWgjwgvdfmz8Ss0QPjdslLkPqbFbxYSBKRCLYVYr
DNNP0PlSIcEMUGJwoalxGpuHFGIRhhjVMC7OIau8UBgBQKNs41mmIrKhWTwFyMojaTrtGRVmKciX
TgrhLVk6IS83cGeA2LBw3C4Ae34D8kRUqFcUI9SCVBeQy72ieQmU5NkqJdEDVQw83xivXSIJ+6aJ
EzfU0tSx8ZWXR8wn8MT1d97j1BOGik4VT+Leh8ex/GRI9YvmHlzO+yHSe1vCIB4+UhxtX9hTSeix
kVMsREHrmBpMEHoZvvorj3Kiep/jID99LKcvLpjq3AJsEjPkuoNhiiYv6Hnlekj53V/KZbEhw+vb
7W/7JnpefrllgosA1h//RSQJUpxAgM6elN6lb9o14rUVC/mGicsRhPSZH7yjb/MT5Kau/hzHO7Z0
+Te54QluDstCfOSFBL9YdokYQK/mqnvYa3k1dbIy9YMwyCqeryd6q2DtfmhHk+aNFfv4PRBy/J0+
5e2KV7+f92PW0rYhdNjm7Z/QYsapLc5oOFIgrOhrBpB38dO2RcaXHFyYR8+YxnZ5rM8kZbnzZxH+
vIMzmoJUY72GLfEHdQD7W7guTdIPF2/B3O1o/98bDl1EcaTUn4/IjTLsi90jvRv6xlqeAe2HIbmW
wHOfKrsBS3TAnRlHKAqWjSdAa8RWo41E/PH2RkKDD19yakLBT7+prPXRKYW22x5lknZVLx+6Y4Up
xsCxYfXeq/V2dvwqux4yCEc0oL0kSY46iC4IWKDZGeWSxUG7m0WDA1+OSuntmmr2fcTcE6HcZaAp
Tr+XGiv+cslp7wMnmgWp6Cb4xtpxLLVCtsgX0BIV4XJ+CjlOUVfX2F44708qafh5omTV0ZOJjcW5
dkOeiRLHuIm9mM1TTKZGGa34Tw3Id4AxSdp4vEY/o17iEpU9wc6fKYchhKrv7lrIV7brJYM+kM2q
Xx9TnLsQtTAJ4nVt7c4McuwTds6QetCiXGcmeZKEnLxdzFbzJM3nk/f0fgxNjogf//3UgyfcLt5b
3FuCfDH/yexKZEUKt/41af/GuL1YvyeZ5+9qtHOZfrhzj+BpMN6+VY3SrOgjIO8m4GhgXPCsCkQN
3/alnDFAJdGLiOvp7d4u7r7c6C6LRVMU7njCe9oQATEaqtz4nf2s7dv/3Nv30k8qIHr6s/9wqEeF
GlTEcUP6WULOh7+TxZas36m355dYlPvl9m1qKSz+tIThALGqSLVTCuwWN8Q75lkzC5ohwNBni9Vp
A/lVTnCZUx6wRcUQAkgYLZE/dhVCB5lfCyDyUVtL6UZdtgS2m5bbw3xOoYPo0838zcVT7qNECMnZ
2dq+BWhB8hMgoR618AxDhPMt7I9fnjSvM5tPlDcowTsY4s0mOj/FhRwGtvR8SSJonbRiUKMP7Frw
Bf5J+/6kIJkeXkwGtNIv0yKG71Skarm2zg3ZoN2lh4JtYHXk6yJhh6m8nV09yP0qMCLZjoCWyMiY
AibRtMEY2oiWllicNZ8RQ6j5YZlJhxdDTPk2kbcaemHA2mqrhfzjMcuE3y2J1LEIza5lXTxbyJY+
sGWnqGWl32DtarMMeCcCMmAGWmRzIt9ADZ/AHTvAWuG0pQ9Og1xOFB7gCEWhsbIpnA+JRjcYDtnq
lQ77UIa7BP0rQEbX734olJWBL5c3CRzn6r2JbXsN21YSu08oQ80PWCxMpHXPF24zyF1Yni+rJ/x0
r9FFiIas4HuJg0g39TtzqiSNA7/tgfG+eePZ2Y3Rqm3UFGNHhuk/9bBdbnW0+IJ62XvOvz+pES3u
lTpItc5FUM+u/U33f4+uJaVy1gsXUtYZ/xSNK9xQw3mGSE4wevnKWS5nDqQSJgr68m6+mTs5i/Nf
yK+VF5w4ySNY53Ivi4bAMvQL5k2zgKIgwrhT5CWeE03DFTyTZdvc9yajxIDV4jL2GjtAs2P98MBy
G4V2+p0uGd9kV044mTehr/LUnwYIPcVl04ifE9j5qtjrIWLumWqbEEqhAHpi7S5b1ie+Xu0BTlfx
T/tvKWM6MJQkYiTitZLZiNm3y2xPgDlTzjmVYwk8EDnA3U2G8f21Ph68dXNb4RbbN2nYO/23OeJB
4wBc40WFYkmpzlr2Zx8bQwLsdhdaKa9JbetWOWSgNu3G8TCjB+yxws++5BhIWABmVi5BWVt88+/v
CLHcKnJbzjguVTubq4QqLmY1AE64pUMMvzgjqeOl6FGbIRmAudvLPo6H83/AN1XpC7CN+KakWqtW
D0udsksrUBJbG2Xl73vSJVXzG8+X5BKM+jcGTV/mEIRSwl6qndVerNlCG6vtZxOExWSjdE5LeKB6
HSPxiFcTC3ZInRaiS9IdP9+p1ZpoBzCXmW2VPyPo2GmyaY0No3N7M3BLDKi2ZepBkncAIzY55EF3
QPMZW+LpLZoPZosto4J2gSTnYYZpo5DWvMGpsNxKEpzLYDt25QptmRPh0/ZgvcdgRdTAGIVsO7s8
Kab0aKC6BHrH0pbXMEBVgyEonpHQKsPDuMc5MjSic3KCe1WafJzGbGRmX/9wKKuKY+Boq+F3ix6g
9rCkPYcYY2dMcKyd2jbYUUfE3p8KM3zFNbph+ZfpEH2VAyRjF2ypETesaEQB8rI31nx9cKIN5FEq
eTFsWhi/OFPfXOj4QyNtvIsbsV9ZzhXw463z9IYYshEDBoCGfWXROrQyzcOjq0LtQRk704q8OxxG
AHzuOOsUPQkt2jJ3OxqS5pXBW2aPBSuFO570TcAGAViyyrvNCBsGp888aE2M0NEYjbMStlOoAo5W
W41VgDcu8cxzltr3rCkj2fv7+L7PvdFq2pUc2Fo4uc/kHr1oSM8krrqXf3N/SS+6H4Y0eV2ejJ+V
YLkAQ3awHYCQrQ/+MQ0rFfDBtfXj0rlYxl1IIMQWeP7Yhioa0sMv2s6JLZLUDNpQqiGuuecarGPT
/nbt5HoXX53QX4dStWa7NEUTCnq8KWR0/EuRrwrAVdiyU6h1RFugNvIdZ5qB9pAtQ98wU/e+G1Pc
HXYBs5mMev7gXW6kjIJvY0IfTauJHsC7vsGjOHxWTGpR86ZRaXORwEGltPvdTyqVr+nO5PrT6Sc9
9h8m5AVuiJSrYVascaAaKmGp7WRGTjTlsowhMO4UzIPLhy2eMR7nGZ1SH8dLyfWqh+keXl+BTnPj
xkTSO23DMeIEXJBD+KMDjxLzXEkywj7yOXntcTBelEyHXliIXbv93CpY/eU6xgrZyJe54O3jlIIz
Bw1q0Y7smvI2rmSEoyN1XHLK3Y4qbKiUFg1v7gUkIYiRXoZQ+aUDcKR0P2ZGCj6U7C4ALm0gKyvj
/4RdUZzmxLlF9+HCti8n9dVSVirsZUp2XKkbRSsh8ETEJFHI1JvalcmiEim93PVa4gAiCUbsHSzg
qvlsco9jI6nYDdE7ZXzxX36VcxGusCfRy5mpHl4ylcuBj0VETx0zr6GZwEPQenO4jRB0GQt5Ztex
AtP3gnn5yBBse0Lw8taN3J4r1NHHG82fddo2RtFPYG4JG/4M+++Xke6Y7FYPvnJUf/pQqy3LX3El
bx0RUtsmTEnCjXPzuKl/tKfF3KMvHB9XGumgVXmEEBSwgBojHCr20L1eB01ptsNYj8NdulsH+CX/
aBTlKc8bz84nsq0Foedg4fqmfx5Vm4lLTupDeNUWPh8PipvSRo3h/HhJP+rzPzvtfGwPcAZtq+Lh
IfKbJ+iDxVkKXRB3duazwXNTIgSMU6X7qecKesPX0sxuTXk8zQTAUIj/1NiDZAjSO6uaMSixcPik
QI0ht2E+wym5FdeUk7BEPf14i+6sSSLOMbDIz6BtBPO3eFmHqXi7m+6x2TpZZ3s9/gYfhM3YZdZJ
xO1sPrTLl4gtMSexro2qNPqUCpOsIRJESFN/yO7KlGVBvF9q5C43mHhHX7nZg7/k1Ru26NBF7LKv
z5MKgzSaqJbPknFKWAy1g/TOJaHHfJX/nDf6K/IVrvlqVAqkPGgh4J6nENcGfyosPEE6auhlblH6
JzRr2nzlrt1uZpzpn95+gO3U34P2UArS2CMNwiU3jblhTfrzoXrBGAnaEREdT62vEGdrMpA1goO4
7tefAD6laWiJF/TCeOQcaAWRWGCs8J9Cv0O1ULPVOPc16pnpsMcae+6nx5thHkt/pyu/bqaOygWU
Od96BVHFpeGc03Cj5sdcNlebfSqKAIRvuf9oC44YG+C1lPigEYGGxziVw0nIjA8kD/dic1ctyCLA
LNdSAC/JN6nEy/fPXF+jMU1Wz9oD+RJ7dTd/THXhXs7kajodoDQ6C29jkGXpUyuoL9qZgOyNxN8q
IZvjUVnt+GI4/DY2eoY+7P8Ri6gFy/9JOz8j9f49YKyaoMOQ+gD3JUsCPuRfBAtBKh/2fPXXoQbN
T9Ry066P/gDv5RKU2VK+wAIhQTCVqeqUCVKnithkdKaW03QXnNkFmsGKWFLOnTLvpriSgOj/PT1X
dpj/9zk72r+u9CFFc4YRri9QtAOzLM7ZW+2GBqQ0msnqAGGPLwFMuN8NxcC+2hiJbnkTrHaWU15a
yPS5PkhoxZazB0nINesRlIwqIzIgfIYWbmINkBPQ6CW6Q89K1a/XZi7vGeCNoN1OHBxzp7OD26ss
QRa/mMF45C/PxHi1Is4jMXrCS6Q/mgb5SRHNUGbX2dKN2cusynRplvtNK7Ko4VeFZbXd6mU+2CYB
WmvsjuLr8U1Mwc8+kmlhp/Z+eCCrfQeGvrCwlJ9DtI6fHjQ9iIewiZL/pUbRgGTOfmb6YJf1PD+H
Tvae8gIuorMkS+dP8lvZ8sCHS4sK2aAZUhOzMfT5jvgsdBj9rB+jmZykBLpC25C4T9yxrppbcz3f
00ZGGfrE/BIx6Y1QxhS250dHnhoVRHNbP/GpTKxONEckBCZ4C0Gf3mv1Amhm+9ZeBLqK/8J+ky6G
U2Wg8uEBGFp5EQWtWnhvaOIrwHTao6afmjEvKImhSq9F2NQgrgU0ilhcB1enIVALVYxonFnNN9Ff
ujZBoW/VRVaAztxQU9/E0MFB7o5R2+Zo54ZLjo+3gLshB++f6DQ3KuvukibK6PPb0HapmJg0LtJg
cIXqXe18ItSYx1r78rBIjpNrVBq/z2vPoWUD1LZS3wUgUMk6xqliG5eDqSc2+N4q8IicAaIfCpOH
t8+QzMJ6Lafs5CTK6miwzrtM/zwtrhsskgQyZ1ZL4cmEkHjMTQ1dTguV9A53y/VqcCm7IFi4B1eR
PFZeOb0jxQG5uY7WPkFpNZ+e0SJdzKupZzAXs99c5qJUdRcqlw8DbbNJG6T8kR4mq1nuBRZjcyfu
e5dGKwVcydBTHYRrLOIny3VYgG6aOfMS8Ec1HWxKzxvhxhcBD11lzdDGyZYF8n3n/2KoZbwc8jHy
jF1TdkIVQr8w+uhOesNn6VBKntHlTZHvt0zwWaelajdjCYP4aKzCZZjQe2T8xSAoufooOfl+YWIA
vYUlTOiLIY0QuL7qsSfalYtGp8enu1LFlHhdSg9c/FYNOJ+kOkCDIGhC7lh/2HX6xCfIVpzvQtqK
T2a+/I015a0B8TbML7ZjeLt4HIAvuoN8WQH7EdbyIOdziUNEycqooBC9oC0l0UBcrvPwVDqFHtUT
OHIBQzZV3y+sHdYUOF5BZ39WcqaQXp+nHjj0QgE7F7aXL8tzaYAPMvAxH15xv5w7PiMsiMtqlTm7
8+o3WUbMdsm1Q5AWWuBwnYHNFPYFpSh8PeBgU3djE2V5hj8+HuUgrZ+c2VNVAhTriidfteNcyFrz
Lj9LV9uNtLPZ23mNVOdp4VU7YKQQwr2ZvwSowexL0mdjMI+0oYaqCt0H/kC3ebqyROaEhcs0X1rU
KQIDeqmSCsqIz43IGrJ9DhNskYblkCOAlYSXcOZcXKzqyx5aDh9rujVtJXLpmjZTilv1jK/7QFx3
m1FfZj7domUQXo09Vl4C0Mtp8uMe3LJ1ellwfNpbhu6iH+4gNpBErq/3wdDnG9iCSH6u9iCkimfQ
lypoyFjLx3G5tiH5G7tOdS2S0txSJSvsozGR+1Q9pEiS/UsDwHRXJsR62mMiSnb0PzegU4nIj1sC
nGgJfv5/evyQ2sc2QCPCR4RvglxGJDy1lkwOWsu4Z4Tnkhg+d9fjf3hMv4KAqgibYi7wcmmDWIIY
MZLG+dDiWA+rjpjsSRjDYfWxJmiDP6MyCW7Q6LnaRF20A75PN70wDXIYBdWENdbJEyV/imbw7A4P
zScLb4J2GNEBuQjzbq9TSTKRJBgN6Pql4q62A8IaOTImhwh9QGbCBpQ3fIcH8w4QXHnnDthm5SR5
QMSq/Z2Bnmmqy2vm0mjhOQpEL807gXvq+PLKB62s7eDNsF6nmNdoMTi3oFVlugyIFf3yOgvKjXNK
b8uQHK9tHEftqiuvNSoGhD+5tj8AWSSYUpx/Uc3iMnb44dE2jQ287kWcW1uq9fQpV46JnQOZjsah
QaBXWC/Adj9+fX+jGRP0Z1+VvJGyP5O2+T+uF83S/OMWagTwwP727i6gdLW2FLdJsAwUuMm1RIRI
2GuBfaURN7EovoEHaew/NYSHf0zvPsYjKt7JzZrbW23ldZTI7qIPlVvolV07YNGNIijXBMIpFw5d
25bO6ZNh2Hr571xqAU1zfOfy3W1b1/XR7Oj81tvXOQIKZTomPvDk1uF98OoYcG1Qt9nWp8p9T8Ia
KRXyH4ZHzRDT4wi41D0S0M9xaQKQ2l2rqFwL9W2TRJJoFLK4aIoPBG9URg5deMigRO4BDCrc76Ry
uMwzAZ8paqVTU/Ve9weBJkP2WzpPQEyEcKr35nUfLIsJAEqDulSWkhQBNH3hMV/6KiNN6qGeOjal
nx6QHqfl6SezUo2uOed4jmTtYXim28RLRhx9sAwlTf4o4j2XHC+StpWQKeCH4B3qDc/p4PPa2Gv8
LP6ARHe+KEk1d2huI5UwfnV3E0wuSYl1eErJEroVQmug9hlp0eGOkKSdxZ9w36puHB5IDWTR8cDg
JZZyX/3T9R4RLX4j867PbmLI3SCiIC+RMti5YCDIrHYCJIZDV/40A86NK/dhk5qZV2VaScvZCxga
rYNfx24dCBa6o2cGRYeCHPdeXNjSRWpECxmRfE9rvBhxe2g4rRUFYyVVvkktNRYh1o5LuhEM3xIm
jgcW6k7TVd0CkyQ/LYMk1LeyAlkMt6wDtIC9td+pJDPw/i2J2N7O2g2fNn2VTUslvHBq7hNCft4T
tbQC+f4waW1t9Y8/X3OLLLDPnvElq4IdPMuCFjQ6jbkuW5jMNPRbNB5HOdRgBKCg8kCPvZYWuTLV
9iM1mGCgp392EihW4YMgWuw8ZK34z+K6DQrzYKC1SnCvQaCwdC0xKd4Q7veZVQIU6eTouACSa54b
eQO9FK6yR4cW/VmHbAszfay8Si1Wsan3SfWQab2EwNasYPK6yT5fNuhJM3Sh0dS4qqiMB/6+HVCg
BMDbixwJRjVuWwJBtABc+UssvOCFXziC/hMSE/HRtNF8Hrv0Qrzy/UotFubK0ldHtoeHtu6Rqisv
B5uaKxzpc6PF/RqYMgaPmezH5v4IIb1e+JPa1lgf646s5LKIOJXsTK8N0I+mhO1MsYtDFu3YiQxH
KB7ExgBtu2JtDcry5ZUN2m2yUWlNqyGAAqd8c3NcHqXgiWgFe4BHJ3d/nlZKQEGXS5FM/MjIMWPl
bCHo+vjS3GUDrdon7RMLZjM6SbPla80kccnmIZ0S16zT0IfnyrAp6DMFR4r/jkHTA+SsW/Ewgkmi
2lQRDBdcj2VCY1EGaEUDhx0KuUAiEXwMY5vTNNWoThYKjHH+C6yPQZ9rHFudnpD98ufJ7G1901o2
OcQNME73P/v7KtVuj/bbYwcDAeHnOiNIq3SZRRv6XzN4KDCrEX3ZfT+hiqhaVM6/z11AxvLKUVEe
b+3wJTMNPm4hdJ5LmCB0X/A59oz99yCoDJhLwVbDi0SyGEWtAdNW4kzgjtL72saKhWWjG91FlWmW
iJLM1BnmGV1C/EwAxLurLIYvCmNYQ3mY0JHXB4eZjA9bdj3/+lABClSiR8Va+dltVsIN1JCFI+9l
dJs8E/gA08JFVAeqQ/Zz5VS8A7HY1YEbLa7QoIDpJ2TmmHYqsUUuM/xKFE28CY1tgqYL50ZOufXc
LpoxvUXmVl7qsFxd7XSokGriqIC0i2QQQ3XYC1DxGfm6CN7UNQaStZVNjqWq49P9kRg5tCZk6f8K
7eF3us9SxXXIdmQ9Wm8fWAkEKoWDNyB5CFEKX4soVj/xjZlroF8MxADyHnQovHFtjZMBav5lEpk/
DvYHXEJwdk+UGXWMSEXJy+6UknOKNPj9prFyKuzZQ/nvrNoygTeqD35OJKycILMffDuGe9o7ABBK
ZsTAFD7LgmPePtYyVt7PQ0qbAi5/eIfPkJuSqmraewHmFjzht9b4O8KwzHKkpXvmcYdYQV7Gixqj
TihFhz9JxsKG3EucrST5noHU9wxQ5Ja+hOLVxzpYaNQsSN4TM8u0BuXov8iUXBo+kLHW3lCXxeFg
2E4nyHW0SSLZnPNU3r6H8GKl0HjcD7ff13t0IZzAvMN6va0khiQIdH04EB0JJfbyMilqCJRUzTad
zfMocv9KQyKnNe9K/pSfq4UV661hgYxGCRi81fdRjsLn5ARjTe/WPVX2prjhQoUVwU7KUu58xNPZ
O+nPZbXfObyN0d1G1G+Dai6nbGIhUldJmTx8a+bOhMn5uBB8ESUd5Qu22oLHS01T4u1KuA6knWpv
WjmT4a2MCB70HGISwRrcoEb+nng990tKukk4YkkOGPLnnmVSkQ+M+IaHFzP48POZ+nT1dEvkhN0W
EyvUnYDcNfEKUG5fOMRCHmEhtjzX3R8y1wPhqW6w2p/JyXOdr8TQsXbJaS8DppeK1sW/+5/SvMXI
sU9xv+U09hE5ZYoL4uKL5gJ9bSnLnShyWc5DggRkKHi6qs7YBNNy0DR/kH+G6oP5AjHBSGk5tvAa
GSxJ3l84obJSuHXyq32B2ZnmyxmCZNjW1Y9cF0MDKgnmgVPhfzeMnYgTrug1g+VC5W/5UzeqWyYg
qLMh9vLoOVQBxv/sY6i2vNWpICptnUYp7hu5AqUGELY1oCOwtkbrK++p+Seqx8+URCidpk/eIg6k
OoHkbdtpXkmhoeFqndtZ0yteEVHWKLIZweaTfNkZro4EpL8JJx7bTVvlWVMDhIxwvHA7b9BwTy4I
ofBiJmadBGh7ioyRZya/BpdRwLhFV97kCHlGA+blkuBjt6WNC7HVqNLVSiE5x9AfWl/JEkbDnXX1
rZuQjXMFRrvN1f6Te0+Ij0fizzGjDGaaE2UFysVVwRwgmPnMM0BVx2vewxqtoWw3OyZ4QRilDMhd
it1tgb/f4nTvQpjxSlbF4dw4vVBm7KQbzSyu9aB8dMTewqZe0WKOE5W/LTiTvyBu8Z3mchFUCahW
KSwXfYI8Wz/k4VnsJwfpUpIMXf8f4Hg9T6qjIKawZvZtqa/S3EtjwfzEoMl8iCFjD51eeNOwC8Kf
hvLDkCMCRERr7NryZ20kCuqP+gvnoCaX6WK6Owotp0T5CWl6KJPXG8EJFOnSdo/ukSDcB6P+zR2b
Wj2/TCy/qUdlaYzUp8T5Ohxy8koaJxVfxYQEOC8h4AXqJihFI28lc7XmWfR4f7xdYWW8EZiqcrfd
SPVU5Pi08AjF0oT0udL5MxnaouTAffwpkyQ+O7Q7r3Gf2Tvxy/nIe5uAYIp0Ua4PW6y+/oGijhlk
s3tsLxu5Jyc9Gc+g2v0e3wnUmo3WbTQeFawoOY+VGMqLpondvMWlaGDilld8f+GcpyphK7FCkjGR
MAvJ8iOzp2cF05Z4uuFOB5k1XnryEmIsydhKPxPR+cDhJ90X6leiWDfssiPf9qE4Ezg9Codzifq1
4jJNa/B6k6RjGfP4gABZsqiYP8sUHOwfB5BHW2RLENtHxSSYONcMs6i8bt0v5b+xaL8DE51Ngof0
gdKkFsn4xF+Njjbupq7h971iAQ8T+UP7fgTuZURt5jlPpjwfLpEphyqo5/0UriphWOOXosIvk/A6
/k98gE7igTSp6vaOauj/5LVZG7ZlGZnimk24lylImpdUY2D/VBFwiE5HfwipmAUMXmx8LZ0eH4tY
IRmopodaJWBy8c8sbdIYshbJsnmZfyKVoUt5pr8nknek0Iz/d9RJvhMDTvRRewXyhveznzKxU4iF
JG8FbMCZv6qVaVcI28I/Domyy06m2Nkbk2MYPAsdaM6HA3sD6o7QMINQ160CCOLARPkWlxA4kTIJ
YnEEYsn0KESP42dhrKpO6f6+ybDRLx0S4ZiG0M1duxAXrWfeELbtYNoJRBLyn1oTLW4NLwaSDNTD
C9WGTZBP8X6+ibuNSp6/0VEtRxa5uMbYk7+8c3mLPXBDt4rV6HlmwnH84eOl26aKDdtgIP51E8Ax
xHOuHwx/o+IUWtfDXIxzagRZrzJA2oegelN0cMkPw2eoiCZll3BuieuSXSPPBnFAtW1eJ20LdO0S
1T09MUkCHrEJUCPPjFFNUpeOHK9A1SBdEmyAHnCoV7kVscF49M57b8VXwjcRkf7821XwKrsp6iw9
u2Or3Yt72ARjK4QedrQMG4451yXLb4lyJHgXK4o9VLr4OzPabm3AACv/OWoeetyl67lfaMSoGVTD
4MGI/Ps/gTlbvrIWAtoNvaZiZXmbQ/JqUVLMzOJHoVB1/ECYaT180jPThSkWAJaEoJaVym3SDKCq
ei8vqGRN8cEMw8XtMeO63AsMRjVWRrHx/Uei5HuhJHTbyuZQyrvs52iNuHhmvkKI4c64+2qxRl3W
zX6V/oS5U9pg7Tvxk/x+rq+0Agw7TCFaFg6ZxHMMB7jDksoBxFgDyb0DRyr2xTdsjvGBaxYKnfrG
FgTjy6r0co2o0xMWSCTW3++Qd2hEUtpObkXrY6tRdQasfHxYDs2/rRyP6KYAHOW+Fl/pChzFD4BR
OGxYE1ZsdoRMRIO9EScc6Xm2adK9jZt1eKMUuYFlaIW01b4Jfqo8FoA+Fj9FV8cAhSi1+VkEuKPv
sIkURADySBgmgLWXpB132XtxMYOyU6Rgytm5Y3ZtThlF3Rm+imZyMC5BGdJEPz4wODu5/YqlO4R3
P5sJEPcNCDkegvi6PxGPx3n8dd+z0kb2siQ3SVrml89neEBlw4kewgMWS78npY3Dg5hdCszk8JrY
Yi3Xf0iCUAg1LFAIuC1w5J2zvzE96EOs00o+u4QWdukts14s/W0wZMCjO0C/483pIFhpiIti6tW6
Vl7JEr1annmfaA0ar9/BD3CJ5harJ3lmelQje9ZJHv/KMcigJay6ImrEgRQkfdzA7xoAE9gtKkw+
d21nvmkpR7ItWmjCfKpS97rnjjLWBTKqNRPckJQN0l87FBr1v8wBnUUXNbKLbML9PLj48ztnSHzv
zNimcZUV1i+XxdA7NbyKf0L/K8+CeBmLbeyuYnWmkCtFKDYuSCWDUbbt/jQQnEQ7G0OSkPGe30dq
buz1OMalOVrPBFoDjsaXKX5M29bVcWZO2Pq364i8l3f7J3vJ5hs3lVN4pZOb4Cxu4lckuF2XsZEy
IM+mBIVIwx0tFX5pR09z2gODTCeEOp5ktgjrKXR0gYpdgNhfSc6/93x85FtG+YT0nItpral3Jt9s
94d5MsoFvUwyjBYS4jQzOM4PIsLu34HTfk/LSP2u9IzES5aw7YHUzxDcP/QgqmTL4fBOJiE36M+q
Q3p+SIe+B+LMUpsAQzUHrMmzI0+9eMldIlk0xAhP7sC6WZp4pqrhzb1Dn2rMJgmfjU9LZmOQ9Y7x
BQ5VKB8c958WXBfKr6J3xlk8PzdYAZwvbTNRebUfgYF0jA9Q8fNHePueEyEhp1XGHHQ5409ktIhq
40FrB6GVPs7nkV3hDsZ1OsL0TNWXMmO/Kpb5dRzUV8A7fBD1C6VjrTC0+uZyytAAhpCUhOHRxV3N
B1CThkRny59aIi9dE13NenaztZqm5cJUNqe6L+ys/CDKUv53zo1DmwDYso8cpWwVj3jHEpnQgeej
ICze3KttV+7PopwBpLrfaagspp8+MbtdaIwd84yheDWjX3u0F/ssHRtUWiY49FfEDPwZQwtKkS8L
xEMsIvTewJmtxQxMiyE+UNui4wEy/eD0SKTrgM2sWKGCuY5qlcx0Ga8a4D+uuxvCviT/CKlWQtc9
WvtFJJGjcdmz+2PNdf7gyI+mOrHSdKH+91XLpizh1pz7Cbx1LPUOo5ITSF5ODEtqs4kRx21kq/VV
0JbinzNqdaAr5TNaadnwzKiljUvRq7oS/F8z+W0Aja2bYvA+vKnexhfmdS/IO7EJ6ebVZAR+7NEn
7JCLsV3fU3ccGvPSkQuZmTe5ZWjviSKRLgWLowFerGfKykw+bvgx5z2OnsskJtXAnMgGxqreNo+U
Ls21PO4eAPA6rAcFFa+szLbKL3Ewcr8ieKDXTBrTDUanA82ZhuW2LbuIrRnyq2xhuSgT6WkAVV8w
nze1cFaiNqe/MjHzlf8WTDcd0Y1L843ZnbDf8H1bf6ztSOQcIVUAyiRmOLr6D9qBYnDs4JOQeuIV
Tk1YvdnIwcpH4aUpqK28WLAzB0gKvp2MVOlXYyk1HKfaqN//pVoEWkcB4WdBNsv3YKMgvAKLlM5H
hL72V2pMkcKJuZYFso3F0oI7QSIpCpluUTCOp1G3KTyDOpE+y46YDpnHWjPqDvrEOUzEq2krba4n
ILVALXRGLINz2vPUMzM0sBUcAb3PGRMCkwK50YyGhvSJQs1VzI67/2tXM+BlCB1tnCfl5ZVNJYTH
2erLvu3eFTmJxEH0DoPPnAKxyMKvR+yqQtne17dfVHhkmAurGEfRs69MHkD6YLnDU5SS4JIEmAc0
oF8S6OFz3D0DH4YtW14sArviqoHC74x2sJcpfFCjky4yznnLjhDKwliWBNx2HRDGKXc49a9eJ0gS
WGgLWMjaE/oIkm30fIIxrknrSLh2fsIoDZ69Me7WIHI7fxNE+/oV5a6+8L/7X0vBtKBuBxdHANZg
ZiKxNwFwrY+LFu5MHNYk1PF+qmQqtyUubWKGdXjI8p0ZWmVhiz61eHM/p9q1T7ip38/DaxAb1IFr
Rpfhg/beyDJESJ4urQLDIYfS65+Zkc8xxXrcJYqi5Hj05HR1PaHanUnz3WMwXRkbenLaJ7hmDJxq
cktIRraQukeup3SvHfLiS8juaGFJBjmA+6RnP4VLxg1rOGoo+PJqjpOKG80pYv6m95RHlKf0enKM
Fenul2nxJ32frV7UvnugO2QpKYACjCd8TgjB2Cl1TDCVrYUflJ8WZE0z5G/0sjyOr52v5OpVQNU8
jX9RU+80JgKANuNrfmDhOQk/q/nO6ZiUSCWSSSMtmj9IlR25ZKfw05oGjbVcfHM81gx2SDgo/g69
aNekXuM57RKxHVLQTCMobMzmHpk9T+FjbZTtvgxYyD/OyrOtfo7QkQwS0vswfN5yupk2a5ChyZWY
u5vTgxkki481Gyr4j9N/a5SZMJFVUfaArCCqiWWzvyMCuvpf0mJEhAOdw7jQQkfVs93S12Lf2Snl
XOCY3mekebDaawwZ1FPcb1+/mYpSQIX8hK4TIJZoz3MlSoS10oxE8GcF7nQT5k3heFsUS9vXsG9q
ipPOI2bR0tRs1SPp2xcaBVfl4HKDaYT72/WDIUqSDr04CZs/eXbAfdbPjiWhuEEcLWASSXEInSFP
CTJ/oXoO8CawqVhxzyvDy6UDGhn6gQRvnNlxftskLcwKWrUOni1PLN5/nbglV8LZXwux/P4T+Rr4
uyFZCriEFdSUNmrM8vpD2rZW46p7F0f4DamD6y9mFcm2vawSGNkTJzzkqv2e1egRCZEoaZ2Bwtpu
CBkEV3xmeSo+K3AW6209yAjW7p7rfMcf8N7XEBBf/MKo257qvFCEssndIZrhHscUyrYCKnGrS2GM
J24PRFcFwfvUqAsjXfnkjnGogY3avt4TCv9hJgvjErJJ5vkRyTPAJNW8YQs9pjVsFvLJYG9LODWg
pdnaVSQwxKLP/xa/aprlk7Fcc8mvrXsEWJyd53W8pqOX0WKajAg4trBiH6u+X/RyZYWBY8YWOa/N
ewfVi5UMzarDr/YLSWh3f7iuR7VMsmOzCJiJQsOtrQLGxegVULMatYFa95lAXsUJl1yHFBChlOH4
sWqUfJfx3ZcyRGXolzWDDStT43sLUCHAQyVVBYaPequSfdFvfZwOyrw7Py8lsRQNNZtwSJXBqybW
ftATNOwrkj1BOf9XFmPOJXGH4P+IFMIL1lRe59sGVXpfEpOXYIJgnyD4OjgHv4kTmJmVbuhEND9A
ykbO5oU0iqf74trcJnLfahQEoU04MUFU5i4yRVFvf+d2+I2lDCEE+AO49oLKlNpp7xVwrIPIdfcR
O1RnGu8vm9CdenArKPds0NdJ0wEacPqKXJ5ASRR5j+dKlpM+WaDgBmOGzV763blR2H0Y+5++xWI5
BRi4Z4WZ31B+3DtxW7fIXrADqGidFHDQfhdDlQKS3K5Q7PIY/N9UFwavujVXpZ1io1hOpDJ6A7s7
MXv/IHGBoQw39wCOyYtgA2tvI/oyW9BMp5ZxGlkykLu/8QMkxCg/sCg6oXXWPS9Sy9ONRBseSO/D
1I4le29w3lquo/LYWiLEur1cuLTp7Y0tKsZZMi/CSvhX4yRTyvNtpKPtUFkORQM5SOF7eH/PRcWG
fx3y+GMnJCJm74cC04epNvtziiHaPpLHvJcngOCEcxAZ6aikof1LkU9h5a9z+s0yPkQkGjFq3rsQ
iUpWkzqOEMSxVPvGawOnkL82V+OHtIqY/3w4LCnvv+URpymDiDFSReH8y7FqBqY9sXCpPpQMY7i4
ve43Xub/yydnXybGpoKG4Xw6feiBxBQCBWx7ECV7hqZ+GNpPmKCjk/i62jEzgVPTqZQ+ck4fQURQ
7tj3t2hVGSUyKicnAPKDbRhnAKMGPrw35E/thhEGQSafmJV4HDX5o5xebTWVJb385pI6AjZhuiGw
4szQBPc6bFWyIfUC8Z5GIXLzl/1UzAWz+ClXwxpYwZTz2hpdgZIAyDoT38fVx8s11QsYVxgAPPkn
oN04QMLb/hTHAcwm8HoxKtD785++LZLK46BA+EHx4Ygxcrkr5dDDYR97kojmwpfOAz7HrNBoWs50
+sGhQ9F44J57EXk4QFluKvPgoHP0jTk4qUW1FcwwRL7msEdZvMWjhLKWmvMAK3O9EKf8TdUXcI3B
7aqX0A7WTbR+s+zB29KAOi35tAORYmnU34Q15cODkvkSKN6/gobh8CE/IOw7I8pPWPuq2xnZEL23
kWb7cQVSU78ejk/evAuLsbAI5zPXd/nX4hNx7hvwGfPe8gCy9miAkjImOVJoL1YpOMgT4F/uiSLV
YwB9SVoJH9FQC+ZxsP/l0cJIIn/+j9mzhlRpyY8FmsQIA6rj22qwCTHZRLSus9jJ6Bo44Nt4cSqP
IcgvW/UVrTsew882OpOTxahVlkG3jCEF0tCvMqUqcC9zOnUOzfAwEp8JdqEe2g4ZSyEZjvJ0W5RN
d+dfchADTUpIlWf9uKKKLY29cvltIqSYDoKOLZzlTFWN2lSaPowdkw0VXMKuu4EOYYtuPFXjqLZX
HzEcySVkjBBnwy+Nbky3aJO4zW3OFZFyIRuXiIO/IdCwAEK2nJ7CWMpx2TVIzBE65jjsryV/QCvJ
QkBlx5eGBxICBjcPXiawcuVOZkMFzmKcBgkxEMAxcocqjirmkWcJCM7732KsWVOrfRdawX9Rf0pE
vkciRcX23XYmXeQNRXdlVFjlGwA4p92+FlzpVDWUSsif59LC2EUpssLkiPpUwGGr2gtl6nnNMhiT
QnN90hzdBlTylwl/OPFF8rgetZVh6GhPpivO/2gj8ylCRQCg7vCqGQ4avLeAKB0KMWhC/Y4mFesC
D9UenlFhTNnxbSESDmViBsQ6rWlvrjQgJgB7dyMibTjm2171Qh1oqe0GrY93k5URANxZR4BPwMWv
zbc4LicxQ4a6Y7+/N4ejSwn4rAQOh13y0YVQdsACi0KxHNj9fYJTV+q6BZZbXJIxKpN4ZdC1VCxV
SljlYzSj/gXETgkUY6hm3dbCGMTM8QS0s9OyEyxsPhuFF4tvTQRA9oY/+H3HhJHzIHrAscCBCqzU
CPGOYaBaZJmHues8f0g6Uc0g2U3mhYJ++Ji3KGqvpVRnumiv5uoj11/KLQbfJHQMxXWOS8z/xQxG
dpd8s33x71tRIfPQRyHGUw5bBzfz5FXXFZdqErgMEQwe+1S/dVm7XWRI9NwzzG8CR7cjBrvPj2ZM
vI8S+zcAlM3NssQFiM1ejsFox3I/gMtOSKdrGGsib6e4E4JYQH6IE/JoMqmZgLjfsSNwouVuQ9OK
bWIF/4F1dVz6VUGVpYSODrGaWR3aYoSR/4W+xK3DW7I8woEMGiZzvTWyy3z49AyKlunJxLNE7nYd
Qp1/M90heW8se/SyqHZdL2N2LUVK5DTGHKon5Fn7PIxa/JAFYos+q6zsbmuUWBKgaR0j/dgsMzYy
wVPhzrE5pxpwks4Yl0LlNMuQe93gxfYQN152/cth0OxwebAg/KXzp8/1gidsN/kzVesXYTyZb/5q
rUzhSmzol9PoE6sn8XkXK8lnnE9D10xMo3Z/YCzTvj8ZO5dHGyUuX6bqXZRUBaOE8yZCLT6U++Gi
+xK0YoN3wrkg03dVXtftWmL9x2rumCo8AU3Afg2AdThTMpbmXXCbnWVjh7d5/Ab3BW9GiP7C6wao
bSB6HN8CHarWWPIvlyGo8AEwhfzu+grMC65X0wB89rWsMpyKF8L74vMPw5BIpHxIJjc8O9GsnTNM
DAvB4nacSd75pLhz9RBiKp1L+rOfAhcAHqSdsvoC2ruhZof+ChzEhiV6r36PRHXa9qYXu+R4XuKr
zyTs4lV0zP6hFOqHoPyGBSQi/D4o1JBWI6LeRK1hGG83ZspE3aledWZpLcl7kG99q+R2+YpkFME6
Q1rkzYvQ8OYlOAm5+cZ0m/1VqsuzMqeUQQaDF9Up6npX8qHR36OR4HZRXDmeJUdmcy/oNzFF797V
/jHgvb1YHnGsxt/780peJZ5WmolkFxt2DieoD7LKFaRgbuh2mLM8g9cSo/tN0MLEnefP8Ypll7iy
AhBR6LttrSojqFwvSVR42LjnPOmgBUUhwyqXVGtgHuNw7EXGJ4ST207y9Us/pRQ14cQZfWl2Nd3G
poVPVRBHdjdPR0/1IfSiNneHlfyRdMelMbOGT5feaiKq47LLGbJHpKFgZubD0h3ZEu9DHaAyqQZM
kYd+Q/vt/doXNFG1WiDF2avjYjTybYb1a0CjwezyuxIVUYotCvNcYUITx8XVONuhPJYPdkgioWpE
LYxnJ6Bdd+NnTeoTAYSwALtgsqJ+0sxyVx/zoUi7aj8f4Scy1sGf1ctMweK7jMbpMpMkuYEnYgFv
SssnhL8m64Fy/xf+3YPPYqz/cuAGUIpbCLuOIKyChN9whx37WwhoKMtYiPXaMGNCF5XQXZuyVvUV
M8wlkjLRrw2fA9k9hvNePuUVYX3X/U3wWQgFYfOGc7c+yI4Mr6wP+FcLVMc/jGYAGKxnEjKkQbDE
CbbkFM+s3fRnP0yCbBG4IvHOsM/dgLROfhn1h1wO3i3pXZgnrOslc9KxwfIcc9SiIPrDhhKN8Vh/
WtuxBlOOkkawz1GG+hVuKuu8mJYS2vy5lTvuJMQwLRCh46wDSppcxZ+wbMRppdFLjHjye6O2QFdY
FkhtvC+v3UXv9qmVSXeUglwzLfilO6s4Otv2L7CWYJgw3zdR8uLw/USD08WEMqw8a9QhLuV9DCDu
9dNK0WO5BO4f+8qU/MyesTcdRcz6fuEUVVXrfOoSudt3EjEOz3pMVee3LdQKYPpRCH4AWBJcLY64
8cFXrxRJkzPjlSnHTCSkhOHN586+XDsnEqO/udsiKqDd28wmZH7QvCgNVi8A9LuBiWnZj/WOmNYR
/ej2vbc6rVxFv9jLYdnykiPPUAWL+Z5w9CmqzTwBiifY72cLxX8yf0FQeM9oqNcNwMq9tOGNAaol
Qrz2meJY4NVhBsbuHCR/dU6jygk7wi2QDj1xQGLxvItFxQIZP9kTR4DbXxCD1pkia6PFkFHusgPl
TFq9eqDTfMigxHlVnSTxnPAr9ur3c5qjgg5ij4SkABgTT3kqE3ORR/QzzvWzZQ6nWXQcBYVU+PtB
LKUpXPSzNsSSnEJNH54+hYlWoL0BodUNEVSvqdNvXn2XYhzqYpHvRDeItTT8qH+NzoLLzNrsL1Mk
3nr/nYqp/eEhjfYY5qX8O/K1igEfzMm7MXrPMrIR+80zHq47zyUZvR50E4hYbF32WgbuiTRSxjSx
Myh643qAEEW9nfafQG7KMT1Lm0qTqlqKvRYGInV9wW8c7loSiWmCKHzLIZaqM8vWevAM2It5gslN
rfUKwud9KxPa8jcEhFV6ZLYohXzyeDgI2rSel7q0PbxhjBbNyg6dk+KFtD8k5Z3umRz0/kkVUPuO
oCWQwkYnoGNmIQ66173+82Z1yPBds3gb3y3xRpe6sXfU6URsYUg8iIPZ0M/uXBoju5MHFu69E6e4
ydkVER8HIo1D6hT3r2NEEoXDflvoRypcsk4x/NTk3i3c1kp3hOM/FwwkIHPlPu1V2Bm+5E3uK2HY
RaCwHO+r9d5yCOdwy6vj0cPqvKGhMIW/8gypGOZ6TAa3URwWg1/rx5/leUz1cHd1f6pjt8jHan59
JZd0w8nlA89H3sDCi61z7pNLXYUb+XTYbJi4nsMkp7wsCujnviMt34FW9ambU59/f7P/8X1/wXn2
v3hUpBdE+cQ9VR22BmEvKUIJziNg8EA4ODM5Y7wlJnvsuaM0m4gXSYf6ug+DYJTsh35lIv2u1Kwl
snHaIVaL1yyM2UudT/UwoVKdBmawG6/fc9EKrbznbFGjyIJZ5uMtLLy85YJp7mC6TXWBYkAcO6hC
Nmr+Kaf6mZs8NCywZJF84VjDcmYVS4a3q32ObliFPQ9c3lo6W981GgaBiSbVo+IkxQutQthS00aF
SWGsTI4E9B9gENo+mBCYKLQCaJm0U44Z141VaBslMRe/YrP9+6Dic+rk4sWS4M3BpY4m5i4IkO5g
lnjNtYlBvGd9qDP+ZfEq+eO+Xpv/v7LIP2DiuOSRc7Ujw86OdFGl4Kbgbzj8ndS97JJ2bA1rVEvt
38dAkRhzEHih0+63Bbppm5e7WDq/6PV6MKp1nfCTy7khjRvi1CpaA/zuBkEY4J3ZBGHUHyxNZx0o
vI5Fz8Zeo/qgHVnEeaHfUrBPeyVHSaxquAH6vXswCBJOZSEYir42SL4bC7JIqVA+qbDtrux13ajO
5s/q7A5+6pZvlPswOY1fmo1aS3ABiY0TDgKUUrx3t70UfECB0oG5P9Lv4HG4Ntt2YJ7FqX5Ns8xd
rHkj6DMfVTi2Kuua6Uj4Y1qhtWfqvElG0rSKpWQCbvoJXEvPaSIi6PZyrqVaj+8PIpoRtXmHfN4M
iLw8Ms2hwHJMzg2ZRgH50mKHvFTc3qohsBfvY9XFku9tZhzcoIncCyLQM1VX1Jg38L7HVRBdz85p
6WI4qO3p3UwTU1TIlNfpwvSwwA8O9kmijeImz2DQB3UoMEdSbnfGHHrz66IRRWid3EaZ7j9umkG1
LecFJ+evAPMFrvR+cFeDEo0oMZ/APBfmf4GEUufHfUCHYbK5aRdxwz5FvJ65AJmfwFP2AVL16XW+
vf7Z63/t7t81u7OnkdJnGGI52RR8+dWrb6y2PEQce8etdVlGDgLF5AFkZUjUZgEYvXdRpTREgykJ
rdAusiJCd3Bx3fpSo1Dr2rzIb+kBxsk9HHRCkBXJJAliezwfyqEkbSX+sxayTjDTLuomLGfQ3FGp
XtIrbLfqrAAJdJbdR1SO343g/QCLLOTjoUm25M1nrgUa5HhBCW0viGAoec6Cyh3SkYg/fGyKfWMN
+oni2oKaYE/AVlQfYToVXBVCRBcGgi78SD6JkTqlHtMURUVlPsSpr4CyjxL1pa/OMqhruf+cybXV
IlJ5AYXaWSMQoaw2GWAxVcW0VpwR9ADP74JTvU3PHGkH3qsb1y21c8mSFBVzs911D/k/00ZiELsd
08nw1vzEE80d0eePELDtvY3t1G+4BL8Hc3UWDXo8I4/9z1PdkawdFB/c48n2OiYFGEKHLymXTJns
aHZW2U2GyW3pfxo1vRftXPrceI72Xaf1nPWAtryCRTHyIelWqWWearrcl62PjZQ4uCAIzMCATgA7
TtkyPmU1LxGLqED6j/X7VAWXsOxATW3zkZylMDyTuBW1RcfxfaiWpg/t/vw92KMbXe7HYU7M3kkU
w5/4JLl/IB1Td1+mdwHNGn013hRdVWXbyltkbybiOJgcrGAdLwc1kCLX7qtXZN2EBxqi9sMV2YxW
8x9CiyVWpwGOWA/+mRSXA3kbd6Ury0FWxtKvyqQ2DisrhhX1jstQdLiuVLqDnlNbMrfXCvjsYQKB
oFhkfg4MtCAycn7fbhTbf6reMC48HoJS0PScbos6ds8ZfCyD81+UcBU6K/UabiU1/T+NoshznjNB
Q2/ErJ/SrRgqtuojflS4apxBCEaasO5VNJ8BtHGq/SmyKp1Ep2swDGeotRevKySKI9onGqQvANy0
CXVKxdCE1caRhNGmwCmUdZm981U//9rCnxHoSJpzWN5tNConoFtiFFZ15etNM+G/XL0P1KE1SzDu
2rHmE/Yd2yKLrD9gUI6aoMG0o6dxtDW7d87hJ3Zm3jphkB+n57JuUr2C/u6bbPFAVAi0jNSCJoCV
3EojiTZSLp1csUb5m302NST6ufkoP945Iul1oBe/H+xmO5XG8AwkmhuUyFjvnIu+DWms/rNGpSIc
XQ55iQdKessuGwUIfANmYCGnaeub7qDy94iuqI/UN6bpR7D/440gJgW2lo2sZ4tyZFvnKtDGJtBD
CyYugIfq838wnHmBjf/3XUWyWAIvQtBWG/tz6IcDwzl2wiPQeT9rr/yJJjjZmoi68k6MVN8s6nED
ZVxGS26u3UjuYaOhpxRgeZeGTYMHJc5c6EGm+kx4Wkpin3HMtNk5pDd+RoxzTTpBWk0yDRKyyurT
0zoAihziNrgLuiOzS0n5QbMul2WCY+MJSXUIxoyCchvX26SSemAau1JNkOY2Up/5RWf0Gr75mG+0
gzLQ4g/J18o9TsXyrewL3mZpb3yu697rREjPr5vlnje6UeS5RTjU3Sv/17D39J7RyhPRXnreaKR2
kmkEiuvNIPOe+MHqHbSZt6hJ0s/VLmR77owlON4o4DtgCsHnxK5SmPDgqCyUjhYzU9yA/iTINLff
ZYzMGvsGPwSC6yuzPkHexfIAnlMXZoN6m2kT+EjNSd6H5rsWmH2apiJxv+h7edj+I+3TE6nzkJ/x
+uLx7Vf4NYd+H8H+DCWJ+It7UKzJG3q1w/UP7KTKVXWxDrOoHTTbthHfOfSEw9BxnvrWWnTpxUkc
MPYntabnbdK1zs7Se9CQgE8f4fqIzrKPOh8XJkPmj/qwLrRvteJ1hYXNF0aKv1sbaZ8RWzut7uxk
jWtApW2xRQfLEVzp8O+XX85no7xwo1+d7NHD7w1Mgd3vAnphUYcK+o25Ht2ViXUOkUbsoUlneaxO
mb4AHB8GrXgXm/Ij6R7gVR7HORaczrxT/xldEg//7skzRgKqKOB8bnTWh8WXdmLLiFkYMk+2uF7a
GEmgquZzDsOSFBu658BcLWau4eK6nf+oi+WtyLu3eslgn1vzStFxyTGl1KNppZ0pMw3jBbm0DiCM
q/1Pvi3zZZu5QsGNwloUKeXSeLO36bCrWmLQrjQKHBDGocUd2dMkbAnjAF8xTm472+DWIQLRl0u+
7NsN2nws5SITPN6pBMyxg82YZju+uYQ0jM67slV14YsG0r7QBJd41OKIuoHQRbyXUAf1b+10grbH
/uN+uGZp419hjpvxekEWqsezcH6VN+XknokVLIzFnuySYNU4GSSH2q3OMqMfph/6tutBG1f594Ix
pjEg4rDPrE6GnOINntym92lnPUOj20d9L6fPYcjRvYeO2xUbDcqxHH01VXJBYcejrAlxGhvV2R8z
xPFaqApvkLJK+njZiMg0ppQmNU2HDL8eexGEpZT6xG41jnSlMCMfZmVAtehnEf0Z+FBt6K2CuCZs
N2ePMMG8EPRF+epfA7ad7KfNwCxExXrgkUtBHXI3ymrWN2zSd9GPJNuvQAPpFA1BfET/Fzqwwenb
Mya4I1Bncz4MhbWrEEqIOk/EcZ5Fv63/Cj7GMxOkvW8YpJUaoLoDHcoYC3JwfACwAci/zlM2sWby
Qp6B64PWR9KTwBfzciENrzjtXS2UDMDFhORtk21M0zDg7RWZh535kcPmpbsoQacMQzlRwnItJ9Tf
JxTamcYs08GEc11oI6jag4fnz6otBBUcL2qXww8OIexL0tFuv5NCplwy10kMLmicK/dKKLF3TOM0
VkoQKoHFYyRVGmoGDqN7blxreEKsRROJDUazhDnWlQydUJQQ9aEEgLX2UGQI+uxCJk4OXRb/MqPL
XyH9BHkUookh4zz/huCj3eAJSPJI0tGrGQPQmaFsSNcZd4QZlz0JaMwddgMWdnD1DFg55Fb1Gy8N
FnIFleWbZAt7o5JAtksv1YgubDMnQ9e5qirzdDxB71M+bhZtVzwWgIHpbFZXbAK/wXMZRCqr5w6b
HcMMdWbLvubKf1llYprwvy4WVFp53wMLrPVimQCQ6FCuOjizY1DKj1REudhuCN1g0hFmXJg/IbQw
i0vcyq2Mnx+iX1nTDP7k6Rcy9vwUFNSkkeAUnlg8B3YP7cg2tf6+yJ0yqF+4ubw8uwRj/ko92pxx
BSeV7anPfXAwdQTLw6s23QLlS0mORH499vuBybu2g9cWQ71RFB4aeHpQvSNPzKHNDf8KUZSQutL5
2pHgQfd90jqcubnQk+FjHzHprrIQrQzubxcfxVB+hnoZb4EWQaijjubjD/5xnQMvned2G5LXcJxM
OGBJjYrZCRaXP9tNaCM6MRUZG2slq1Rp8p2GSpu7MvfMeJDBbbtUvITjI2c1SLmq1Sw8EjGda0qI
ARRyoVXpQd/qKy9t7YMaxPDTPkCWYP1mPk7SVofOQEddWJho6GGApC79ClDlvvAopQczV32nb11A
YAfJymTC4r53KhAhmlhAZzuOgSY2lmtvlfCThEu7vmJPvh5A5HHlzxOxpAySmCsr3w3EOmXkUrEL
kSHxpT9S8TWoq0BA8GpPY9ZULwdJREHAIHJ9jKp6aAf2O3g7UtyiRtHIX3e8ncQW9ds5aWM0JVH8
VmLQL/KohvMWoAioLfJ2EYrRA9TBWeIpPDAyEujYaDlWNgjPx98mbuG9vhm6wFOmpuCTkSkZKKvY
XvWilsrDAyrgcFJXxAa5F+XbTjraKRzAYnHgPb/dhoy+he9r6c36eIshGhX3GQlXiIYsfLG8sJrp
YYkg0/02DKM1qlzdqwGU8SUvgywvWUHTnAjpmf5O/9I5+R4AIcH8gQFVSBLnPWcfEpYbCSkUdoj2
PLsAO5KjDTo42cRkfQfIlWNpcXq5OS5WRHlHC+pMU2sUSCAlQndbihcE4AZdC+9F+R7fUESP0bnP
HuExF7Q7cDq6NVoaibz6o/ELnnowFwMQWNMhB3TbwnI1VXRKZDt92tGNq8tgUVRz4GMqBqNksMxD
jE6kbvJOrN/AeRnQNjnrIRwZV9dYpB1UT9SkPwtF/PJ5qdRKj10XnYWelVUkG/TKoUfMQlQztPMG
BzDsST8McryWODIP/ur9zV0GaCUZfw1cBbBYvMY6RD9YNYOoulugzFq3NODvpIBEEC2S5OoZsPTv
XpfnOQesP29XNPYGSvNdHfIMcWLqdhWZdky2gqtE0FMSLSXWBR9YwxdrWSvLvsZa2vaVbtJ9v8bl
ouoOeHtycq16Ysar0TlyMcFnOAnzvB7dhCWo5ht6uXZf/1Ut7O0oUAD7iekJMc894M5PoVaU5AfY
xY9Mum49VDdrySpO7nVBtmrGKTN4k9Tgz4Eq4kaTPj1mx1HYKBeeOlQFVPgM9AdwMXKJyio/Q5Xm
2CSfC2audXhpqdGsEJktSDjd8lOErWUbleQBlec3VDidniU7o9L/fPCkNrvzF0lSS2qGEk+OwfxL
VphHo4p7cs0lTv1yBiCwVP2tKWMlulH1vK14SzaIxyr4T5OXb9IuYa7lHsU6fbylrxZbdgHnNZE1
BqwpMLBF8QWx5pIuuhNp0UTjXbZlkvFqZxlh7kZCyeqM2UtfMN3Uwd/Ok41i7qcPbw7qlYlKhQ/g
Hc57zGNF2jr4fOf6f1jZVWc5Tsv/wPf9PiLarhxDQ7zX6xtWX3xEsWysv/dvNwLRGe0V5OedO0Of
Vlo02mpINTjfT/mbynajYeIVu4HZAyUtqJj+D8S5A44LZX7veWLrB0pnQLyY+I6MyIIIVhI6xIVL
9CadLxR5SqjFGBmek987IZR/73gI3zlASsxYsGGb5rUkJGZooE+2/xCBhO+xWIovupHfsLKgkU3q
4F0XzaqzhMXH4QEOkByGv4xwYGZHch+N5VJmcbSPfNbOkDb0beFWVviWL2nxGFZYP+vZNBG17nXq
Fs4HD8NGhxnNfeF7jE6Wy7E1lllpmvI0DW0JyvM2UPWpMjrngSnHI+SxSfp2W125Y/8qN+ycSGb2
J5ZREiAVd7ii6GOle1RaiPmoS+ORjLWkXC8g9MrhDFsB3nmR2yjisU+9cdd976+Lz73HiA4VS7Kv
L7l5aqDZOKmVLF5aodUHDUhFsRWN82kJOY3Ps4rQyHDYx35wL3Li+3L8WnarjtpMD+1fWoQQeYcS
HvSrUjRTVWtKKGPt9zO/JMZzKjCWEhM23WGqSPE+rUlzF3ogBDz4TKa+n/gv9VuBYAvgtq/oqIDy
h83s5aN4S7hKYAijRweY41cko1YTWVD+SEq0VMKwV/ZmG+NLEAQ6o3LDe+GaRQwK/dPW7xM/GjJQ
KtngZMROqz0ppo8IML3Bas0XCMiaKR7JQlSAVjLeqgVkALmD8TvielYL6SLjaoodfLR+yXU+bwOF
8zPvc2UDZNNcagvfdF2hL5GLVEH/bBGdvr693TvZoJXGhwuRB3zB+2FVV/568OuHn52EzAj1t4NQ
LdjNGfRshPDIctq/IYr6GgraWyUl75RnQgr9erv5k595V8kl7ehwqy72JHJe1NILWJ8dgykmeIxg
cu86TObumUyncFiQ/BlwYNubXvHT5DhAICaBEq2ZCO9AdMMOFB4Cb7qqEBe00YknVlGDi0wZOsF6
asCWYhkZSjeRae76iKV0dm+qqH2U/nfjjXjWrzn8Rai/u0QrD/+R+TkNLa6lpmQBe6wMCzBd4HRm
zn6illtT/Qur/BimdVEhy/wy4hlRkpf73PqgErj6jFeU32IMXm6hUvQEMO6A/khvCI5HkXJnhkWi
Iv97TBe4UpLZfU7ar7ZZz32kE5DX2oPQJDAprIQIIbWOw+3ZAYLvHk0WCNHgiffG7trgNdAKwmAT
gTTS8ws4+Lwi/G4j62xECp+mKS7bRY/g1KXOJOMprpd6nQOl7q4xLAdfObwdZJD8baSooU1x/rai
mitJvvZCMy/uprrc1jY0PZRwO6WTPV2byoNmTCh47O3CclVXBePglbxzan4MAet7Pv3+jlYx4XUa
QqrEPqx4DUWWELqvPFoeXlb78pG+gGyes6FCuQHVT5aAmjM4Gbp0+p/3EFo3IcgTYI58L/jkQh3+
fFvTymgsQM/iuEkw7J55kKz6n5+nEsQtdLdfF/O3XgDY8z0jGxYgiSkL40iqae5OUcWGWJcpZQIu
l3PsPXe9mXW91M5w1XOob8d7YYnBnX5gJeW+G6dXEIhaB5TrD1r8s9snWVtaSC6xGoSl6EEWqXBM
TWg8bichLW8b53EUaZw887WMQBvwRvshm10No0WIA0dSt8EmzSgFb9+l0fZmv2Ka5Jm5Nk5P8Sug
jNuJy9tPsuwIv+E0NiV2puDG84dZNyp48iLXURLMYLPNZ5desrpcWU1j+PXZWjp9radjnqPxcYU2
5Rab0FmLmGI2SsTX3E/CesYraevWW7qvJuILFTHTEIXiq1br5WHhU6njDmgE05eAOxjDOKMvBzhp
hnQUMYwyN/qvFdBCOAJy7R0A8zzR2aSdhoUEh2wcJT4lKLcfOmO2MyCAHpMFDF19AQF7lhWXjR1w
WxkUYFSkUr8CaEJcBuBjK8MV8NY+tUdHtchUqmTV41ILBo/5FGpX7a/P4eF3tVr2RPjYU7hEsWbY
TMoNccxS1D2INLC3cxu8gNxBQ49AxBmBpvalgSjw6dCEWG0soBvGrCrpjNzwgBzEnETGJtVHhEyT
hGc5S56C/ads2Gpf9V7W2JMqaWAjX4nmdxGpb6YeGe2TylY6Oe6lDkkw4QiKMvyJhVUTbU82C874
qh5WhKa6enbDa3eFOSlJ1VT0ZxYcnb0LsexE+BloHNzOXazu6vLd3OS7ehCtsawsIekRC/gtW24+
m0RWdEb6ptJwy9L6wAprjBWQ7gNwjgdUG/OmzHPGEBBvq6ci35pDuDJtfocK9bqcUYkASHzrdfpR
179VZtV+xcjp69MPkAZZIn5pgPfjMfWJVe9zdlC/xJW0cGgSNzSVNzJJKS0iuIuMWoqDBQH7vsY4
B4qqMqErhGDAs0EyyWH8/+Vsh14L77/wYOla+jHz+HHWieryM0D4JvVorCFNxXyDyT6bTa423R4R
cxq/U4Fy79qCV+eHBPd8ILUt9HC3DVy3sFArcbJvjGPcBrvKPIaNKGwmkyzQwFshYfIIXNyw2LzB
Iya8lZCP4ltRUH/Hnmcrd4+vGwdttJCb/o9SjCx1HWbXqDjle0+9ZPK6QtVAGMevYMA35HHeFKXW
euUsTouEORY8olaqufSKhPK3SvHlS1KmZ+I9kbnxrkMvWzIXh5DgnvBwRBzWlPltXD+FXyRV0F3s
K5SaEWno7zCM+S0p/XIiO/tR9F1lyUJsww/6APlQXOr+e0TxTHz4Kf6rsdwaFKI5fVUvQWLPiFbl
M/cBZYZqBttWVadzMYbF+Tpqap0rwy2mNt33zmNCefAXJEGSrAr/dPmWQrn8Fu4U0+YyysuedJyk
CmjbFbOwMKxZkfEbdlPWBMuhbqr9We40Gl5hG8c2eMAGmsri6WJgkwfR7EvN8LQzgazwDqNP0fc+
D+bMiOmG8Y4LNEDc9i8b5we9Dt4zL/zdkLOiA+VhZ1w8hWwT51BnBBGg/T5UnI6wPrQ8ejigHFwD
BXKG2+AfEntfkVs4d2oeBbhk9afVD/y5GSTxbTsryVEeqXkV7OWX/9Eeml1bT0/szSVi03NR6EAy
YJOq+hmz7nzhPLr81C/6MYtsWiTuse9LkmMOLgqiu5uCKSPAezd4V0dXIsIRvoGOFNBUX2fPFYwI
1LhHGuJTcRIsPqfel2aJKP+uZtru+BIRvQUnGahmOHvEJhz7qHqGTtr/lIWZCZu7n8VxTm62cA7v
UV8cRHrzI0/2s0vtnyn100xgsiDMnZ/YXCd7YrVRDNsmHVeapmj7o9L5jvfQoTTf582HzwG7+Hef
5Qw8tL6nlalmcYQqQtXHWc3VxqVM0PX3/7FJW/6P/NP60qDfwwa/oQuhSrpOAc18/sf7gPIUM5ed
ES/8OJcA/U9UFjn0VBWhdnRMwsLYi83Kj37ExO85URPwIruyI0JgQKIhZaXDArRDAIR30kWRaWzJ
9vB8DfiehxTD4Oiq1wRuzIkZLTOhvO0hcF7jCZMqMX1uw4cvSKdJKWmhbKcs1KaOXXl87+vfrYY9
BK2oblcOar0l90Whll39tTQebDBXMU0JZelDgd/uEUt6z3MF0sW/uuABRexJLzcSUl06CCz/mfLE
Qf9be5gJ5sxSQLZqqIM1nPQykwSn9S7ScpDzWYmmaGtXBJIuimgHj2xGitXdcJM11I2HsaLYROmd
M1lVusfHswChN1iGnRE5z2Abn5qxO2PB3DVY2sjZZ29n0nmaiMrhl7uVPLv/OZte4yPzuKtJYr6s
GNICqL30NqIG7CEMjKI1RC/GqlN4ILiEQfQOeKAG19767+L0eAWsdh5/QEDyCAGarHK0hapvxT61
gjj9XouQi9IxChOb9/0diitqt+ktEpFGdR4tXOTEtecB+paP8Qwgrqo4UCnqDp1m5HxLjnlSp10q
0dlL9ozcvtEZsJD64i9pSGATSC5/8h96x9Dsq4gMNMlVW8cudbx5zjw1c/GmShFtS4mPvm0G9khX
21HCNbe+Y9m6Hi7q1szId8AiMkevFf8mGNdpug5dDVGyzk3Uk1ocf89lzj6Dr0HZ0rvKCEeUg1F7
BUw9SEhV3oF40BZr2kJOXTdsKQbfIJ2UqrGgKrkrR2TA0ut8qLnr6aqwBtiKxn1aiCQ7X0r6xnKJ
JAzCdscr7CsCOXn/Dy6qQ+4rM1a3sz0ecI6KxBN7mcpdS9n9S+vm9tis8rGls7PLILTVZG3dTOsL
curmHr/IHpME2hwGL6qbM2bFYMg4iGavWKVXJabpc5Szh12LkeXleySjo4fuZ/BcpgrVxaEz/RpU
AQc2WjD6Je7rKYHe1F3O4m1heWg63K4jnuDL3/iivNklF5Nhl3qud+E6n2KUeUTalKIqO3lJCc8x
MN6aKkruQefn0EW9/kxiR2oOXQxbbbDAIZ8V7LIs2pMq/c9AiNJV0AiDFm0V1AKaNp+Nn3qRomyv
gnZZ0ugsPaHSBsjhZyjibcC6gzxYkV8+fBOnNCCRNStUVtTNtiaNuPoT4lVzNpsEMTpXOy+I+4hg
zzvlc3MAMQL2ua0ySqhp4qhIVJ1ruxEQjE3QL6/zh9HLi1Nh/JaMxKre3FFJu3e3ea9L2wr9HHHK
NJ0ctmnZYjKhr3tKixC7Ooz30RuYbD4QjA4yJy+uwHA1V7ZKsvhIp7qv2pszONtib5NJ27Ccy4uR
gRaLs4d2GY74DRVZ0FQbFPGsPAzKP09lW6ZGmD9fpR5LHIpG4YJIYLvU8sA5EZXr+p3Uk155ePwv
KYcAyffq4LQEdNfQNFYROjbolbd+gJcvYH0J0bZRql7+2e1VzEap5HfymBDtIullgxEOZXbsC8Cy
jGha3nkzWkcWXOu7BClfMgLf2rdOimza3is/+s1kHhpudz/jQiAzJy4tcOI2VhmfTew1fikk5KWZ
03851aopH7cbuXvoToU2ZaUtL3nFc44Fs8J3M6QFNLzQBbJx7iDgrKJ6tBspCGhglCYBQcMmqlhe
T76j0WPeSXN54/T5Cl8p6geFdgQDRf7A6dyAU7grcYjJQHOOr6e4IpaKlatWIov3vrdJh+0m3Gp5
BVnnjkfaWZFg1n4KgeDklBP9Z7zL0R2kikNw+oyFEhJd5Cg+Vp205SoUV8vrnH92M6crkY3kA+bx
FiDv45KkZs5eCEpRbk8Wl4YT7HNMAQnSqyaoIXquPcGvMDWLQYui3d79wH/MD50cAXTshYPZo51+
IUXCzlkOv+Rmv2yXi1oO86x3Qy55onpmitK6jjNYBk53G+3pHJuwpLz2g4gRbD8AW7oN9r4URjzV
dSrTgGHxLVZjgMK/86dI7gTT+X6WckZkjaFJtZwK2hgaHQoKl9lUMP46PwFgmxXxcjLGUdRe/3bL
+5TW+HnoJTsht2XMNzNtKkvQn8bh64tQf9CIWCjY0s7ZDwgkd9qkNvq5Q4cdHl4T3+sMVeKReTg7
Kr7ddsn/O/Us4UAmg011C9cC5DlsClmUXeFukMk5wDKHrRxzS4oVhuBOBLje9NJ0uvcpAKJbHenH
9oRn3Zph8VDUdRqcSQKWnXaXZTdauiGSqacodxmKcloq8UMvJx9yEELnFYCXv6rq+iuPxyqi3wUm
sIVzf7htw51Omjs3I6q0ZuiVeY5nF0KyHBW0K1HqibUjzxT13WS+0fwNNLRrnXdSpCCVtZhdhLoo
4FBI0QxdKqxXpyhVfmsncobV/mWOqV8qnnIrQTwEp+wzUmJWZNKDPaytcT0KiJpDacX7OuZofZh3
Wak2+TmBRm8zTOMEt++T10u8fVr69Ma7pANqJ4zj5Y6UX3rA8u59bNmWSTzsCgxiVPQOrBR3sUWQ
tBljm4+FbhA6PWohYBwqV24Cd4hKmAbFyMrRoKyKQTB4PFMu7rjXB8HP2eF/YXsecTtPtnDDTdgi
GBiETWaKRq+C/G3ZGIQm80Ja7rbIknAjASYdyVNmDT3OAOXzI8WWreeP17p9OQxBWloE8iUN0aIa
iJe67Q3DCQqmLx5jhNjbrIQbg6pWRymuppKHSI2nLaXhoH2tK4H+JeC+Ldg5WKU8doTsp0vm1Oil
rQa2cumMjVbAxLaBoZ6iloBOwQvhSg1QrvD841PacHNSU3mzTdhyrJl9wMddAEX3ogCNgHLFcUDu
abBRMPB6qlQdeFAhoQWxxOs/kxgK5jzBjOtlu+DYPwqQV3gUhkiFR46u342udHH20wLLwpJW1rmJ
BU4GdFqgBl7yMEZzq7owmnsYBKHflZc0Fz2GmDRIPGUdowPqW4Dx08W37E0ghK2GmJnNFvodv2Ax
yNDLFbZJdxlqOVHSwEFP1+PWLKV5iHwe8m3zZiWuqTIH0gVpjyS8jWm+URU+kV2F6UZzZqL/9X+Y
pSlIrDdCA5E2e3XBdo3BIjYWdJap/JTGDQSDcFKPpbmnuRThWL4/ebz35Jl7AEOFsbrCjlKSg7+K
MOMm3CKhnAM9950J3zTll71e6qZ5rt6W6aPIj0WWCbaVVsdUbli/gMkeDdzHJotY72XrU13Rxs56
GKQAPMj6gAq4a37oUx/ZS/g0ZTmar/IX3FmGtLYl5p4YaXADErprND5xBnDfsYtszx5f86q2+iUt
JOr4/ot2awy3w91U3Oj1BHqE2jh03zOZJaeNMmKIu2hh60N7FeDobilTVxio0gwfXKsmfODhbmmk
IsV6lY4EkftOjBw+98u1JuXRueocGDS5yg6hwpFEowACuXiHJAP4oDMzb7iyGQ7+jn8fIW1zrxFe
3yAE0vOitoXWn1Vs4cpur8qaVkbeYXfSZfBvfCGdHko3ImAdvA4DZCP+pPWqw8MdoRjeh5HNos8e
uMspIDyQAt1l7pfPg9gwF+xTioGdpMls+2ZEoTCz27BEAGmQ5uDhe6lN7eE5PlIW1P52xetYktPS
/a9svIk/34GQ4rJduNnbQt60Xcu88OyEhOtZRpqYP8jWFTUhJJoTTsEDiYP1QI26PV6SkD0GIqyI
hVHPIbX8nzPMtBYTtq3zytR0Jw9H0cnIq7CBpG6bEyWIO6JiRPYtnrcQdnz1H3P0UrR4y1clCe9H
z8FxShFMJMkLPBOPU3mGfcvzdz91e2D6A1V8FwfETAreQAW7WbYOiglsk/RqcG5VCNk4H8hXopxA
FjSwhse02+Pbba2wrpcac5U7tBwaPJhxE+9yd+gccbQrvDo5Bm6iHqV2CrheSXLLGhA1oBP9cSeB
trvzB1Rp/QhQYqOD38SABsI6M4Ibz5ZR5mwSjQMA7lyuELWgq3Kr+JAFFre7MezUBnoR+TNiqgNz
VDCHFff4LVLFfkReS8cJ7uaGZwUNzM6JewYC+vzXNoA8EMMh+RRMUWOZqHQri3iIvhQcz1LKk0J+
UJYwpR3GPXr6C8mnlUs+Wux+3fRt1qoSPqbXV6/r/ac119mG76Z4B3cSF2r6oEkEbEb6+Ei7j4wh
3PAuXk6Eo3HOyElFFWkaSqeM3YXRVgyXx36/vD2U52fm6V48x16F7UehFJaqxPYxN4a2DISqUGed
Lm7hW1iLcRTEb+i3ayy5QzEQECBt8oKlOzZCtP+jKJLAOfB53BqG5oLyV+Ot8L406hHADHTP5KWU
hHf3bwde/jW1CwMS9e+sf2Y3RD/2uWTt4Iz+UY4GhAmcaYJ+CQPLjgNdI52aEyDBMmoQG/TUYjUS
Xkx0KUcDHw+nguZei8YjJfEst73BierB1MGGM6UkvvvpPxun4j6nnhujidUc8V91J0CV9gv6ll/v
HY2vUE4HMVPDjeNWw2WTpXoATfIlJCWJ1mHJ7OCkPooWQVtvgH7YIaXKgwU9avnUeGJK0Z05N1fp
li4BQe1Deb2NEYqkweMtoRRv4WhhUuCzowJafEf4W40BQF9mazqVwS8Y2++xR6/xHTYbIgGOW9iY
WGvPgbsiuzcOiigSC78ddaZkVaQNW6a03U+4TgCvFzAzmlOc0n6hY+cv66i0iTDRAVAYVf9EWlKp
RkyLSlOUGI5ktnAi2nBD9NOC6RQOnibJKE8gL7ZuLmOunfmz/vFGpjvfOmXxwvPGvSCZZ1/ZJz2k
2UrvLMNZwv6BgKrRfN24CqcXTxbK8cTGKJU7UGtKejQm11fuxsS7FT3VC74M8Q9tqV0GGk5pZ3CG
KcvsdwYdgc6Ynih7EcAvHeNkAK1uAk8+PHLJh8Gvr801s34e2V68uQhlsNnXsFMeTIBYvd/X2+VQ
GFrl41tEmJFkIc/s+z65M6e6WERJc3N3tsIPb2vvPSPHpfOi9deDkZfl+tHmQqYvVV71ikF+Ec8M
qq+JmeemFmf2v9rFw1hoYrraSjLT+60fwNDuRGUbBF2V1QEeuitgBaP7emLepZdxCFi10F+d7t16
mnEDluWuxQVJCFxBUC07TEnwFO6BGNUJ2dlN5H5hGGB4K6shm/Tit5e6icQXlysKdJXq1rEGr7+W
CyOMunGT7Air/8SZOtZ3RwpZuaqHQndeiZs9antZMRpi1dFTxJNCpogRh92ppQvL9ithj3JxN01c
hnLFerqzb7nDKfjBtTR5fwJwW661lK0BD5zExdzlIc+txmhxknc1oUx9HSuAS8zDO9y5dzJJUoBD
udVzZC65BXQmZmbRpRtfWayT1Qk6F7Xa+o4uQgyWAoyc1Dzx9JioORa1mgCMG+KUOI/BCXL3Rjk0
cPmjv7pkcAffXuzdVpkBDZpEQxEqwwITl41ZezWQZxq0mqBTs8ZvUNGjCuUPWVB7FYmaCp+hwC+h
95MViZDOrC46GL6drcfRSR6nsgZpR/oOkGXjKkwq1qPlriLHZwzluL7m0xPIin8gzgScYPiuW2fZ
0i7RS1nDw0bCLL3pFDLaImdD7Rw6qHvo14NABtXZSuuysqUImUAk+kGxVwQ+CeW+PSv3RJXXjTtw
371Fy57nH6Yb3PVLD4gHiv44/0A+8wKosoZJhFDfhM+mJCyeqW9ISj70ngrseceQOi6gfrz7WgWH
xfpUu/C07MjpnNgWsK0zS7bhvFpw8aVaisWlh2uHHMZ93D8DhNYTyPGATMn7NCatez5iU/B4fgDI
jnFvJU/kLRuL/4ZwQQLaMMN4qQHI8TVDOXJAtMk1K9NKLqfyYP/Ht+as5OZJIMS5J9aVvN/FRihm
0JAgDLilsr/43tXrwDKxwXtKvmyCZ6OyE5P/P7xKsyfqbpr7ugYgaVQWyUN2rs10BuNR4SPx5y9E
/nBR0fJxkgsfeczsJfCvBJY9fPfF6JQnKaqxoejtHAzQMXecLq+N265x0d8ja3jUfHPNrxF+bq/l
OzA2xZjx8vhVimvquh0X8pWPnSJgiBl+dB7aztPJDoiIouyw8uIW897kHfWcjhwsQCfooG0ww30h
7/cY4pYycdy/ajI+SUXUfffNdKtTAp9/7XGd07ou3dWUpzlXjt1yrISM7/Q9nStI2tUR4ljTg/fT
Ij5S1sO7UzuDz4SCUirJl+4koDk2fsAsEu0CLXiazHCtD8hsaFijwrblRoMtewKmOk0ArbdLMne6
RiQUBeVThCeEzmuLsY6g+RUrZabV5a84VY9Z/VchyYRyK44nmDmQiN0QtYvnog/b/W46wJF6mJ/m
Qaq7hNZN8/EPZEgm2NzFsiX4YChROW84ipI0Ij0EMnbBJ6YaBgyNA8mOYdHwKd8gtB0+KzUmExsk
ykfzVuJyAQTy0UMDo4GH+jXF39Qz4aLoaHOJxpWs1D2pAGFdZu+1MQ1JURxvVOdH6jLpqRjqv6NN
vOJQcu3l1ViL9F2ybAMWDX04W8XVJG0cY2LXEN5cVJzbpz0jQBWk08a+XTCXlylmTKPFPZsncAWl
wtKnjVftntrb7PLDGLpXEY/lKUKT65Fb3hHLjFuMkI/tW2AqBv1bg4E93i8ShcqY4rsk3Jra2i/U
cqUrJN59qbib9q7ydC2sFcXzMdGwlXBYiz6/MDSvG6e2zI56pTV5lthkbhTP95QZoIGiQT/cLnp5
HD1kRUV9Xuaj8HBGB/Oayrl71HopsLHjf3B4j3VY0SyPovFxspoLtWxZgO/kWBmlWVEif6m1DRcp
IlfjcKJmp9l0UA7W4kV2IGBvAvftbEfYJMp1e26abxu9883Z+0TcFZEUV0XHQ7rlnEykDUgMRAI3
cYwXCycKFUf2hYYjzn6r4B04Dyv87GK2s06yKosZdUHXFXfF1fOLwFQMN84D/qqC5kRUde0dtaUI
WzMFoWEP/frsTlEzwpMzJ2tctyWotRDUIlLwk+i4ebD5omK6S4tR4SGTk6gpt1xHZDjCm96M1LOs
lV/Lqdn3XZKg9UOm9LgaEp94UfbTzKEVnjF9pEk3t2ZEX1HrxC0lMBKtkb20qscf+dwL1BoregzD
XbkNx6JOB4CdFuWsiXmjuciAloQsZpCH2947I+timrAjJy3h3crtltSgT+Nshbji7NEQuw3juBnH
+zBx3ToNNg4dZ6vlVpv/DwCFAqmLRsHlE8bM+m4Q7iDUDEesl3JVZ53v94Q4e5w7Y6lmd2VgUQTK
ciCoxAwm+hMKlSDkAd1VlvoxApnwmcGoA1GfoA9Sb3ul3MehCQ8bW+kR86eIsWbULFRT1PScrn5a
Vu4YMKVotWsmN2Zl6oCbiKt2NLl5Rjo+AI2/w8Yuwxd9PtPhEcjjCOlHd7sUBiWjoY0fw1xucquy
iWHivVePMERXhYU6MZFyi5o6na/rvDCOYA5ct9/oAqksWW/1/mw7yuBPZFY8rj47wDOftDQTTKIB
2RDbSNOhz4YzbGYKnWukrmtgwHQEiA9zK9n1AdqgtZMQMUUGxyLPGV+iz4dYUJCljmgoDZtd2IU5
wbTZ4YMqGh2YAQ0gcoBa99sCpLvzLGLWTZ+z1jEpgS2YdVn/IaYL3aMLr2Wt5njAK2MxO4xwBg+l
FJPa+hzIUyLurUejGO4Jxz25f2FIl38OsiF+uoQmaQ6Z87o6JmoJmuk1+GSGU/1Qch0RUraHrSBa
OQAOUlneFH9GvwfLRFBywGsFE6TR8Y8NLhS1jsr+4kDBdTg5Qwr0xWEec8WHU4R6CbuSuVErhjGQ
Sn9kuJ7H7kK8mCVUEMnMYvaArrOcNmt7ATENtAnZYSpkW7mOKkFce1YCSBTSdmfy2l/dGoZnQb2Z
iARNK3A5CJ/5VwxGg8aD2lVLkCIutsgfZLOA0yeBxtNzUdLnF7AwtJBsk8E/aLcCXQeFfO+p4mTu
WcHOXZDJyENxSoM5bMUjZv1AN/TJ8j/Mbxa1tpFit7SezngTmJiMaK/6XUqM7mi99+ysQ8mv13QF
m+vPP/LrKq2paF/tzuynwiDab0kHas9YAlJlTNI5MTrqyokkyWnIkTldWScdS7c2GFoGKU9t33ya
6JPuZdhGVAzZafnpPcGctkjbMc/lHwuW55jadqLKyTu1s1qlb1IuTkpUHmcH36AICaEMmatnUDYl
dnFKhrC9sNe1tdTj7HmxdRuOepc690DwC+VIlRoSs+hkvY79MHEufzh3pWqk4Fnwi9fxTQYzyeiu
2IwuOa3wL9v7EZny6lkKqtk6GFOy/5k0+cJbfvkYpsj3kk7fDUbfH9Zd3fS9lw8Bk9YML+QBVmWK
w97Ol36/sCb9Zmp47y/oqi8i1iCjs5nQwpbMbyXd36F3Q2GL/N2o6Qj3ZeiOhcbFeduAfvx9D7UI
nDML7BD6cgMwJgkyo6JFpPyPwImtixmqJhlW5cU6JldHBAOYu/OtxahZtqmdxciFQh03sWWNvWO+
ilEzZlcSwLqAc5Yr3ZND407lq8mO1E3MiBOLTZtOr+9d6LGV87phVCpkiiXDBYRNRyvGd6M9N1ZP
wE/Ru967o8LP93LzeSBMQE5D2JxNkKPBN81FGY81xluia53DzXNFuxhchy89dRm42VJg3Misq/+w
oe3PP9h/38zCPbS6ngKZiaapVvyXSbk6Mh9kqkPFm+jQG9KM1ou6cVdBUchjoyGF7+w8fcUvSWsc
nRglTNrpBFckIm6PUyF8CIZ4DJYElWtYx/i52/Lp6e+qc+NQcimytW/NUtjgeNb4HfDE8cVXN1Ck
SSGm5Ux3212whVAgmsbuzh4nzIzfdP3UbOoc+5o0F/da3HhXhgk+AxxsWGw+hN6zPXYkq5aiwN1g
vK5x2a5rkwbJ/2zeLGJyl3dNQdREKYjWfrmNbUX2EprDfWRHavN/Ff6EQzGKnY4VNfcmgAaffmE1
F4HFI6qfTmSYZHQJF2LPapWPfv/hDTg4EPlUT3NSq0dQ2S9gmEUhjr8y9DAAjMIpKU7H4Am4Wdd6
jgJpVC5a1PYVCmvFsAR20Vflu3zsT5TDUS/0j6SIR0Reo7lCK4GUFO0KZme3CKzjscZNsmBhQXJk
CTyyxwZn1Y2zVUnkGjfHwvtzHWAaX1hPINosEgkTcy/u5n2YOau/rg1u3qa8VwuCjmoVCY9GTjEv
SrYLX5uo92vsxDHP4Q5O7EDP1wTw5MCTFRi+oEzXOz+CrWCmzBNXmq6C3VhUfYKghUAXwZ2YbDIc
q6Io6NDzI8vuIk037yBt4xPiAAyzL7nQEeSxkgobI2/GvrPoWdW2n45JQa4cH3nXEcsc4Z908JuB
4I/gLss3QlyQFWglLdK/FWXeqGELmhfqy1xS58N5R23XUv61tvA4zZ0TKw0C0r8/tMNqJ/lSjaMS
TAogQZEQuj5PQgK4RePJ1xSNaoOZvGKStV6fpOHenBB9N18sogfjCNuCMyqHZkkj1z0QX8Rj490/
fVLkRq1yW8oznjJya0yN6s8F3dDwN8hoZIAcLu1LVp8XSLwAKY+00C7S7TxMe7TxfUL2QWvQoV+C
FQPc7NS+LrKt8LU2jHGBXR+5juXJiS0HKKTSPacBIDukcVWb8jRvDE+IhRJjgz003acr3Irnak6h
19JTLxgo39tt8W4BkczIspp7UPJ6KYyYezsY7SqXTykIJeC926x8Tul6j9LpIMc//DWtB/wrbYHZ
d0apo5r/vNeqDDwIAgzv0aCDpFRDeYDep0rNUZ0b16UBSAvnQ9vgWrS+Ncdo8ZXC7DrlGYejAhyE
ANfMVvsjiq9DgDa2dTDp40BvG3CKj/DlC9SC/nKZyazeYgc1+5eKHx0DWHSnSJu6RbB4irz/7bUU
7aQvS1gZQYLIlom07R/fH21ocDGLpXStO8tOt/H2GnASZ9w4TK1aSMrQkTNivmw7Br1z8SSvZ5gs
ZZarI6k4iEug+fhAinkATH/7OZGXE9Rz7P8PkB1pUQBLc36qjnAmOX14pd74U+EOL6G0iMu2dUOp
4uvVgdfC0diJy9WAyVRS/d/RJmPmZ8z03cfXtYWFr/bCjefnvfZmoOSuMDlEHWrxA5WDTscrg5sN
FEHYD+4ARvCWeEXq+iLu4YzQSS7f/tHa7Tu16zaV6Fhc+cE9QquEM7fCxBOSabbpK+fRF5HbqiGn
VwwQFPba0MvlXhTg83tMevYlP7x4FC/VUcZ6N2/EJPANuTGe1a7G89Sxhdm3XownAwsK8sBbyb5n
NjUGKigEfAzOEwsiB8Hq6EqTlaiQdOF0DqqOCi9mmukLmw0L0dPgrtr0Yt5Wk6Jo11Yw0lX2aPp7
iCkiAV2q7dRkBq1ChqNuEVfBvbsQw9LFGY95q7esKnobTiqcgKsuCAosruT8QVf00ZXzGJqVugXJ
M2CH5V504zoePZs73eYKT6MkUHmrhHk0nWI3Ip+NOURUBX4HSByUkcJny/vQaZ8XRlQ4f7gXhi0P
c08NN31NiWXwn5OlQt6TSqZnZaY0wFXNa/HHwZXXaXbUZesNqagV+HRuK67sdl6EJsTheKq8c3HP
lGAQLtnaB7cnFucHAZQjpUk11mnyBNhnrjW/6SY2TNxKsLDZqXeYcxZ+QaKQKyaI2L8XLc0lLAHt
hJmd/rJlkQ7lSAs0XgNgPXxmzJD3vo4arkPRlxcPL9m+gO42MAy1JD7KJ0PscSHPEkOnPc3dhX5z
4rSYzBs27s9ghhHvzils8o1Op4NOQwyISmgQ/zLkNZFvnLfP0EFdV0XoscEAHwRaEiJkySY+uJWO
YYs4WlLGgj2dvmi2A2b15bbdMcIpmljCrixisdZcUkztpVe7dh854syIg0AL/OzASjn9AcVYnNDp
0FjHQ4r50mwu9Diq+Er8ahl5O7di7EoUBWD6K81c5TTzn/RJQTpREUoz3rTebaghO/8P8AHXf08P
zYzdmnAsIo+nbYtlgtyylUnWOqO25nY8l0U3tyrvJH5sfGjLi/vC6R3peVfR1i4uFck9bxZk5TwR
qscYBYgxCNXPKNfoWkHfLPI81O2h1eXGl68rTRn1gVfP17O6S9ujeN4VDCwIt5tTS0Jg4wu8SPD6
EhkLzS8jD4mC28kirURmEJkJBNMuUXTA41CPkbfXfdpBCw7zmw3vw+ugUuWfeK+YrB67WIQNtBIE
utwEVL6mGq1BVqqwR/7fiVb64fprSUtmnYAa565bVSo9BustXCjKqJBOcA0S5Q1tBXZATNNFeBBh
9aJorsKwzdvgpvUOJjj7tMObzZWsXiNP3lVgHbCfYUyHVlpXYJYoIes0ivVQAXjWlQgCGO5EOYNz
v1TXzqOi0gH5EK8elPutXe34/LvpnuLE2AOwsXdhS95CUQetXts6aKSsfwyhu8d5dvjice+ruoN9
AlT4Hgber68H6Sh/cYOEOoT8tYpiDXw7rIw+oDNG5k7K4LvGPA5JzYkMyZOcFlj3cEdrSVgF0uEN
dnhck1MPBHq4PaCRQEXJw19rRJO5u+tjw2wC5a7MWVcJtZxJwv1824fJx9xD1ZU9EUzPhKw4yS8m
d4f0GqK+2/cNEGW/3+RCpcrqhLnjAjzPCkPseF9zGz++ioQS+JqWKm2pFhthLvUz4B61ZYcORI6U
CXSe6ZXHnbInL67fUC41Ng9zMTdNyB8XXPL0MdQPZCE/00/NMotCJVChrowOVs5FCMPqzC36MCA2
O39J9VWihJBSpKNeI8FCCLPkr4ksSARpYYTKrURo02R8eQgYfEv6UDz8fn+Ff0crfNJH4HBIpk/a
tMc8RRYFmreGw0PpK4xVb7MtWcmRyDkLPXiQ2ZPUCW5BXvyHimeaM11wmZrF6H82aD0uHcdGAQGH
yUcibtI7n3P05iMy4sB5wQmVsbTqdpwD09uXx9fgRo4ZUUAAIkItLgpvZxiSAh+VMB7KU6bhkTHK
uR8ptlUv31hFYnnkWOWlzo5q1/0suytcMjfm/rpw5hl8VWJ4Xxhfv0iqf+z2jH8YKvAL1w3Nu/v3
uCabKZMLbejGmiYc5wser9Vw15f/vQr1cqXXSJwC8d9dcklyqLtpYQ2gPWgJokN28gfrAvSLOLeE
Dj1EceVn4CcAvtSXJJLNhDE/0jMY53fwQvUKJbMGkt69xaZJo2GT7ppPg+ZB+uDYhDitzC/q24KU
D9wvVOYqTaeAwbRXIpqNR4CrsEerTu+oRjGKtC1md3s5E2KMvdH43oeskjjKSNd3tV3kpLvpqC3S
MoluxEyfrgwnPYIxwVks3CB4vFLjvP/fTV+r3nkplUJC05gxfur19mdFJFmlatVZ4OO1p08e3QgK
kjwRrf7LqHEAqmUCUGnTqEG+c8sVh/GGHYXZRcfGwYxFSD+9CMv/vj9S7yBA+Pj1lMcuaKPopSGL
vhvfxfoTvK/R5KJba21G3FINMUXWlLdPTtMPhOstmdulsVfm8Fx5OtKZhTnVGRem+re3JCI8LW5G
RupPNkVGarhj3mkyvlNP9cIUQRn518ysrR9NN1IQLYCPjZ84sK1pLmNoDrZqhjKtvJwwV9Bm1nbb
J8u9TxLQV9DLiVAuIE3ZS40jP0ArJP4t2FbseylSXTJ1RKT2lV9sssxS0SPMYybPzEvVwKWDSs1/
5Y3wMtkpfDB1vs4ux/OEWAeuIMqNsYqYiNsydQNE1ZI6C1fFmRxofaaUiM4rRr5VYHic6XSYGr7E
+5BREn2MchuPLWD4ygZvB59ItTmTAYfNcZrDQa/4vRO2CatoV+DdtYbpyIhA77p35hZtyoeJ0TKQ
zdVxOzMjuRDWyx2txLP043BYAWNwTPcYo/RZq1aBItKBYhtaSWONLBdOfsfpz42u4vwqtiRb9guv
j8p0jmPF3c2SYxtzSebvjNeLilwWJ4Shlco7eC9fUaAPSFKFcK/Exl6me6ePogQ71RIY7WofrlRj
KbMygGWuIOCIGCw24Gy8O5xO+cx0wDCQwzfoaORoD6RiWWeunDiFORNaGRzI9umDw/0iiYftTDn/
G5iVLQzVyBgj7cwpmbYwHujTxhT9/HZAcx75QU5uG3C/xlQ8Mey5olq31Lq6gtC2UggFd+yX3rt1
fAnrQnPKK+xKrBpn3j49PihqjPYZzHI/V1AJ4qaabUZDQy5/Y4DXzQm61E3yX54g02/EFy8wkGxB
WctKUhnrBLzg0babYe7mStjE9zj2QiuCLJCXhK0fR4XXuAtb/b1fhfkIejF+aafD4cF5XYDk2Wx9
9LRIF7ceiMjv1gu0a1JRK68nYlYvXCgfqmaAdl7eaHakLRbt8JYGEu+QeK+zUNPQKrnZ/ZjfSs7c
E4zW2eoawoIdzMV48stnnG+rs6Vm72pz77AxJbofKOvKNB/zogrvsg5Yh7KadxtXcTpQ2OGmSx6p
IVXoV5XH4byo7inzNcoTwPaqE60NTQEKbf51h3PP75OK9u2jqiHTumlT/hD3MFlALyRR4vb5OqEb
s+ngUON+OVYVK8HZP1oiEUQEKFvkVXMqnF0nmaO+y+xg51Saiq1HsprUQYL6vYNCyXgKOiCCWjqv
WNctJFCQ7LTeiT1TXq7xWc3CWklmGjJNN8SfCfD2kNBUfGmNYuGW2NpijzH29YmYZXKGYRY1pIge
eGqiVYUVEUAO6GRmGWdkMfwsu6MhF9vqn4AAXLX9DWiHerNOGGb+6z8lV38/sPI8HsvNvYEloEZl
bEY/tbkMhBZHE9HvIsCtpCMQF4WaNlXL6nM09yxewaPGLPi2yTyQVViRqivXVJxfogtp9e/lcCpa
SOVMqeN3yJGzX4S8E4yaB6x10vARd3vUnj909Yw3eYXyt662Elo0aM8aHgvG7P23QFhmC/l2lFr0
x+wRk3c3LO5acFoTpzL/ATKYHzdUkInI1tGZQQkGA1rgfY2hVUaRhML6lExSQvIknSpoNKdHi30u
GETjRIK5mWZZTkJLigFH0AoXcxsL2e044xJyQaxiIxU4O/KSKY4rBGQ2hbMhCCThMukfpEA3iBow
uc4TMx0pu6OUuqsBmuXGaEuyKopgo4Egd5by3XBzw+wje88w+g6oIMQvmHKaKC+VpvpFXQXi9l6V
brnlyz2GFdLnAOIUbglPKcGhYh6fzhWZn/WUN4Iq54O94ZnEnyI7a/7LbY/xSlRZgtE0xQUHQspy
c0z+8pNfkp3hAXQUMO87M3fm1uWdS7dLkaVStL8b8dS0UxNDIvA0yCfoGXen3E0g4nLeBuANR3Iw
DeFqTaXPHMLDAVQ4R5dKBM9O3u0rSp5UHfuC7dQ41D+HmQOV9I4fpxO5+rTiJNbw8mR9loWQ9AiA
fV187SGMql9SSLOsQV1LN+wDoxSlHjEzeAtS5UH7mliA7RiQN5p0I/2gcNGS6Oi5NaohCFaXNZk4
H30PlfVM9iVBZR7kWO7JiSOnBjKJmfYp/MUXJJg5+ry8jGwmGGfigH8M1R4t+zfA9PFEGWbJH1sw
9i4QzxzozVDef1MyhFRgVvOSrwvD01J1/0u2U9Qt5I0DnXC04/oH5IP0pAZg3qs17bQFp3UC3mNW
N/5QT5Ox2Z83B8E0k//hjsJDL4AAFtk/AmMb0EidIrzrYL5mfxhbdbwcfFH+iGWOR0wSa8UENhqC
/7iA7LgBNX3xzSW26yUOCXM5uTBBTsSmo9fYJKEKl72vbb6ogi/bbAo3XA8LLpdaACrUBjKR6w8p
PqzOeoLuCbCksZ4d8N73e022h+nbnRsUaY0F/J7bOTOt97Rj7ld9rIwxNQjCm5R6R5GkusPar6t6
PtCUvom6juTv3l0H+XiYKYo4vkm8dXFzUfu8HBkGI2rKYvjFS0XqUWzEMW/XkFhQxduCbWcXgalo
DtqtOkFT54IKqTk7wHKEpCNASPLQPemYXRe4xs3hMQ/US8YAHnMFzGqQh5kvaTzH8sVz1977QIhC
aRhTkrY/f5oVO/CM/q6zzek1f6/6WAxCz7YwDo5X+XmlBUhY86IVJQjhSMWtg46catmLGNYF6ORS
fVek7ay+R6XrCrATVzxGglpGIWSMCX5QDz1XvV8xis5mUiBDko9WhbN7yqygd171J/jyX0p37aXe
Ylcih65ZUCkiQrMqWxP96NauVZaQFaTlzBZuUxCSZM95WkCc7aOuaR+Wej/Nbrfi8e/mdTzAfqCz
YK4mxL8lWJ3SaLaaXObF+mRFJMOvzhzm/sYbQfOZX51aoTH/u0noIip6dgsVKFZkYOeagtHAvmz7
GoChxSzzQttFPmn0w9jyZOlny7i05JE9oNtpuND77PojOAioxp52woUyi6oMdhg0j6XEmiNx3JOR
ZU3m0ZrpH3bUZUsiZuA7krqx/fMfw8LIVaKL9rl3vRrHZvfx09qjF3Sy0vB/5PkachJkdrAchD7l
TdT8A5fSn63ueDgP8cmEtsxdwuV3GDBFxQqI1/Bm96jrPSxXAlRBXHTaB7OTnc3porNq4yNmjj3I
6Af5kBiio6klQ3wSOJ/v6uSgJfknuTArqOku4Mx1qfhdnYiEE3/JInedWFA1DjAG2WIOD00C6z+K
99zY+Bq6/c5MisIXQ+S/B3Pvx1ztkwsHOovSvWcwuNYtqSo8Pps+kJam+SGFVSlIvHiM4Zi/05Xm
dcX2L4/+VI2+IC0tlJWgt4+7uRELOgKJCdT+I42Qza3vUuFsozgWzy9Uf4jcP9UlaJThlafdGL0a
ksCezGA/iSOX5YpIaYdBfRvgc6OxOI4obcHn+f4/8K3kZMQezWnpF+RJnNFX8BNNmrV8BmxBXGmQ
mc7wUt2y+42kyCjPwAZ8/dk32E6zxQ+q2eTo798yZakbMbT6PyB1X0+dBjTrqRzsZw771IyMlVKq
n4vYO0RRzQG/3dAeV25ze/z6zQNu8dty4stwPASgwErG7Umyxgng0cuER9OB4cfNtWsV564esnXD
TKjkZXZPg1XdXuXyZaFC1Vtl+Q99PTKkg9g5vi4VzZKAkQ5RFaFYZ9x11BmRt1BaGqC1d6qxCoYN
VbAJqNY4ReOI4v31HBUkRj0mwl+qPAbzWvCOHuVRiSOCNM7fp9V53fmQmHkh66pH5Q9Js0OPnCOH
bGQq1aZHt0m/IEbs7FtMyyvdjsP2r09tCCDt9z/sFJ+DmFW1MKFuJABZOGOTF0ifKBGxfNp7WseK
JCROKSncHovXtU3iODYWmOCxwo8soFrJgCKxUlWtrsolXZV1OR6Fte3VWXNM/cVfXF1pi7rvMsVd
JugjbQFRkrVTrTiwHFGVq5CtFQHuuayU1uf9/++d1gLG1mO/nVIl2tZCADe2Ql/wrpUXPAITT+IX
wSTOQTsvmLFpqF0M/+i0X+SQ3wxGz4ofFrnvPTCQlxj8L4Zf6PgPBMtUe3gYX7UPosDjvoNA1WmA
CeSH5e66E0IzqJGwhH5geOXS5URHfnECxjf/1VIV9YJFUvG/QLnTiV8I8IKUlBg7FJ0klJmABQ6a
BcQZkYbKQrxZEmE/ndujEAM7YF1P73sCrcqqM6hqHHcqaM2XXHJXTeawyHewpW9L/uqn6DkEU0dn
7KBNLCA39IhM0oOhKo1l2cZf3DR+BWlF9w1EfC3IMoyNbE9gv723PAViLvxn+y2Zo6rUUgPTYKbr
gXHEfHfXgImUqFPYmq/BcvpGtUC45eIVz2B8L2iVwvNNY4CD6zjtwFmx/Yr66FIgnqIOJxX4OiV4
5Olai82C/FLbaEq54OKDxpl7c8pdwxoC2VmPxnKdsMaeG2VTfptbx8tBKN0HC16bxQvvQsH6t2OT
hO0AyN3u+8Hbo/51uXoYcxqztqrtrf7i/Z2WHFQTIm7nomuIGWkCqZtNIqJJswFyhxFGx8Jh/eYG
mvehdkq87PN/aVpyz9Bzt+6IIl8dclXc+s5GAq2NF3BUQqCgRX/EOj+9b25TH0TxWlKu3pHpBb+l
JkvqU5RenSJnQvGNDZMCnhCD+Hn8e97OQmItxYAVv8eBbEJAoRLVHtS+p5XdLdimb6IE7LsUXaEL
P7+2hfHralKa3gd8Q6B0zrOI3VjeHsZRYYWkp/lA6Qpb6Jh/DNx/5XefVFm48PzYQAE4xqW5x1Ub
9OzImgK6mxePj3zzgm72/twVApuvW9R78svFrcbfwlcbP4HXcobTWFFBZpqaPIARjStc89/f0Z9C
yZW1yaxJSZ0g3IjviIkwjwQkn5lMrYGn90pWu1g7GA7JyP0yc8tRhY/tVBW5U4dXdaudrubl9e4b
DS+LaaaP2ILqQeit9l/tGbQJxhIFyFSrkqgki/euxcVFTUk8KF7QQr5JBnu2nA+RgPN4t15TL94m
11YabjJol7klMM+TqMG8o0CGhqXKfG7LGGm5fC+j04nltq2kk5EKSmgNRxLIO+t/wCvNVsjzP8OY
dWvAeMnTWFTsnTJL5QPKQwxrOGFECdnpYgx3CX7cR7/6gACyzuH5A8lGCzT2/Lx3otdSQNOeXYfA
2YvkY7gpCrGj3Mu8jZSJ9QnlcxfPi6ZuP38P8AuaZhKEJp6L1lHPltLCDX4sVXeLwaESvZVnUhG4
YNnMMZU0eh3ZYHEQNmamLaDS3+78P9AzHA0iMe0bQcp0RT43RoNhc9MX2OjVaZqaGmj5Uhu9IlBv
L0VXhFDiTbeYJb7rP/G2EpAIE2SqgnaB6VEZG7Pk048dBeuEQa8WMl0Q01q3BdjkRzcX9bePkfqc
QLpMBe9tfqtvsot67BJ58QjrPK8z+b0arQHoeGnS4zJtsR3ftBYYnMYZ8n1ou06xM3VLgH6fpcGd
SyPU3dgRUybRJKdEE4T2Se1ayQAy5RmoFh6OZoXK75mrGyEUug1wEP/uKLhBpsZVcyksNfNstBuY
/7Xm4yKjd0iCBBZUK2deprXpWRMc5h7P0pfpdTB54vUzrp8SrRjGMz+haEHnPSGnyiX/bedwbndF
Oeh5HeriQ/zEyAaH6fxaKL7TsKMWeC6Yg76qfRhbSSgzfnZSECjs+Lw+br7qr/WMShgD0yyh+IMd
ViiIDi86cmGQdj7C3os3kqoaiSLhVcnLGdSF/5q8FTtl4Ox7GOalRXSYKv/PrlxrPrjSS0uSp/zq
YmvUJC6vViVkCGXGaWKa7T63rLXan6qCnqZ4uG6fT6YpVCnvEKQTWUng69XCjj9he4wtyND3TxUX
LM7HZCsKHcn8KAN6EHiQn3MGgfdi8f9T3mnUK0FNbYIe+iN0m0VPUaDisDmGBxGm1z1K/37j8R0q
3D7VBDTcR5H+3BTJAtVg+Xpt7Lri6Nh55+jCQi4fA5iPKSgIalK5PvkhO/odrvlo2SrYi0efRoKo
uKa3Ylgu0iPuoVZJqC+GXELO5pG8b3Y4HjCPZFKUKXj98Zdyuj5UdPXTKdoWo0LNBg2vkYlh6+6p
fpqGpnKslX0RNrZSBe2Fn97gn3LHegWiwbvC1TSNKd6va5nDJPU7G3SFaw8q443tHwajZRCvZXNt
cUmGZQP/7q+VdGfQh7zSHQ9wvr/HoXifeVioMc/uSIplh0cfBR4mL0jZ8zg2u57Qsn7CkW/ebMiA
TVHFWhhYW0bQhMvhUgXyYiLDq2XYN2PIyU26Ejk0mut7G7afETqQlZeYwA4rG2MBcmRxdaP+5jD0
ZyoyJ8mG7eIWTlHu6/FIrap47J2YOjRF3EfzisuYvb3/nzirTtPAyElaxUGMkCsdRhpb0LPPTJ3c
CzBvfBQyuudQCIqDv0VaWI0m/A0CgtFPihlZir1TUuWn/DXmuImTsSvC1pPMgHuAgvP9F66iNDsV
18z6RGuou5j8ORolZTVgbJ+0+lpHXt811gt9hWL1nLQoVnm6v04SSbp/cKJypLnFXon08NxpjXPi
RjCBT+lFwfLAsksHU5Ekr7muRC0JVi/vBbrwWV8H+WkUw5MJOVDfgWk2RHg+9QNnYxI82f8sYyfL
Aki9v3DgfoK47UdIJ3Iu97ypA34I+kYQp8t2s3At8a1PqmAtU7VvVDNAFdbw+pQyn7Bj+b3nuCIs
RKtomRKQPU7OKbVYl+oAm0wa7EypBHmzal6fEqA+7EPMkLeSpcQGtyAnPrFpQ66nCvZmUduaSO/j
Xi9tZ1mxCZn5FoRBZmYVz2J6quSCWwQEOyB64lfiX44yaiaBzSEOde5I/VyR/0yt/iv8rYI7Z6Up
jU0ZplK0oDk8sQVaeBCKMxk6PMmb5YNMmzDZ5S4YpPn9DOGIP5s23XzEbZihpJn8dI3aY1SL2p1v
2Bwgr+E/OmQXlCzvtF54E1RJor+mytjijd3mHcGKEwyW/xckVqbyQ2p/Ic92coxmVW45VGXad+Xy
9Qcm1Q5ssjymZnSASP5DmDkdIZc96Dkc4pbcK7gE9aD6lKCyAcHBBN3DVeL3GCOmwhUSnJPTl1Fi
us2wo94XTFfpEW1WWxEgQLfgqCkwcHkJgKf1OYiG8rwMBui2iHGondo6REwH+D8RfGbqOTgC4V7U
DIc0UreATrPtLeQ/BY/f1NII1xJMcKYLjv0mFg0s9hLPgZF7SmY/A3+QEQB7SUei5LcKCVZxddS3
LH3HT0anNT/GELOx8A7cB7V8DUiD679K0HMLw0ke+i5JGVVCbU7J/J9U+tOp7v8w3RY62MAmVGb5
wkHDenwc4KTq+imybdMNVPK3v6wxCVY7O7+1C02XvqMdHq7/TvI3hb7uXziTdwyKpgu53uHjaqYj
lEqxNO5OQuoZ1Edo9ZvN3tkA4YyARNqQ73d0fPHH/X4EBbKMOageaNVjNnBxdatUBmkuRAg+LL3f
Y3Sh3S3pkOwJs+bbuWdaeDMs+b15V7ybLcnwn1P2v4dt0QmVLuEh2wGPQNbJlu8h/nMW/gsNzOwH
A1JlcOuBqR8wlY7oAWyF1pgJ3IB7ai3MAQ7X/WZUHT9cDCFmM2JSUppNEaKPoqkNUfmm7KQNRVMr
D4MQdaTWdXZX6WI9P8b/D+aCTltDvkHdOomVwx1q1CPEtdaz8dAsSc6/IQnhLqwy7SmTl9goQRmu
cpUNEk10UtNrOB1KGn5QU2HUq2aejuLNls9zpa2AY9jdl7uV+ma6JPT1x+N+Ry4o44cfsKrtmCwE
bmAPonUHbh8ibZad/52jeVkDkNbAK3d8JE5i/mZE2HgW1MSbqj5LOO+YYBOxALQXsZa4PqxcM2fU
DY5esYBqjbWXB9DoxZM0Q5Lfwq7e3ulmbRuIE41ES4xJ/tzLYjPhopWYOQR2JWFTcWH0zxpeUg4c
480NTqf3eoyfpTk0jVypB//Wwc1RU/8X0vpKoPkwjrgXr3byY6hjij1rH/rQHMGH7EKLI3hKmtum
aBw5f5JwQTPWL6uKWwU1dKGsPVra3IACMn8oDZSQiUFSymG9Lv0hPBhNpub29zCb8tLePP712yPu
rBV+6EsX7qCaS9wgCUNh9VRHVWEO4p6Q/C+20ATz9qT3Q0sQsMMm/qL0dxJbhWJg7zRraFE75N1v
mB0v2+DcOsu23yYqhvCxyFY9nRMcCU3A8P5nO0BnEoh6KQ1qdcFL42zkOb3LJUW/1zeidgRJHyx5
bVmvY64WjQE4/2jJ2rGRHKpnkFTrjvvKtRDw4Zqn25rHeJvm/Cy+JzN1btYByD7oRBW6jOjD/AGP
OwbZHM4lGffgulpUWLeGcYXAYbazp43cEVdFR0rocjQBww5IxkYGWPUzE741zUxcuhd3/nZG8FRc
Mn3lh4oPjnbnYn+SVFk4sqarfZiIb59u9m+ThA8Lbm1z3M9HjswXm+wKkTSELYYyISE4jospv0hA
aWZyy5yqUmKrXulGu7yN6FCyOaX2BSptZb4o66+zZnswAJWBsW7Z80aAhULqZEOtKrh2hg4sAz1O
Ax2zfiB9mKSFZF5Me18ouLK/2lQIRsvvqB5Kp32hdhyArD7X7pD6R9A+PnU0BQF9upmtyhBPX1+M
Ur87aYV2QKB+7T1L1fH+hS90YDksOcIV+ACLAjYf8QrIASw22jW+aU2p51hpt55hfxg71UxO7VfB
uGxCymXcLViyAMFkmL4dXSXvwEiQl17NbqjTSrWUmVN2Iq34XZO++fl3vrNRMLmpsF3pc8x57+zA
gFxCByH3AL3K9Bkk80oFf5b7kilVt0oQcfZ4SS10Tylej5QRhuFHtM3B9iHvVt9MpD0ee9DInTuC
K/xAY3szb9j1hwvniVnQy5nn8v4DIgyoJAMe4k2HJN4q3ZRaXRnjkNGooanmd0PcAtoTiRgFDDCi
x+HuFodraMlVREGsdoX05gkGAw98FWRJFo8Ow9x61cyAglVRBNFFtDTCiRqCElWuXAMZlkCbTfgN
zx+Uh+kes49hr702tw7R5mr8QHBsa5IVbN6pxu/iz2li5fce8kivXWRk+QmAbnDMS7f2C74Dd3oj
xmwPrWcTiPDDVqqQzOJwEdoD2JUrzSpqnh0YAklLKacOxF2EK+scFhQgf2iJdGU0NAYBqLVUVzA5
w1GYwQ0neQTb0FiZIowFN1vwN4LH9kVbWumUgcuiA2P8yizysNDt45OPsajWftP54hE/DxspAIxC
3Bz8TTNAbEhzrRBviEskMbSKQ4ACN7Wpgje2D9WJ/+5UVe1iBPEl248YjeudFaxBd1fbTsVXZ7cR
HrRwyAYXllvJUyUDc59DzpFoJFqUtCNvu6hYRhO19irZz5jovCFJupAWsNSNqullXyAx0diTCfJ2
qU3syF/3Ld3BTmXreoYPKXji4/LLcSlAzrE6ispjIEN1+YRTjzaOb2L+th7hzzEO7XNeQtGYxrSO
lXY3AeMo9NN6JNkBeJqXc/tuJaexhL7igO8wAB9qLEt2G6bobFD1kBI+gYe2qVflkfkdyxuncohi
b7XjeLpdZ9W1sL+SUpfYUK9qD7kDh7w1u0XCXCtEL8K9yGCWMwSQcqjeI6tJ8UQ0oebEENjlQogs
CAIGtQcb806+oiII8vcVc3O1trNx6hU/O1HUECBqrcGi7xMCtDxcPU4patMJjW/5qxMO/DWfWPw6
/AWeZOIZ8em/O68UeSyRb5lEqv25hQrrFSlej5N+nn46D9xhwXaILTfN0Z7c54JNpC7REkoz3T4P
az2Zh1EXrrTCVnGgWPK3Fn3FYg80HhC3+Xa2a7M2bzgCi6YFAsSAnXKVSdGlsxWo8D+fR8ogfrap
xiQ4o0oJR8VB/fWTLiWDHdupfiYGVlbZHvRpssU437tRuLVmW60ISYJnVeJuddvC/dxgtOwfU4CX
8KxR5bgNo/4LslT7Kyvf9YfP5spx+66xpzh/7vhSDnmFEwUZRqLBPiqTKGAhiL8OjXze1hTlUwKR
II9zA9vE4KcvWjTCfvFNFrk/Wh21S32ty9zOqC4AZbKZ/l+MQHBl3tKsuZJI0VsGSFegW+WGXFmt
mCKtVFvT9FYEy+RkCAa410l+0MQy72MJ18EeblsqrUDPaW7jU6s3vie6XA235fTLuVsrQUNcjaOW
75/72I+tZGCcdNAz+BypvTJSQAki35Ia9HJAVEYPLImIAhGjcY3Xo+blnA4PrCy5Ok0q9/ej+mrI
pJB01vXJ7UzBsVcUeqidGUn+sHvjKCs3ksZEYs1RQjdtY48i6tHCHS21iN+V4h8JCQv+zILLsdVD
5UOFMFVXyI3jadT7xImtX90FGbtoe2lRHhx+hEkpsoPiI3hnFQ3J4GJV6rBk1LUAE2uEn1XkWxNl
ff489uO+yNnFUdpjTwXBBKA//m8NVRh7Empduha9xHQTfWCOrEqDSmRbRRrp4tWzBTHaMic4p23o
KtsqGwrJqSjzSjitX0lDtp+Zc/JMB53N69WWKZMRbz83SrhYBO8sMWWjihMNVJ8Kd07FwL2tsqHF
4dZwE45mU/DLt60GNtrBzU05xgkJE6/ibLqoKrFfdYL7NXKpO2a+kP01jHD0A24HawtNT/RZdlwZ
wIJuoQWxgZC5+vUjlPsQVZP6s5Zj0DLYQWv+6tGCFQMrrK35zEixBPB6x8rmwx52b5rYDGYAolIF
vtERvfCbJT9WdDtNYriVTE2JpHJYyvJ7EGmrX7E91dvMKyL4p+4osuKfpx9hziisbxNB0xz+Sj/y
qUvu76zDXTuaG2BsYkYlL4SAVEDg+L6kV9BWb74UH45g4IqM7VcP0HoKqUM6T0h/rcM6xsc7OCPm
KcbrcXLOyyp8EP8jnZvgMLONfjffjE2V/gNqoJBlrhkr32a3pZet2QWCnB1NfM1Y5c3hW+k6BZiS
nByoi8IK2xaTz/rTFpmE5LZJD0RHBWCEDPnpUWx/C72z2fWDtZyrQ+cxZzpKsPsmVt4kKA9B25u9
VpzNBo5yJbVZFm2wm3SkXQTkC2Hv+Y9cAg2UgmiyK4rMcD44kV7kr1BRZQZaTUD2pVQqCyUDA2mu
sa/m17q67UMtxV4fwl8ZNOYu6xIHRP2bSREUqL7iZtVufg7Y7YQXdoQO3O50u0pH/v7J9mw0tBfQ
nW2awzSx+t+tgCsZcsL1XNFRaOOWT1qdF4TeGkil70M3Xz/eQ0MwFZrWMExMA/VTV9J5MpYkGWEp
iz8eLo8WCfXM+9TS2MXidg4W6yDOc+4Xk5e9OwCbThRn8Wt7NVntjStRno8rkv/Bsb5XxtPYN3W2
kXLgKU/WY/u74zgxABbtZaYyZDq3OX4OrJJ9tXgCridiBuAG2H84svQwx1XItwHII0lgtkNiFik8
QNnBUC3urFyeb1dyKhZdHdsEmWmB1fLwfmm4WGjujrpDGPsKmK5pJFhr9kxu0jVoilF/zi9m693N
gc7Rrzy1A2R+mTAi6kSNiLwRrAlxhxcqnXQ6s69S7dVKDdHFSOwY05/sioGObUllY93JaggHbX/7
RUs0B+U8I5p1IGjaHQFnOeQfJik08oHRuA/FjKrJn7iU4FYcThwhyPRUeh8ehtIfQZnO1NQzrLza
Qod76fbB5dz7qW6FlqlFGWqJcSOPjGcU8iuxR8pj/Im1LfK7Q2ZbV+FeXARU4uC3whvoo+69fzEo
yTg6j3p2251kT9MLPgbPe0BAJhm0PrXzBpzIZgNPCD1Pn2/LX3aud+z7Jw/3wqykDzLdlj34qMse
lJfpLQrrAnMOoqjVc07ME8vK814dQZFauPF4Y51EAu4YvSUcBOZl/NxAEPEsiRg3a0/eLBIdvuTb
dWzZNIx9HY6hqbx8cXqrTqKpucX9nOIyn4Hs4DFEEV0N/zs7UvC3Skzt/XRU35tdDY6/KuT3Tpun
hVWzcZeKvMeqwPs83dfv26/orhzMZsLON47OBidF4YaXa0ulTn96hOAPfr224LazfFHFVTDqfd8S
fDxHCuv54AouQik0nEKM/6M9K1/niRs3Kd7v4vAvGBwsoJVWT2bIoBhxZUQed1fTmWimoHq1vb1p
wp01Ch/N8w9r1rPtD3I19kgSFudscEP4ZLJ9O2wPhmiQ/1bgtU0XHOEI2p6u85jm7O9E1ULQr62A
XP9fWVg7V3wCLskXCjG9xq5z1mV5iEztZfkuRYe7T65pWsnl2CCk1UFjYXKtZGZOM1XN+qmoExp2
WKvT74S2232oSmNDlge7tA+8CiExfo7mQVGbIGU2Cibs3sECbmuhBETTyNAZ8t9i5poEwo0mvzoJ
rakk2rUJVab8hFGe3/zSFg9WVJ/YGVaUEc/DED5smjtVJS2sEvDuEtPsByaV4EeaWmBQQD6eQBIj
54ABs2qaWKvCPnnYkzIH7o76bZrNrxglOG2FLxX9SgheYFfkCPjmy5iciR5XT2f6BzBQM9noyJP+
Vanye60HB7psii3/xPrVyLTMbrydZTaKQRrVj3on3yWB64rgSwBHokpmyF42caS5Qfktwvb5LAZq
+d0gP27fCqEyMotc6Ei2GqUCCmM8pV1v65EZNhXw7VawEFz7A+UaeIbcRYX2OeF4mMHoUW9SLJ14
auKOFjhFA6Q+UVIYKR50UyzUAC6r96uKKlQktJHtdbLAZWry+T4x9jgsBLT/LKvTgGikXJ7W3pJx
VU9c3BnNiKCqKd4WpDDrsBe4/aV/H/XuXmzw6l7zIPj7A5r/NM/DOr+UZ6G1lUKVuX4qq/lRt5Cg
vm/Z9wEZpMIIC0tSrOpdtihAUcjdmM7YC+DuG0h/3RlTQ6hZjVhWqoPHO7nHNPndyxQMl0i0IClk
x2YflFcEWuXjKZ7TSNWjCxmPPZaXFjF+MbIKdJx/9H7e4XwFahleIqZaHXGHW8kNE5OiAwNPQN+N
MuPAIFksyuGbOTJSVS8PfZFkkxMPDIp4QD7C0wp6SqSthPIJFpAKR4OJ0ZR2de8I4aoUZCH0VgA7
/uJMSwTbXa1mKsC+kZd56nhV+EToZ3yloQNrI7RV0zdoe8OdHBvcr8G589UP0y28iyL0BXea2/Aq
wHCLrexy0ppzQ6lzv4oIY9/C16dFyKN8QR2/7Tlk9ZncUc8djVHN6PXTj4gZMfo5wbjpHbI0FOnA
891CyJs4EVVhbigH63qYaRqDTpIIOaIveclRWLAbbTTW3bPxYiR6pGtIOou0NskG2vlHDs6GtN/M
g9H8vLiumo6twSr0KtQRGOVGOuHRdGS4IxIH9neK/koBnXxUeFjCvAX106TkdiQk3xTn6DokYpr1
KEIeAiioOiBQ9pTSbDapZjzlzDuoUOQtJyGQiYcMC//GZ9QSRr0jWU7Nv2RVagnkgcyrg/KGzgLb
L5NneksbgUW3Z5G6c65K+MdWC30WW3K/j5ZFG3ygNJf7dInQZQbn9CteBZue7O722FqBws06oQDc
n5w+uPjoHomAlwEE7poGsAFHQHaUfOX4SNwsVWh4xaM2Ettk7wcor2YwKHRjlqN3hK16urA/H+oV
R44Nxk26UzPyMyFTq6nEvWGZNDrS4VqwroDfTtUYM5zwVitGjY+pQ//3svbkKRQzZnidOUyBcK8E
2u7usWLKvOmljS+b/hQUW2AmWLJkejgQ811rtctsYrtFcnfeJk/TjtjWDPSmB0Dy6//5lSQnFUFN
/lQFoTxYkohMRGIuZFw21g4fBO1D7aIPYj9qaNvinT5jkGP2n1cPyoEU7BoEyIOv7iRCI6GmkXu9
JDHTGREgx6GnYqXgb+ilWHK5ITUItUzEKcmh1zLB/W5SLtbB3J9tR4Y4kW/MqTmFBHCQ4wMqQWdU
W7etQiak5RWqMXBoDJyefrKt0Zmdchm3Lr7q1QQBek2Pz3kRMkQltK/7NcN2YiXuAdflZ9AHzxrn
7ZPm8ranxqT9xwV6aon7g1Y2JRiaRip8Rb+1ejG1d2ZWL2ROVpbnu/Kx5p6/jDo+EbeQKyPRuVIJ
x++sZmC1YD3EDLVnroX40vbXNis2qL4+xyu+uHj053Tal69kSqzuqjOSojG/gZEIKTGUJQD9+Ru7
MPjp6nMOMAY4fLYoa5x+f2ESm524+wP6EymjEJnfxHme3PntGg3DYs9TLK90nj0Aoe3SHcyLaJh8
6/NYyR2zjEH/iXfw1rx+IQLsoyc/lE4liPosnkT6DFisuGnYstnd4IqcA2C20yTtSe6yR6pZ8KI6
VPmGCxgSIYGCXyA44iPVfC+6gv9IzhxHXLWPJq7pWGQLBSpkUlysMuuT4Fu27Bh3dy2ThE/4NzEA
zMueMe6pvLrx7MDZjZl/Fjl6EsTHiVeA+lpwibmdzoSLymI6RjLUcl/E43cpsC/5q+PuZQ5CsTAQ
BQkeShUc6lLYIcPOLl/fPkVA861kRx3jfgBIYSmx7WsT+a8HuQBjxSMKd65bXSj6YkTJvdqwMiCn
UW4/9oOFzLywu1Tvu2kmHPvXdo8Iy7VLby4ffH97uMHOZjCNGROmpv8OzXKPadZRYeqXUxTyQgE+
T6UMmzFa9EAYFs6ZZWFB5zhNWrErXUh+Ul7DHt7ansL19X9j+e1m1I5U8/Q1hzp7+HkXsCdWXHHn
caLvIOju6Cy0szgVtXGBieWjbv/goQ/gj6+cIhg8k8yVl+lN1/Tgjzz+VSin3CAUmawmV9zVoCUF
4MV5EJopumH1xFt95ruueRkdpagLQ+DxtPAzVZn/gSJdzTPss4nwLr4SnoWma688jBRaMoOm2Z6R
I8dQz8gAO/d5pLwOSvikpl1UsjU3bpNan3p5f99TbtTqzf7omMbupU/kNPuGxW9j3/YHGUAlgvno
7k8xQKyUV+CnwBLNpWXh1R5gRVPfv2a4w/n24LEd9XZejPcLxUFzCt2QVKJVtVfUIbmmWgJ/SypF
/mOzMhsWKbeJ2auHNM8exidZPAgaCiVuNj6isw7OcHWKwopfFXEyn64tLHgQX6ubS0FAwDKQ5nah
g1ogBXxwny65mzexxtjbD7/3Zc1tj/XbLNd0tGfXACkduUbNo+44DRF4PF8yXDXLrYirgIjSyURx
S4s0D9+OhDJ3T+SItE3NEjCIm35smux19p7ZkIvkNyk8y0dmlgeMXm9prgC7gaGl7djAN7ifvn7X
dQKzzUMWIxYRXrUTDxyTO4PpgSXQXAOXFVZDGHssSdKizoEsTTKOIC1wkpT4FFjT1PSt7MmqCFEc
fHTgdapEiRO7FXcR37WNrqGgsOcw+qk+KnNzg7CqkO7PyxX9fR6xjgQro7Cbs7y0vIiOYAdGVJna
jmJhy+b+R/OGIUvPQrPZlxW859YZiLTfrQcS6F+F+yDeBCtACz5zIQwVvTuOCg+wpJx+dfx4x/L4
tvUTSkM5BkE2oTxfD2R0OFAAg3er6UABKJaYGsaQH38yWSDzJK8nhnYjtMj+VM7PZeFo7jZQAu7n
HgMXcWQvTr/lMDeQh71Oxp42rUYxcVfCUE2nYwHnBw8iTSo2Sm9/zpZxZKD+fg0uZA9luqWxBT6z
v9Cxi2jX/pCYm23gL1PcXthz3Y61XkeJfjsbbWmlrW7PNOC96iM21RA6wJn2dA89fT1GUuErcAic
rvVu6EW1nGW/GsXltR59QKwEGNFGxXTQrn5Du1SGBrqw2fmDaCqxWHQKhbl4mndD+1P2VdgZos8w
rMzSZKX8tgyleSNh0aV5Dyh98bEltPwbufpU9FxPU1DKmhf6bKbi7SkBqY0dueNB0cdtcKDi1psA
ZqxsBIqA/dksBBL0tnwcKLOvxh+CTZVGnBi0e1CtCym7wg8ZDTdTgKMv0pM4zWEXAtYDq0BBPyrH
/RUPBtWBvOggEXuz1+UV6oTbIEUadN3fgMAR78umrl2jT2oQxNBAgcAwCeai2IQ4jhekfaBsA7U2
PdHNNQvhp2wUacOyxwgV4btTXM1Sotr2EYy0d9lSAml2k4ZzHwtBOhox9vCWqcfyQMrIe2COCWtu
48XjJZdY07o5IWOD9tVwwQGkciNa3Oag3OQNO31kO4J0xmPNzI+g+2dfMl2UqymdnSt1pGIGaCq9
uA/FGthc9zgZKk41kCckatVY87CVzbW+gQnplFTtm3WmEew3WtjlQPnTru2Yf+SNterwHhw0crfx
roE6LJwjuPCAxVpvTtiHF+SCOYpQAHS1O8A6Tbh6KAiowtMVEgKROgFoqgn8+KpKYW1Y4qloHBBC
Lu7q5rK65HjyICKpPk8pWwb4KQvftCWE2CrdpGeysCbxcY/gyFK096DiKm82ygqgWRA+ut4bWnBI
s+UfqRY/hD0ZUHIWqbn8JKITS561CwX4XuyrD6rpZPCKiJ267qD+IjGP2NzswMtdQchfiqDX/pPM
hYFhOKUQiGp3GkCSM4KCkGBj7lvBJiLs/w9qT0LDLkp5G/BBHsW2eFqj1YQt2PfMBf94FBG9FEH3
2km7ku3cmVhPh0fk5n3EqszgxsRpYnR/bPhAnkyjXGEk27X+vhQnCC8Y7cBtHMkWT3RaJy56XuFD
3fz/m2xGZs3scMZtUByjeth9+jtn2/hHvlQvn6yao+lPLsqYMf16NjF3TVYOMo6yiV4RlCOpOUTt
61fQ+cfGFAjNPRmX89zqPYY8XuW81nIKtTGeF4hBmaQ1SWSw+kfiN5vzG2OQtOxQpcHoI+J7YVgx
dbhwv50Z0y4IgHTTbCk0ZAzF/tBewbRvcpzf+B9cw2uoiD0hvdHYmVQYCyRlBHkW5xceTbybLbI/
bx792qMXAFg2KKND5XFpDwyAt6m+sS3VyQ+Mvi6JGUkPBKU8rOLpX1mDo3zZw4I2KNAIAM9y6Y2M
VzKozRFDN0ERY1XZqQLiUgq1xCez2zVyD5u1eknCyKHkEGBeOGoH0H9kTMmf7dyUFaMVCejoDuzb
BqHH/vpvQR3smg8aZBsqfqYBsUN+8UheKLsM+o8Y2yaX7v5PK6bVZXWAjDeopazbtyoIw/lhTFOT
iBNVry9BffKJPdG2QVqb1P5lq2ypkK8u5DEpRKsk6KiY9tP45tfLmjZ08c1zS9itrwLlH3r4vzWU
n72vHG7ANTSj+MemnNeXYB8MG0sDbXen2Rfyc6Grc/fQHZH8bG3dS+OlS7g+fNmAXukWwTFKA1Xx
o6Rcbk8wlROhv9d1+2ghz2uzKvhmxuHKk/3PNith/EbuxBm+mnjvxXcQwNpfYsff1qIGdN7M7mla
w/ziYG7dkB2+6BiT0osQ9ngUnCr3VFn+de1UqLasofE29OM5q1FDQGbzCURxfXTE/u5RgwJgIXPV
yjdtIUlfJOVckmuyNdwNIUJ1HpjmNOQG72rFFlwRGtaPsIOc38qfA4ndjhDbYWBrt2NkhvJgoIkW
VEfHf53+/Ff3mX0oboWNG5vdZPjQvnY82fbIjwNHroA6G9Pr551yPi9cgWYwjQKt1CQXVVN9lGUT
wntyx0NALoDlvyYtf5FuYePQGAt9GIvb9d+6Y+gfUZwejYOiAGsE+TGNUI4BqnM6EpLcGbJ9LVc4
Pg+riuWLqVdc+n4JD19uOMCKzE9ABPHKr0P2bVzx2U34wbSIDnMX92m5nkcE/zuwaX013BU67bEI
D4nCwDQaH8WnELnuWYMPPfJCXHRK7/x9+Kme/WL9m5qezyrxqacA6Hw7f6Gs0zVnlJKpxDvyPl+i
sixe0bI+Z7dAe8jStyF7GJAIEdx/EZ7x57x8mKhn38j6d+TExEHcaclx9ow2FXNEs8hMJUhXyQeE
DPOY6IJsTm/3I/8usYVLR9P5x32LpW/6q8Cq5xiAqTMla0ySP2QJXOY4DIru0yQvnhdRpFcQi/e9
aKJ7iVuvaEB8qhZCsmrURofrRWUv4d2bvfMXo7A+c/pYPvFxx937PXP31PYg41JTDzDeCjxe1AJY
Lu5bCmfvdyQr73pwcT1WvesQ1gaLNFs0NdZe9U86Dv1lbyApBXyS6onFLjzPMRa4POWVdZal46SE
Ovus6TnZ02PwS9c8zY+9k0d3Pf7HcHbM1x3HGVBqUxIXcvzIgpifWBkxB5gj4K4qAc7dCnOm1KLp
PJB5oaDJhIOw7DApEaQnB1ZLMcvXktIyFsIEIj9URS3fEWLaMO0pdgrJ8t0lQLhFUvhvX9g1Bqvr
qryPucvDNN2WRweuvwNH/nHlIvOrmRJmrKIq2z6V+CyoiciaHEO67hr5NJuM3PKZCITD6f3TtRC4
ba28mx+8Gp8p15sRuiBZPpyZxTehp0x0KzWGqAjYeTzYFnpEZNsuOHVqB7GKImJDdptkm4ke9MvF
rzXGRtKWbwtqXk4MuANhgiL+6AueEPg1c3F19KVrIZ7pIpgeWzFEuYFPdLKhJCXBvL+pF/xsWCEs
St86arFXxR1wP1/Hzow7bqHlORw3QhXw8ycqSJkzcXNp3EZotDFsAus9JtZEvYlxR/Nzn4hdczZk
5D81JShVw/Pzmb8fzMgkzciirvaQFY6x8Hb9jD1TAwO0yzB7/nmf8eQ7NNYjJbIUlZsLuGidqWXN
pwBG1Y9gR2AtJGf9Hz1aPfrWQNmCx2X5W+xsmJFu1shfQdPGepeCyOv9B1oIZ92G5Cz4d3mOpMZM
1ssIubC1liLNrvI5cIl2ohyH0wtzR65A6055sOootAYrxZtEabI1dVQJ+n15+jaol4dJ69wJsFtv
42vragdx+0U4dQkUMTwlBAkKJIihWJMY53JXYycfEisyLyszAVGFb54VZs239WmkF2jFLUJUYPIv
3aCQRt2uBvxNnRaPGH45mbJb6CyTGtU9jAaX016+UxkmGA8nGpLanoNn9CVdS1sDT6fsUw+bgI7O
rOkVBn5wW0aPkr6bXInZ76R+K9D3kJnfcFgsNOLp9fPkvjcsZMbs19xpDqL8LvZNCY6dziOMBgxF
E0yjfv7ZDmsnXysm9CFTwJ3+I0X/+H+3mzHNg5nu3Hm0b8uUbLqUx9v1rz5/yILjOlhe1feM56yL
puC+P+gfFOshsEC/+sMKgK69jSoQx0EzMr5QxiQX7hx/qdL0LpSbVOz0PH9+z02aJMtnLNbOPbTz
UhyhRNCKTTfWWGGGpPjTXFEb4/wvwsk2m+cvo80J5Q3rOFCM8ZEerRKM6jj56GYe+Mj3NfYwYBaO
8pEj76bIVa5BIXMBdp9JYt3eJK+RXFuCA3obJLIowqL/ZafvmRUWKSkaZ/vWkmqKjOMLZMceqJvY
jLopwLTX5gObiZh/BKM40tboose3/2YA2eUuLu+bw+rMrVZrrvK0IMI3GBWzcxrJHYE51CIfTm3A
9TNj4UwJTaGCUuUJ/b8eNSJ3AwjYpnDfd3QONIBNwnN2pSQAG1ngKnrQHa+Vk97tj5QMrRjG1gkE
0dZHa5u2EcVU3MbCULSzc7pjSqkghV7czYL4HNz3Y1gJSwYhs+i4gkDHMIUV8n2bnUacHs7nWFpX
1R7Oxh0EV/ZYT0xjhfcDmCzM33kqcZH9GZHU2t81s9rmTPBRy55n1UXhGUCzd+2r7t7dOUN4jjNd
rjCD2+zjQcdvmRhVBfty3ZzBm1m3VU+TAoZQPZCVm36f/gNqkw68YT+F4TGkHIRnu3dh3GlF1dam
eVln3pgJJw6Z8DhjJuFM648bVm8wDDQcxZT5uCM8LwijpO6WVIGe2TwTe/VKsJvm/lxz4zRXC+ZD
UO14fTzfLfQM4utIJyb6h1DiIWOlc5nk82tQhnhqNEifVdpy2OYTDgRBSswJgg0lDm9F6p6ncNUd
qJQfutzVnxUuFzyJE7VAtJM45Kjl9uroXII4GsSooEvdVpYsKwkGq28pNQrIV2vRIuCJB6Mm/+El
aNwaxXbrU+8fPZxXZSN6VIrNI75TO5d34gOO5GqArM2d+HPCVuDGcoOziKx1fwf+lnupwnvrd5TT
BU636IpefXCM+6ZzsUAD+F0OsQfA0SLFR5FhHcd2whmdZbyrQ2V02uyLM+l5ewozm78Fw/ZazWhV
mSdQNT0RT1dzflljptJAaj15tSUOS4hdg6QteDEn4myk/L5MFGJp2BGsN0Edn9S8TRCoDSUKEyAt
pzZHxZfJLLpbSk5IB6ElzlQNjtsFSh5yKMiwCmuckUNLcteJV/PON81n9B74kiox5zf9D0+N2U5d
jriU+TN7mJGcSgzB8b6FpJJWTymhFPd5xpI4OxLOCk/iLV046E6kzsrctdSNwY77AqbuXCzaBi5K
9RSoocyO4qb04p2tSBDI3gOVPU+lYO1N5DyrurrFHiUpldS5/ZHkClbMyullyE2fpOHincWYgCY0
CJ/xCllNB0S7Mrdgu32T2qkNBo8MynxtXNwNB7Bg2/VjQgZN7Qajon2vfpxZQVBa1hMxrmzqByDf
qJ24/D0KcwlHDYvZfvsYg5xdemE5HLDRQkXsbMZsbwElrX0n1hGt2ADG568jKgmeFPfSqsr6VtVW
PGwD0OpBfTaRKIeevYvdCj0iMmzmUaDXyeUGGC1U4PhClVyHOuYEI9tZyDPl23EoUQwoudRXCpqa
QG4j/FLBVOWLpvu6xQ7JuWG8+AxJf8ftwk60Y04UtIDUErXPNAIcEKK5wye3FnX8AeE/lWsSgs1Z
OKFwIbPb5LxDZN4sIU5NswEl8M9/hD1k9bqv+3FDxmRYoBsWb0brQaUc3ffkABJyL5JmxGmy+o9t
57s0fSzL0e0iGmMrKW3szTFEAJII0zvUQ0Mgy93842NV7bU9n2/cQ8zDL8u5zb/Joat9ernAcrDS
pVI/JmWtboTmf+u6IrzBfujMECLWrePq4B+n54stHwZEruGqoRysKQB3BqAY5QgfqADmYdzosTB1
SUDg2cy0Yj05XUTRxIUOHU+gLYrLGh4W4cjWNh3koHUXx4gg3qBc1mVous2IzHVCjcmLhdk4eSRR
Xss37YxA5DnTY8gzfCHqpSomnM8/rnDoyTNepkv0PDdHgRzDovP4blW0AL9YV4ln/fDgc/qEClOq
1S/1MwCuSRNmPWg7DKDKhpbr0QLaKPqijbM9Mf6wIlTADHg4GhJqj5coP6fNXu0S8jc1ThqJa+XD
WaKB7gHEakkQJ+Kh4uggYRxB+8OH+WO5LBY+58Be9M7GsA1+0Bl9N7pBC1/oWFOZaMWwNyqNakNO
yQD2JyVoujfPdcpTC7e6SKeIY5SsSBy3pDOf2kcxSP7UmGxhziDJ6Tw0X3pV4/j2TlL3l+HBRmPN
6DXBkrozoniYsVv6dvfAAn88Z8qK/j6crwnQ9WlpnjuqgTO1Qx9wcEx1KzI0NDPxD8RhL7jY/+QV
5jr5jbjnZO+iAEnm66huvjOH2sVSqCrjivKADwbK7ro+PClGXrW/qjpf9hQIumKFBht/upKT8L9R
1i4NrZYoPCTv1HdpPeBbAv8d/wFQFXHiK4W/t+1lCtqCLqPKA7Rjj1Mcyb8Q1aFi2RUygkETAQa1
5yDZ8ykrxc66JtK1nvO0OUXcs9+2GUPeUuEOKr/Qt50qyJGpBZ4FQHy6g1UxRcQHQ9fvvB6tFL2L
0u0GxXm15WZjwAK0Puljbep2a8Guy4kFRzVWJh62o0ivihf1wIA4mfJN8PS3pKJlRlM/lHeGTcw6
uIUbyfLoBVpZJNuwFgP0AHve7U/Za8WEddcm5tjYeU1AbXcrZWY4fxE2tzR9JZm3ijDlraH57FyQ
6gkjjSuHIdgTL3SBxiPOnJEI9owplBUtztKWgMngriLlb0c/vzzZrv956mfai8mM7MfuEpkujxd/
XF+vxPc2SKzhA3TxD7wrJKgYcStd5ZzfwPvEU6AY+zn0TaIRFfPsSeNzA58UCrKRukE0HfFAqJ5b
FF2UCVywSqyjECFf6oOUehmzi7zKLCcbe9MxYedxUktXuY934L5UFTUxJeNAvfmzb0sDCpu0RWXt
RNCBYRiNw/+CcKeNRcNIp4ZhOViGOKQO5H/tFxUypf6mZxfB7eZ+pcPbBqhgnkY/01EjJHd/TvdI
pj9hDsPooxcfwmPyZjHqucdUb5731RIFWmB3k5ePsIi5y3M3sbiZ28xfYibO+mr4COJYqDM680YG
aYdkjqHeXZcxPkqufU5EhdpqWlYQAxDPZm46tZ8u4GYl7yZFJixBRIrIqS7i8ylwHKKH3qvi/VXt
g/9rdBqrOxSOToE8VKNLSN2uL0kO35gmWYiYYVt/BcaN99l5pwK8urg8AHv9/cMYDV0Jv3hTB4px
bog6RJM6tqPNvol8kRG60yEdsP1zKnMwNVmkh+VYfzLN+sElSkGFh0Al/Wge99OB49ujUxNFVVRU
kbwxgVdTOCZF49/86Y/YzKBPFouj/irRixIWIUcu8XN1zzMsp2vxHgN4HazV+Fj/VPRbjLvhlxbW
i+LXoGM+H/OkTu8U9TS60AsOqbZ4TW9L5anadrljGcCIdbEPQz7lIiRHMn81SYrn7fLTFH/0TgZ/
bAOEYrlIm7zQXhKhxUN+QB5n29hZw+ScAn/OwbCjQIU9ZxIEeuIFhP3YnoNabQLt9Ra8p16Unyr0
7YLkNb16ArkxVver8P0HEb5ANazqOZARmcW1MfDyolg7hnt/hxm7G7kQkG+MzGYV4DGT6ShDp7F1
xjxlA6I2U92W1IiRIEnNwfom0R3Fm6Sq9mR06kdnsaZxRxWT6EUSnXSisu6+n0vAeZrbE1tf4+ss
tHl0PQJ2ODtbPKms1HonfxwXg1m6gBl9Q9XKjpmCTy5dMHb/c33GEk4161iNOLx5ycP2zdVhmQnO
UGu21EKx4R2L9OJ53q3WXs+79jKqxPTQILM7/NY53Jn17VUjalj11lfe4hrZoAlmXA3V8ojkPrp/
TsevjQY3hTHDRLt868Xc406sKXkvombdGys8LgVzKQbsktzzECzaxCW0D+SvvHo9zFOXEcYRVkmi
1EcOf+e5rgXP2zGfOyhSUCySPo1qzVzVDFatPwJozOPsHNws9MMxMbG0av+mtB2NaeUIiaMJTFPm
Bq6oCos2n9EJXi0HPvC4Y+80sjRDDVXYIip6P3PXp5jy8PIFBMppzpJUYw1GPGSLHCl1X6vtOWpY
6nz1gJHRpNuvml3f/Es+9M9usqwUMYtyO2HTMCEN90KQIF2vP8yvbZkmZHDe08rv/o+5h/FHUd7F
hE9Yq2axmhZtlkF3LFnUB1fw8CPPgzw9uMX44hd73t2meERwvZlw2nWf69I4rfFHbXpRaSIRtnyS
sgu8XyqnJnN26YC9YObMTnERtwf16US8z9IXnf10MBqNIXM2cL8U/eNhZMUk4FczaTcfqNBDVZxA
NxzRNsVbdyGJls+DqZ4ZX5TPrxT/w/2gKMb9V+1jsiUSWrLLd3YuI6LdXaLtc5H9BU3ayf1OHKab
r/3EgXUSmdEFgacpo7VtetcL7kESN7V2jWf6SCiZi9zFjaPyaDWpSyXcwMmgUTJHW+iUjPz9Uxhh
USNEYAEgaKPHC3D7IeJMkq2KYtnGmNSqrz2briX3eGRuihSMxkSh0gTgJgipvYKWNDD14s6tsRWR
53kP0kx8dGTIFmI75SoB0GM4GNkMH2F2OjnE2ELQYtNITmK1vRqntJrWZzhjwemvdCq1/ruNlb9x
OApCdAz8h6Bswv9VGaSw18P5QczhQKTIIZLnfoL28fuIRZxE2XVc743g207rV6xal79HVzdIlZ/R
bG4pKGTMNXGJ5YfclhIjJZdUj/yO/HpULpCMfQABTfNZnN7IDCcX7UfNLl7Ey/ZVtLs9rWDgACul
LlxdGvpjdaq+dQBNr7WhM3xo4JX3MxJlgUJ9z6jh7t9s/rQFE5ccd68yT6Z3FZVP7DdfiPEnFz5x
vGHKK/hCT56C5fROijzjdMio0INIQHWAfUZzOfD8rTb5u4xV84PueWLuBP79sL0rwkiXsTYz8q80
/Q47wqF/ArXvF1DJbM/OhkKxzJ03BBlmDXOusfp5yK3RB/VxghyScWDb/xWZDE1a15mM3C2AXBmw
PY9pXTyrbdd8g2ikD7rrImetrQtjXjK6MRK3mXG9AfrVF/9PF2lD7XqF5BY6aIu8m+w+vnjCVDJF
poq5PymU05YA05LyPRHIyhZYr9KEPukV94iB276AShhWMc2txTxufhFstDLj6QaqgojBOKIev3DE
hClMMqxskI7UGGo/Dv64ynvWBpzkHcW0FIcC0vpmo67vnRTL4kYNX5PatLakNej52W7+d1TJOWtf
VsugIVgVdqbs/PnzVTxceqnbUmT2gzNzrqEMSihGZ9g/LaBhVPZb+c1KPhbpx/4/JkSULZV+o8gG
W/fFJKMZgY9rFGKsO2vjk87o5Z4MZTsp8uY0VZrAsOei6zX2qReVK+Tj4RJi9oiJZv97g1SLAeep
4xGw0F7tILW8HclqFcjwnmUaOvolDLDiKwg3YkmiGY9TQkeyqk0HvpsfICqJwfw1j9rFVHOcmc9x
TMJ7GgJRV6b+gUjNASXRNjCUlRMtwdbJdvD7IZQc5yqff0EiLvaZXSlsBefdv12ySUDs9y+FmuIp
rM6UvklWZI4XYJX7gjkwMJicKGumGwjAwTXMjpVWAyUsi0ASw67DS3MaM2psFFOido24C9koSQ2o
Ow99vGFIp91sWf9m9HmIo9Ee514/Pxuhm3rgirxuWBKSnl/A4LUNALZGYox0B2FfhjOQcYsop9QS
L2/I7iXRNn7CdzIAz34hbR4/QRLcko0UdtZrl+p5whxnFn4UvwzWbeYNbn7dzVs5VYNmGMNGauRg
y5OplCEjCu3IpJf03SeVfIEi9dlL3VoYUJKwo29ZzVwc5gX9LjlSBT6Uc3mi4K54aKMzQK1w/9tp
6RRhINF+FWQpc8PDYlwQt7ZuTtfzZEflKPQBQTboY0eHkXsDEwQ58bT2/cyxHmsBb9iLyK4qVjiB
i9w6B2KVqLM9Za2iet6DkIeuvRQL24zlviDSxaWW4wK3VVo6S8eb6DQ0+JiSH7Q5rfWPZzaD4MDP
kKlkz+9aCr1LAJ0HueiGalYo2iVZ9kXLlMDiwPUsYMmeqLH9EurBsAtQfRqXiUmUPITnuePTNhms
h6+v4yKY51AxKm1WgieZ1et6MmVYNbLJWbw3BATKuxTvN6hZz6FkooXUNzbJDUJb0uNYSZllKvZ3
cb9TczYnfOXMNhqkhRwHgYiLEbc4SwwmFFWkicAHZLXVCbaiYNtL+Jk/rKcMwm3R+bowH+HxGmFX
ld2CugLobQTVcgUZ/bu6AuthE3rtKl9u4vvLq65sKCbIFYFMsyfvwisAF8jwgWr8X3zTr1vzcnET
gJidmju+TUFPet5MDZZYo36KZBBRxHuFwIrJOyQ+6IT4N7vVN/cZjpjxnv0Nqawj+W1jc7py+z/7
yUMLbVTM7uEppgN2KkKQlcIEd679mRD2nvhG67P03IuRImnH1MRmFbSXltvlYE/5wL/q7uTcOpGL
GrPi2Rp5QuOr2Sx2v1kfoyPmNZvCcdxTqJs0Pb/O4ooPoHrgSbxuvttS7tctEj9VtJNODrLuI1Sl
DgmW65CQcKfMSIxwSalcFulSX2t4n4ZT3TFNGgjfNHWArAABj5lCJcep8D89dT6+SgK3VWMhFW2F
xmJOizosYFMnWfHpYcig34eK2nuz5clJIq7T71p0mIT4QIAeVUUxhEOlI8XGksmRm69ynsu5uSFB
CzidtrmTlYqkAIRdAtF5RSS3eyy2Gal7NyITqsVhxw+uUS4nCVkcu7CHyS2scRyWhBTulP7qdcFu
iFO7DMh35+rUcwefcp4y+Pq1mcH31fW7Y+triPa4kX/RXeMyR7P1tHD1Lu99J0QW2GyhqVn6gbD+
h6HU1fsFmVsuIXl78HLVTwAe21CZcvnWImFq77fLPpn9zCMBfj9P8XrDy0OjKKy5Zgosu9Tkawug
TBaZZ0GebQVDM1RLN9j3PEg0AfwhfXY7nq6ZhXS+QQa+Wd9FhtkhepV0iyKrw9Pn5Tyzv+Vydtc/
m4J9jBbdoyZb0U2O82S8AaM9KzbAsf3F06SAaoe/rmrCLce7TQaGptkdLe8OlWnNbsy/+C/rrxPt
mA34AvekWXnhWpw612XA+01Q2iqq1MDrIpBSc4Dwv0m9WAaCWPE2Stf0MPN2CHk8nq5uf1AUT+OB
wnpNj59v5PH4sqa/S8LDPlLFtUNnimS2yoTiT2DTmbIb+ZvNzE9cah6vdrJMl1RkIgEVu0yfpZog
PT1x8Ald2u9KrmUB3hmRfGF6PAnEpQf/arW8ntGmRAHf7fvmmiZzU44SadtqGnV+9PwwBxRFnp4g
7LSv8s3Dwg4j188Y9z3+OssqKhAiFtV+c/wFD0P/P0awvekdBuYW1pIGJSBUOpYzFF8n2UkZNZ36
uzYA5uwG+mBtXREuy0H7eTF+ZObMCo0BHFwT8ZTKoHT0RXCu3jngt/4qhtsnOIkl+myXbsybQALg
IbACitrHi/sakJ1XgY8coI9rTFuuCaeFcwIKt3X1mhOw+MRunc14Wp1mqOd/JfmdQS58wopBEipR
PQxsn5evSUnG9zXS3U7VppeB5mVp43SD2SEQqH9qZQOkdkEkescj32eCykgBab3vOuK4/VDOnHU3
VzNFPfLwCrol9MTA9s18dUOB4vEUUNgoBjPxUvQm7p5kWbEEehWy9/ilVYGWPbAhYELkX8GQG9+m
f6SKe04VJslRKCbOxRHxWtg/IQjALZJU1CtJCk3h42kK85ECcMxT3Ub3Loksto0GEKExhklRuvqF
LradiGNHZpGzQyVs3etps9YERhweKmwYTllbrEeic60u5NInuqc/j7LFCFkNufoOVL5HC8/Y7+bU
Pzc8DUzT9scVev8z/S8i4PPhcH7u5y1a2dLQt6AhFDVwV8jNCVRktvNaX6KrYsf+DBMmt8t9NCvg
lBQRZj8luKba2eOC+eVmjq6ikkMiiyjgrkA4NVA/bc85DhcMHago3e8xzgTNl9eB4LfAIq4Ii3BQ
0Bx5afqCCXXR2y2ne94Gvdec8OwDELrukNv4FD58hQChw9mVHc2kLej2D25VkIwdP72wbFB9bJL4
1zqSVEnxjuo29sk0C07ALv28ZN69DliXikL/bXty3Q9Othc1JJeiNu7a7QffUERSzeOVlnNRGNce
+tHyJMAVksvcN7LyZtBp247dSI6J9UsuIIX38CIV2Mvzy1TS2bqbb0dmdXOJHlSm64BsbgueASnz
4PgskDMB/W4gicYse5Nxf9iHiH8dXgv2dbdrllP6WCI6dJq5aYm8mEmrOglJQzT2i15RQ2EYSWgD
Ot/Kl0i76lLc7d6IXTR5fl+/Y5n316A4zMAPabzoSilBD5EgN0HG3Fjv0PfSTqwGqw7A1JEdSbc6
6+pG13ObeiKXcVWw/QwiaynXO8Nyzd8a1WuuvkrjKYG2KIQfVxMjQ9QqYy0leBy3A6xcS1kZoD5x
z0Fuc9XP94sxv3DtH+jlMewIgwwBQ0dU5qYzi658cE/iK/Y1Eq7qjBZ7FiJPXflz3RAjE94TDlmB
l2OF5q498n6vDZ/f4m3Z8iQc43eOF/2LI57abdxJnid4qOFoFEMjuxpN0/RQGtFXefk3KGOOAlss
R5g78arSscRvt7WhPC4LsxlJ7TaUhuKICEcugaiaz6gq3Jf4lPtyygPmpmVF8wbHr40zky+R2jg8
iq+3ZryNgXJqojj77ELnnhWnJ6s/FN9Fgz9IVvLZe0bcan+MMHbd8e7NRYxEDGNBmXdJ9y8D81bZ
UPScuMBa93U9IIMYlNjvvDjybT7iAl8gJOXoE9lbTAzJ1GZ3JKivaHbkmuz9XH8twJ35Yh0gXfYy
W6ooKH0+7+7lZaj2UusB5wjyvhRpSCiyKMlqQF8ldp5lw1sB7RRZaoKPm/Q8Wl6nDdcNmcW7mkZY
VsGWuMce35lOcCg/faB9gEY8ZDHHS3LtKgATKPrqsUnqczBPdWAQchB2hUHinpLlyYYiQXDj0uJo
sICOuK+d2Y6PruBXTVyoW0GNMClEYdr0pTXLw4t759SHJm1zmN70C0/7/xaDx6GORS/ST/QLYTGk
TIQYw6K4U9Wz8H/DS0lpq0zSvcvjuMSvwQpy03NmLz07Dp6B5tt0V+e8PM4x0I3AVaL8OSXTaKEC
5jv7WSlTVh4yhmu/GUAskfU5bZRzsWkyIHcsHSDhumbNCMVqMGKa5YMoxX512coFd/IB3LE+9iWC
G+YABxqdQG0S8LNKFTb2JgcjUEVNGiQGHFAiGGomA7vFO5g11rCUiW/M8QSAfYeazG7TGluJ/Kit
tkUG6WuYTWNqqWUO1G6qoQ1ho3VLmuVpqsht4+Kb1Hd79aXQ02O4Rb1f5xsj/r1G/6+VOb0eEpvK
u8HcKnSSFzaiUHk5fsYumkop0T3HdmjJxeD1VfDKYi4XPcsjPk9yJAPC8jiHORjaviVy4sKIKzAh
8kD2ORDQsqPDFvqn75/xK2ao6lTYFTSg7B0Vnws5dCooLrnVGa8iyk8Psb/ZERuRAI1mlxrUu3ZN
+5Ylce1RXwo+uVe+XyPcSixzIxJjJxNRgW1nm6RmsH37DV7uPZpcblEGEc/+hJNWvR4IiaTOrsZA
7PciZ5KELzW+LDgpmwAx2qiQBII1LzKa37z1TrgP+xjP87QcTu1Qe2ao6L/v2og9rYTxLptszYVv
ed0nyECyPS0eRpliggEUkbLIuOJhWxounpF6itkiU64rKmEmDZ5xP33IP9fbODymt6seTz9A/WKL
Iyr5rNxyMoqGtFApw5oVn2cp9tiwdcGhJd9KieTuhJzKz4P2xz1DuQQDRCFDmp6mnSFWkw/ZFgD7
2X1D86+rpjCCW2vKeYz8FTIGKafR0kBAJW0BE3MHYzlJC58Lj056r4+LQVkGVa2fdMk9IiiEQ65K
xP7sHpeRnSzBSVuJ0mgwLnpi5wJM4pNX2V9d
`protect end_protected

